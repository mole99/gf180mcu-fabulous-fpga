magic
tech gf180mcuD
magscale 1 10
timestamp 1764324363
<< metal1 >>
rect 672 56474 27888 56508
rect 672 56422 3806 56474
rect 3858 56422 3910 56474
rect 3962 56422 4014 56474
rect 4066 56422 23806 56474
rect 23858 56422 23910 56474
rect 23962 56422 24014 56474
rect 24066 56422 27888 56474
rect 672 56388 27888 56422
rect 3614 56306 3666 56318
rect 3614 56242 3666 56254
rect 5182 56306 5234 56318
rect 5182 56242 5234 56254
rect 8990 56306 9042 56318
rect 8990 56242 9042 56254
rect 10558 56306 10610 56318
rect 10558 56242 10610 56254
rect 13022 56306 13074 56318
rect 13022 56242 13074 56254
rect 14590 56306 14642 56318
rect 14590 56242 14642 56254
rect 16494 56306 16546 56318
rect 16494 56242 16546 56254
rect 18510 56306 18562 56318
rect 18510 56242 18562 56254
rect 20302 56306 20354 56318
rect 20302 56242 20354 56254
rect 22206 56306 22258 56318
rect 22206 56242 22258 56254
rect 24446 56306 24498 56318
rect 24446 56242 24498 56254
rect 26014 56306 26066 56318
rect 26014 56242 26066 56254
rect 7410 56142 7422 56194
rect 7474 56142 7486 56194
rect 21746 56030 21758 56082
rect 21810 56030 21822 56082
rect 1026 55918 1038 55970
rect 1090 55918 1102 55970
rect 3042 55918 3054 55970
rect 3106 55918 3118 55970
rect 6178 55918 6190 55970
rect 6242 55918 6254 55970
rect 8082 55918 8094 55970
rect 8146 55918 8158 55970
rect 9986 55918 9998 55970
rect 10050 55918 10062 55970
rect 11554 55918 11566 55970
rect 11618 55918 11630 55970
rect 14018 55918 14030 55970
rect 14082 55918 14094 55970
rect 15586 55918 15598 55970
rect 15650 55918 15662 55970
rect 17490 55918 17502 55970
rect 17554 55918 17566 55970
rect 19506 55918 19518 55970
rect 19570 55918 19582 55970
rect 21298 55918 21310 55970
rect 21362 55918 21374 55970
rect 23874 55918 23886 55970
rect 23938 55918 23950 55970
rect 25442 55918 25454 55970
rect 25506 55918 25518 55970
rect 1374 55858 1426 55870
rect 1374 55794 1426 55806
rect 672 55690 27888 55724
rect 672 55638 4466 55690
rect 4518 55638 4570 55690
rect 4622 55638 4674 55690
rect 4726 55638 24466 55690
rect 24518 55638 24570 55690
rect 24622 55638 24674 55690
rect 24726 55638 27888 55690
rect 672 55604 27888 55638
rect 22990 55522 23042 55534
rect 22990 55458 23042 55470
rect 21634 55358 21646 55410
rect 21698 55358 21710 55410
rect 1038 55298 1090 55310
rect 19966 55298 20018 55310
rect 3490 55246 3502 55298
rect 3554 55246 3566 55298
rect 6290 55246 6302 55298
rect 6354 55246 6366 55298
rect 12786 55246 12798 55298
rect 12850 55246 12862 55298
rect 18274 55246 18286 55298
rect 18338 55246 18350 55298
rect 1038 55234 1090 55246
rect 19966 55234 20018 55246
rect 20526 55298 20578 55310
rect 20850 55246 20862 55298
rect 20914 55246 20926 55298
rect 22418 55246 22430 55298
rect 22482 55246 22494 55298
rect 24882 55246 24894 55298
rect 24946 55246 24958 55298
rect 26226 55246 26238 55298
rect 26290 55246 26302 55298
rect 20526 55234 20578 55246
rect 2494 55186 2546 55198
rect 1474 55134 1486 55186
rect 1538 55134 1550 55186
rect 2494 55122 2546 55134
rect 6862 55186 6914 55198
rect 6862 55122 6914 55134
rect 11902 55186 11954 55198
rect 11902 55122 11954 55134
rect 17278 55186 17330 55198
rect 17278 55122 17330 55134
rect 25678 55074 25730 55086
rect 25678 55010 25730 55022
rect 27246 55074 27298 55086
rect 27246 55010 27298 55022
rect 672 54906 27888 54940
rect 672 54854 3806 54906
rect 3858 54854 3910 54906
rect 3962 54854 4014 54906
rect 4066 54854 23806 54906
rect 23858 54854 23910 54906
rect 23962 54854 24014 54906
rect 24066 54854 27888 54906
rect 672 54820 27888 54854
rect 22542 54738 22594 54750
rect 22542 54674 22594 54686
rect 23774 54738 23826 54750
rect 23774 54674 23826 54686
rect 19630 54626 19682 54638
rect 1474 54574 1486 54626
rect 1538 54574 1550 54626
rect 25554 54574 25566 54626
rect 25618 54574 25630 54626
rect 19630 54562 19682 54574
rect 21198 54514 21250 54526
rect 24098 54462 24110 54514
rect 24162 54462 24174 54514
rect 24882 54462 24894 54514
rect 24946 54462 24958 54514
rect 26338 54462 26350 54514
rect 26402 54462 26414 54514
rect 21198 54450 21250 54462
rect 21522 54350 21534 54402
rect 21586 54350 21598 54402
rect 27010 54350 27022 54402
rect 27074 54350 27086 54402
rect 1038 54290 1090 54302
rect 1038 54226 1090 54238
rect 19070 54290 19122 54302
rect 19070 54226 19122 54238
rect 20638 54290 20690 54302
rect 20638 54226 20690 54238
rect 672 54122 27888 54156
rect 672 54070 4466 54122
rect 4518 54070 4570 54122
rect 4622 54070 4674 54122
rect 4726 54070 24466 54122
rect 24518 54070 24570 54122
rect 24622 54070 24674 54122
rect 24726 54070 27888 54122
rect 672 54036 27888 54070
rect 1038 53730 1090 53742
rect 1038 53666 1090 53678
rect 22430 53730 22482 53742
rect 22754 53678 22766 53730
rect 22818 53678 22830 53730
rect 23538 53678 23550 53730
rect 23602 53678 23614 53730
rect 24658 53678 24670 53730
rect 24722 53678 24734 53730
rect 26226 53678 26238 53730
rect 26290 53678 26302 53730
rect 22430 53666 22482 53678
rect 1598 53618 1650 53630
rect 25678 53618 25730 53630
rect 21970 53566 21982 53618
rect 22034 53566 22046 53618
rect 1598 53554 1650 53566
rect 25678 53554 25730 53566
rect 27246 53506 27298 53518
rect 27246 53442 27298 53454
rect 672 53338 27888 53372
rect 672 53286 3806 53338
rect 3858 53286 3910 53338
rect 3962 53286 4014 53338
rect 4066 53286 23806 53338
rect 23858 53286 23910 53338
rect 23962 53286 24014 53338
rect 24066 53286 27888 53338
rect 672 53252 27888 53286
rect 27122 53006 27134 53058
rect 27186 53006 27198 53058
rect 23202 52894 23214 52946
rect 23266 52894 23278 52946
rect 26450 52894 26462 52946
rect 26514 52894 26526 52946
rect 1598 52834 1650 52846
rect 24658 52782 24670 52834
rect 24722 52782 24734 52834
rect 25442 52782 25454 52834
rect 25506 52782 25518 52834
rect 1598 52770 1650 52782
rect 1038 52722 1090 52734
rect 1038 52658 1090 52670
rect 23662 52722 23714 52734
rect 23662 52658 23714 52670
rect 672 52554 27888 52588
rect 672 52502 4466 52554
rect 4518 52502 4570 52554
rect 4622 52502 4674 52554
rect 4726 52502 24466 52554
rect 24518 52502 24570 52554
rect 24622 52502 24674 52554
rect 24726 52502 27888 52554
rect 672 52468 27888 52502
rect 21982 52274 22034 52286
rect 26226 52222 26238 52274
rect 26290 52222 26302 52274
rect 21982 52210 22034 52222
rect 1038 52162 1090 52174
rect 1038 52098 1090 52110
rect 1598 52162 1650 52174
rect 1598 52098 1650 52110
rect 21422 52162 21474 52174
rect 22754 52110 22766 52162
rect 22818 52110 22830 52162
rect 24882 52110 24894 52162
rect 24946 52110 24958 52162
rect 21422 52098 21474 52110
rect 23774 52050 23826 52062
rect 23774 51986 23826 51998
rect 25678 51938 25730 51950
rect 25678 51874 25730 51886
rect 27246 51938 27298 51950
rect 27246 51874 27298 51886
rect 672 51770 27888 51804
rect 672 51718 3806 51770
rect 3858 51718 3910 51770
rect 3962 51718 4014 51770
rect 4066 51718 23806 51770
rect 23858 51718 23910 51770
rect 23962 51718 24014 51770
rect 24066 51718 27888 51770
rect 672 51684 27888 51718
rect 25678 51602 25730 51614
rect 25678 51538 25730 51550
rect 1598 51266 1650 51278
rect 24658 51214 24670 51266
rect 24722 51214 24734 51266
rect 26226 51214 26238 51266
rect 26290 51214 26302 51266
rect 27010 51214 27022 51266
rect 27074 51214 27086 51266
rect 1598 51202 1650 51214
rect 1038 51154 1090 51166
rect 1038 51090 1090 51102
rect 672 50986 27888 51020
rect 672 50934 4466 50986
rect 4518 50934 4570 50986
rect 4622 50934 4674 50986
rect 4726 50934 24466 50986
rect 24518 50934 24570 50986
rect 24622 50934 24674 50986
rect 24726 50934 27888 50986
rect 672 50900 27888 50934
rect 26226 50654 26238 50706
rect 26290 50654 26302 50706
rect 1038 50594 1090 50606
rect 23874 50542 23886 50594
rect 23938 50542 23950 50594
rect 24658 50542 24670 50594
rect 24722 50542 24734 50594
rect 1038 50530 1090 50542
rect 1598 50482 1650 50494
rect 25678 50482 25730 50494
rect 23538 50430 23550 50482
rect 23602 50430 23614 50482
rect 1598 50418 1650 50430
rect 25678 50418 25730 50430
rect 27246 50370 27298 50382
rect 27246 50306 27298 50318
rect 672 50202 27888 50236
rect 672 50150 3806 50202
rect 3858 50150 3910 50202
rect 3962 50150 4014 50202
rect 4066 50150 23806 50202
rect 23858 50150 23910 50202
rect 23962 50150 24014 50202
rect 24066 50150 27888 50202
rect 672 50116 27888 50150
rect 25678 49922 25730 49934
rect 27122 49870 27134 49922
rect 27186 49870 27198 49922
rect 25678 49858 25730 49870
rect 24658 49646 24670 49698
rect 24722 49646 24734 49698
rect 26226 49646 26238 49698
rect 26290 49646 26302 49698
rect 672 49418 27888 49452
rect 672 49366 4466 49418
rect 4518 49366 4570 49418
rect 4622 49366 4674 49418
rect 4726 49366 24466 49418
rect 24518 49366 24570 49418
rect 24622 49366 24674 49418
rect 24726 49366 27888 49418
rect 672 49332 27888 49366
rect 1038 49026 1090 49038
rect 24658 48974 24670 49026
rect 24722 48974 24734 49026
rect 26226 48974 26238 49026
rect 26290 48974 26302 49026
rect 1038 48962 1090 48974
rect 1598 48914 1650 48926
rect 1598 48850 1650 48862
rect 25678 48802 25730 48814
rect 25678 48738 25730 48750
rect 27246 48802 27298 48814
rect 27246 48738 27298 48750
rect 672 48634 27888 48668
rect 672 48582 3806 48634
rect 3858 48582 3910 48634
rect 3962 48582 4014 48634
rect 4066 48582 23806 48634
rect 23858 48582 23910 48634
rect 23962 48582 24014 48634
rect 24066 48582 27888 48634
rect 672 48548 27888 48582
rect 26450 48190 26462 48242
rect 26514 48190 26526 48242
rect 1598 48130 1650 48142
rect 27010 48078 27022 48130
rect 27074 48078 27086 48130
rect 1598 48066 1650 48078
rect 1038 48018 1090 48030
rect 1038 47954 1090 47966
rect 672 47850 27888 47884
rect 672 47798 4466 47850
rect 4518 47798 4570 47850
rect 4622 47798 4674 47850
rect 4726 47798 24466 47850
rect 24518 47798 24570 47850
rect 24622 47798 24674 47850
rect 24726 47798 27888 47850
rect 672 47764 27888 47798
rect 1026 47406 1038 47458
rect 1090 47406 1102 47458
rect 24658 47406 24670 47458
rect 24722 47406 24734 47458
rect 26226 47406 26238 47458
rect 26290 47406 26302 47458
rect 25678 47346 25730 47358
rect 25678 47282 25730 47294
rect 2046 47234 2098 47246
rect 2046 47170 2098 47182
rect 27246 47234 27298 47246
rect 27246 47170 27298 47182
rect 672 47066 27888 47100
rect 672 47014 3806 47066
rect 3858 47014 3910 47066
rect 3962 47014 4014 47066
rect 4066 47014 23806 47066
rect 23858 47014 23910 47066
rect 23962 47014 24014 47066
rect 24066 47014 27888 47066
rect 672 46980 27888 47014
rect 25678 46786 25730 46798
rect 27122 46734 27134 46786
rect 27186 46734 27198 46786
rect 25678 46722 25730 46734
rect 1598 46562 1650 46574
rect 1598 46498 1650 46510
rect 2494 46562 2546 46574
rect 24658 46510 24670 46562
rect 24722 46510 24734 46562
rect 26226 46510 26238 46562
rect 26290 46510 26302 46562
rect 2494 46498 2546 46510
rect 1038 46450 1090 46462
rect 1038 46386 1090 46398
rect 1934 46450 1986 46462
rect 1934 46386 1986 46398
rect 672 46282 27888 46316
rect 672 46230 4466 46282
rect 4518 46230 4570 46282
rect 4622 46230 4674 46282
rect 4726 46230 24466 46282
rect 24518 46230 24570 46282
rect 24622 46230 24674 46282
rect 24726 46230 27888 46282
rect 672 46196 27888 46230
rect 1138 45838 1150 45890
rect 1202 45838 1214 45890
rect 24658 45838 24670 45890
rect 24722 45838 24734 45890
rect 26226 45838 26238 45890
rect 26290 45838 26302 45890
rect 1598 45778 1650 45790
rect 1598 45714 1650 45726
rect 25678 45666 25730 45678
rect 25678 45602 25730 45614
rect 27246 45666 27298 45678
rect 27246 45602 27298 45614
rect 672 45498 27888 45532
rect 672 45446 3806 45498
rect 3858 45446 3910 45498
rect 3962 45446 4014 45498
rect 4066 45446 23806 45498
rect 23858 45446 23910 45498
rect 23962 45446 24014 45498
rect 24066 45446 27888 45498
rect 672 45412 27888 45446
rect 1598 44994 1650 45006
rect 26226 44942 26238 44994
rect 26290 44942 26302 44994
rect 27010 44942 27022 44994
rect 27074 44942 27086 44994
rect 1598 44930 1650 44942
rect 1038 44882 1090 44894
rect 1038 44818 1090 44830
rect 672 44714 27888 44748
rect 672 44662 4466 44714
rect 4518 44662 4570 44714
rect 4622 44662 4674 44714
rect 4726 44662 24466 44714
rect 24518 44662 24570 44714
rect 24622 44662 24674 44714
rect 24726 44662 27888 44714
rect 672 44628 27888 44662
rect 1038 44322 1090 44334
rect 24658 44270 24670 44322
rect 24722 44270 24734 44322
rect 26226 44270 26238 44322
rect 26290 44270 26302 44322
rect 1038 44258 1090 44270
rect 1598 44210 1650 44222
rect 1598 44146 1650 44158
rect 25678 44210 25730 44222
rect 25678 44146 25730 44158
rect 27246 44098 27298 44110
rect 27246 44034 27298 44046
rect 672 43930 27888 43964
rect 672 43878 3806 43930
rect 3858 43878 3910 43930
rect 3962 43878 4014 43930
rect 4066 43878 23806 43930
rect 23858 43878 23910 43930
rect 23962 43878 24014 43930
rect 24066 43878 27888 43930
rect 672 43844 27888 43878
rect 25678 43650 25730 43662
rect 26898 43598 26910 43650
rect 26962 43598 26974 43650
rect 25678 43586 25730 43598
rect 24882 43486 24894 43538
rect 24946 43486 24958 43538
rect 1598 43426 1650 43438
rect 26226 43374 26238 43426
rect 26290 43374 26302 43426
rect 1598 43362 1650 43374
rect 1038 43314 1090 43326
rect 1038 43250 1090 43262
rect 672 43146 27888 43180
rect 672 43094 4466 43146
rect 4518 43094 4570 43146
rect 4622 43094 4674 43146
rect 4726 43094 24466 43146
rect 24518 43094 24570 43146
rect 24622 43094 24674 43146
rect 24726 43094 27888 43146
rect 672 43060 27888 43094
rect 1038 42754 1090 42766
rect 1038 42690 1090 42702
rect 1934 42754 1986 42766
rect 24658 42702 24670 42754
rect 24722 42702 24734 42754
rect 26226 42702 26238 42754
rect 26290 42702 26302 42754
rect 1934 42690 1986 42702
rect 1598 42642 1650 42654
rect 2370 42590 2382 42642
rect 2434 42590 2446 42642
rect 1598 42578 1650 42590
rect 25678 42530 25730 42542
rect 25678 42466 25730 42478
rect 27246 42530 27298 42542
rect 27246 42466 27298 42478
rect 672 42362 27888 42396
rect 672 42310 3806 42362
rect 3858 42310 3910 42362
rect 3962 42310 4014 42362
rect 4066 42310 23806 42362
rect 23858 42310 23910 42362
rect 23962 42310 24014 42362
rect 24066 42310 27888 42362
rect 672 42276 27888 42310
rect 14130 41918 14142 41970
rect 14194 41918 14206 41970
rect 1598 41858 1650 41870
rect 1598 41794 1650 41806
rect 2494 41858 2546 41870
rect 14578 41806 14590 41858
rect 14642 41806 14654 41858
rect 26226 41806 26238 41858
rect 26290 41806 26302 41858
rect 27010 41806 27022 41858
rect 27074 41806 27086 41858
rect 2494 41794 2546 41806
rect 1038 41746 1090 41758
rect 1038 41682 1090 41694
rect 1934 41746 1986 41758
rect 1934 41682 1986 41694
rect 15822 41746 15874 41758
rect 15822 41682 15874 41694
rect 672 41578 27888 41612
rect 672 41526 4466 41578
rect 4518 41526 4570 41578
rect 4622 41526 4674 41578
rect 4726 41526 24466 41578
rect 24518 41526 24570 41578
rect 24622 41526 24674 41578
rect 24726 41526 27888 41578
rect 672 41492 27888 41526
rect 10098 41246 10110 41298
rect 10162 41246 10174 41298
rect 14354 41246 14366 41298
rect 14418 41246 14430 41298
rect 1038 41186 1090 41198
rect 2034 41134 2046 41186
rect 2098 41134 2110 41186
rect 10658 41134 10670 41186
rect 10722 41134 10734 41186
rect 11778 41134 11790 41186
rect 11842 41134 11854 41186
rect 24770 41134 24782 41186
rect 24834 41134 24846 41186
rect 26450 41134 26462 41186
rect 26514 41134 26526 41186
rect 1038 41122 1090 41134
rect 1598 41074 1650 41086
rect 1598 41010 1650 41022
rect 2494 41074 2546 41086
rect 25678 41074 25730 41086
rect 12114 41022 12126 41074
rect 12178 41022 12190 41074
rect 13906 41022 13918 41074
rect 13970 41022 13982 41074
rect 2494 41010 2546 41022
rect 25678 41010 25730 41022
rect 8990 40962 9042 40974
rect 8990 40898 9042 40910
rect 15486 40962 15538 40974
rect 15486 40898 15538 40910
rect 27246 40962 27298 40974
rect 27246 40898 27298 40910
rect 672 40794 27888 40828
rect 672 40742 3806 40794
rect 3858 40742 3910 40794
rect 3962 40742 4014 40794
rect 4066 40742 23806 40794
rect 23858 40742 23910 40794
rect 23962 40742 24014 40794
rect 24066 40742 27888 40794
rect 672 40708 27888 40742
rect 2494 40514 2546 40526
rect 25678 40514 25730 40526
rect 3266 40462 3278 40514
rect 3330 40462 3342 40514
rect 2494 40450 2546 40462
rect 25678 40450 25730 40462
rect 1934 40402 1986 40414
rect 1138 40350 1150 40402
rect 1202 40350 1214 40402
rect 1934 40338 1986 40350
rect 6078 40402 6130 40414
rect 6402 40350 6414 40402
rect 6466 40350 6478 40402
rect 6850 40350 6862 40402
rect 6914 40350 6926 40402
rect 8194 40350 8206 40402
rect 8258 40350 8270 40402
rect 9202 40350 9214 40402
rect 9266 40350 9278 40402
rect 10434 40350 10446 40402
rect 10498 40350 10510 40402
rect 14354 40350 14366 40402
rect 14418 40350 14430 40402
rect 26226 40350 26238 40402
rect 26290 40350 26302 40402
rect 6078 40338 6130 40350
rect 1598 40290 1650 40302
rect 1598 40226 1650 40238
rect 7534 40290 7586 40302
rect 12798 40290 12850 40302
rect 10882 40238 10894 40290
rect 10946 40238 10958 40290
rect 24658 40238 24670 40290
rect 24722 40238 24734 40290
rect 27010 40238 27022 40290
rect 27074 40238 27086 40290
rect 7534 40226 7586 40238
rect 12798 40226 12850 40238
rect 2830 40178 2882 40190
rect 12126 40178 12178 40190
rect 7074 40126 7086 40178
rect 7138 40126 7150 40178
rect 2830 40114 2882 40126
rect 12126 40114 12178 40126
rect 13358 40178 13410 40190
rect 16046 40178 16098 40190
rect 14914 40126 14926 40178
rect 14978 40126 14990 40178
rect 13358 40114 13410 40126
rect 16046 40114 16098 40126
rect 672 40010 27888 40044
rect 672 39958 4466 40010
rect 4518 39958 4570 40010
rect 4622 39958 4674 40010
rect 4726 39958 24466 40010
rect 24518 39958 24570 40010
rect 24622 39958 24674 40010
rect 24726 39958 27888 40010
rect 672 39924 27888 39958
rect 2494 39842 2546 39854
rect 2494 39778 2546 39790
rect 6974 39842 7026 39854
rect 6974 39778 7026 39790
rect 7870 39842 7922 39854
rect 7870 39778 7922 39790
rect 2158 39730 2210 39742
rect 2158 39666 2210 39678
rect 3054 39730 3106 39742
rect 3054 39666 3106 39678
rect 7310 39730 7362 39742
rect 7310 39666 7362 39678
rect 9550 39730 9602 39742
rect 9550 39666 9602 39678
rect 3950 39618 4002 39630
rect 1698 39566 1710 39618
rect 1762 39566 1774 39618
rect 3950 39554 4002 39566
rect 8990 39618 9042 39630
rect 14018 39566 14030 39618
rect 14082 39566 14094 39618
rect 24658 39566 24670 39618
rect 24722 39566 24734 39618
rect 26226 39566 26238 39618
rect 26290 39566 26302 39618
rect 8990 39554 9042 39566
rect 3490 39454 3502 39506
rect 3554 39454 3566 39506
rect 6514 39454 6526 39506
rect 6578 39454 6590 39506
rect 10546 39454 10558 39506
rect 10610 39454 10622 39506
rect 25678 39394 25730 39406
rect 25678 39330 25730 39342
rect 27246 39394 27298 39406
rect 27246 39330 27298 39342
rect 672 39226 27888 39260
rect 672 39174 3806 39226
rect 3858 39174 3910 39226
rect 3962 39174 4014 39226
rect 4066 39174 23806 39226
rect 23858 39174 23910 39226
rect 23962 39174 24014 39226
rect 24066 39174 27888 39226
rect 672 39140 27888 39174
rect 6974 39058 7026 39070
rect 6974 38994 7026 39006
rect 1598 38946 1650 38958
rect 12238 38946 12290 38958
rect 5394 38894 5406 38946
rect 5458 38894 5470 38946
rect 1598 38882 1650 38894
rect 12238 38882 12290 38894
rect 16942 38946 16994 38958
rect 16942 38882 16994 38894
rect 9438 38834 9490 38846
rect 14254 38834 14306 38846
rect 2146 38782 2158 38834
rect 2210 38782 2222 38834
rect 8306 38782 8318 38834
rect 8370 38782 8382 38834
rect 8754 38782 8766 38834
rect 8818 38782 8830 38834
rect 10098 38782 10110 38834
rect 10162 38782 10174 38834
rect 10994 38782 11006 38834
rect 11058 38782 11070 38834
rect 11778 38782 11790 38834
rect 11842 38782 11854 38834
rect 13122 38782 13134 38834
rect 13186 38782 13198 38834
rect 13570 38782 13582 38834
rect 13634 38782 13646 38834
rect 14802 38782 14814 38834
rect 14866 38782 14878 38834
rect 15810 38782 15822 38834
rect 15874 38782 15886 38834
rect 9438 38770 9490 38782
rect 14254 38770 14306 38782
rect 7982 38722 8034 38734
rect 12798 38722 12850 38734
rect 5842 38670 5854 38722
rect 5906 38670 5918 38722
rect 8978 38670 8990 38722
rect 9042 38670 9054 38722
rect 13794 38670 13806 38722
rect 13858 38670 13870 38722
rect 26226 38670 26238 38722
rect 26290 38670 26302 38722
rect 27010 38670 27022 38722
rect 27074 38670 27086 38722
rect 7982 38658 8034 38670
rect 12798 38658 12850 38670
rect 1038 38610 1090 38622
rect 3838 38610 3890 38622
rect 2706 38558 2718 38610
rect 2770 38558 2782 38610
rect 1038 38546 1090 38558
rect 3838 38546 3890 38558
rect 16382 38610 16434 38622
rect 16382 38546 16434 38558
rect 672 38442 27888 38476
rect 672 38390 4466 38442
rect 4518 38390 4570 38442
rect 4622 38390 4674 38442
rect 4726 38390 24466 38442
rect 24518 38390 24570 38442
rect 24622 38390 24674 38442
rect 24726 38390 27888 38442
rect 672 38356 27888 38390
rect 5966 38274 6018 38286
rect 5966 38210 6018 38222
rect 8206 38274 8258 38286
rect 8206 38210 8258 38222
rect 15150 38274 15202 38286
rect 15150 38210 15202 38222
rect 15710 38162 15762 38174
rect 1810 38110 1822 38162
rect 1874 38110 1886 38162
rect 4722 38110 4734 38162
rect 4786 38110 4798 38162
rect 6962 38110 6974 38162
rect 7026 38110 7038 38162
rect 15710 38098 15762 38110
rect 6626 37998 6638 38050
rect 6690 37998 6702 38050
rect 14690 37998 14702 38050
rect 14754 37998 14766 38050
rect 24882 37998 24894 38050
rect 24946 37998 24958 38050
rect 26226 37998 26238 38050
rect 26290 37998 26302 38050
rect 25678 37938 25730 37950
rect 1362 37886 1374 37938
rect 1426 37886 1438 37938
rect 4386 37886 4398 37938
rect 4450 37886 4462 37938
rect 9650 37886 9662 37938
rect 9714 37886 9726 37938
rect 26898 37886 26910 37938
rect 26962 37886 26974 37938
rect 25678 37874 25730 37886
rect 2942 37826 2994 37838
rect 2942 37762 2994 37774
rect 672 37658 27888 37692
rect 672 37606 3806 37658
rect 3858 37606 3910 37658
rect 3962 37606 4014 37658
rect 4066 37606 23806 37658
rect 23858 37606 23910 37658
rect 23962 37606 24014 37658
rect 24066 37606 27888 37658
rect 672 37572 27888 37606
rect 8094 37490 8146 37502
rect 8094 37426 8146 37438
rect 1698 37326 1710 37378
rect 1762 37326 1774 37378
rect 2706 37326 2718 37378
rect 2770 37326 2782 37378
rect 6514 37326 6526 37378
rect 6578 37326 6590 37378
rect 12002 37326 12014 37378
rect 12066 37326 12078 37378
rect 27122 37326 27134 37378
rect 27186 37326 27198 37378
rect 16606 37266 16658 37278
rect 2034 37214 2046 37266
rect 2098 37214 2110 37266
rect 8642 37214 8654 37266
rect 8706 37214 8718 37266
rect 13122 37214 13134 37266
rect 13186 37214 13198 37266
rect 15474 37214 15486 37266
rect 15538 37214 15550 37266
rect 15922 37214 15934 37266
rect 15986 37214 15998 37266
rect 17154 37214 17166 37266
rect 17218 37214 17230 37266
rect 18162 37214 18174 37266
rect 18226 37214 18238 37266
rect 16606 37202 16658 37214
rect 15150 37154 15202 37166
rect 9314 37102 9326 37154
rect 9378 37102 9390 37154
rect 13570 37102 13582 37154
rect 13634 37102 13646 37154
rect 24658 37102 24670 37154
rect 24722 37102 24734 37154
rect 25442 37102 25454 37154
rect 25506 37102 25518 37154
rect 26226 37102 26238 37154
rect 26290 37102 26302 37154
rect 15150 37090 15202 37102
rect 4286 37042 4338 37054
rect 14702 37042 14754 37054
rect 3154 36990 3166 37042
rect 3218 36990 3230 37042
rect 6962 36990 6974 37042
rect 7026 36990 7038 37042
rect 16146 36990 16158 37042
rect 16210 36990 16222 37042
rect 4286 36978 4338 36990
rect 14702 36978 14754 36990
rect 672 36874 27888 36908
rect 672 36822 4466 36874
rect 4518 36822 4570 36874
rect 4622 36822 4674 36874
rect 4726 36822 24466 36874
rect 24518 36822 24570 36874
rect 24622 36822 24674 36874
rect 24726 36822 27888 36874
rect 672 36788 27888 36822
rect 7982 36706 8034 36718
rect 10558 36706 10610 36718
rect 4162 36654 4174 36706
rect 4226 36654 4238 36706
rect 10210 36654 10222 36706
rect 10274 36654 10286 36706
rect 7982 36642 8034 36654
rect 10558 36642 10610 36654
rect 16718 36706 16770 36718
rect 16718 36642 16770 36654
rect 19854 36594 19906 36606
rect 6402 36542 6414 36594
rect 6466 36542 6478 36594
rect 18274 36542 18286 36594
rect 18338 36542 18350 36594
rect 24658 36542 24670 36594
rect 24722 36542 24734 36594
rect 19854 36530 19906 36542
rect 2606 36482 2658 36494
rect 20414 36482 20466 36494
rect 4722 36430 4734 36482
rect 4786 36430 4798 36482
rect 6850 36430 6862 36482
rect 6914 36430 6926 36482
rect 10882 36430 10894 36482
rect 10946 36430 10958 36482
rect 17714 36430 17726 36482
rect 17778 36430 17790 36482
rect 26226 36430 26238 36482
rect 26290 36430 26302 36482
rect 2606 36418 2658 36430
rect 20414 36418 20466 36430
rect 7422 36370 7474 36382
rect 17278 36370 17330 36382
rect 2146 36318 2158 36370
rect 2210 36318 2222 36370
rect 13570 36318 13582 36370
rect 13634 36318 13646 36370
rect 7422 36306 7474 36318
rect 17278 36306 17330 36318
rect 3054 36258 3106 36270
rect 3054 36194 3106 36206
rect 5294 36258 5346 36270
rect 5294 36194 5346 36206
rect 19406 36258 19458 36270
rect 19406 36194 19458 36206
rect 25678 36258 25730 36270
rect 25678 36194 25730 36206
rect 27246 36258 27298 36270
rect 27246 36194 27298 36206
rect 672 36090 27888 36124
rect 672 36038 3806 36090
rect 3858 36038 3910 36090
rect 3962 36038 4014 36090
rect 4066 36038 23806 36090
rect 23858 36038 23910 36090
rect 23962 36038 24014 36090
rect 24066 36038 27888 36090
rect 672 36004 27888 36038
rect 2706 35758 2718 35810
rect 2770 35758 2782 35810
rect 5506 35758 5518 35810
rect 5570 35758 5582 35810
rect 6514 35758 6526 35810
rect 6578 35758 6590 35810
rect 11778 35758 11790 35810
rect 11842 35758 11854 35810
rect 4398 35698 4450 35710
rect 3938 35646 3950 35698
rect 4002 35646 4014 35698
rect 8642 35646 8654 35698
rect 8706 35646 8718 35698
rect 13570 35646 13582 35698
rect 13634 35646 13646 35698
rect 4398 35634 4450 35646
rect 2258 35534 2270 35586
rect 2322 35534 2334 35586
rect 6850 35534 6862 35586
rect 6914 35534 6926 35586
rect 9314 35534 9326 35586
rect 9378 35534 9390 35586
rect 14802 35534 14814 35586
rect 14866 35534 14878 35586
rect 26226 35534 26238 35586
rect 26290 35534 26302 35586
rect 27010 35534 27022 35586
rect 27074 35534 27086 35586
rect 1150 35474 1202 35486
rect 1150 35410 1202 35422
rect 5966 35474 6018 35486
rect 5966 35410 6018 35422
rect 8094 35474 8146 35486
rect 8094 35410 8146 35422
rect 672 35306 27888 35340
rect 672 35254 4466 35306
rect 4518 35254 4570 35306
rect 4622 35254 4674 35306
rect 4726 35254 24466 35306
rect 24518 35254 24570 35306
rect 24622 35254 24674 35306
rect 24726 35254 27888 35306
rect 672 35220 27888 35254
rect 3826 35086 3838 35138
rect 3890 35086 3902 35138
rect 4286 35026 4338 35038
rect 17950 35026 18002 35038
rect 6962 34974 6974 35026
rect 7026 34974 7038 35026
rect 14018 34974 14030 35026
rect 14082 34974 14094 35026
rect 19282 34974 19294 35026
rect 19346 34974 19358 35026
rect 4286 34962 4338 34974
rect 17950 34962 18002 34974
rect 1038 34914 1090 34926
rect 1038 34850 1090 34862
rect 1934 34914 1986 34926
rect 3154 34862 3166 34914
rect 3218 34862 3230 34914
rect 3602 34862 3614 34914
rect 3666 34862 3678 34914
rect 4834 34862 4846 34914
rect 4898 34862 4910 34914
rect 5842 34862 5854 34914
rect 5906 34862 5918 34914
rect 6514 34862 6526 34914
rect 6578 34862 6590 34914
rect 9650 34862 9662 34914
rect 9714 34862 9726 34914
rect 10882 34862 10894 34914
rect 10946 34862 10958 34914
rect 17490 34862 17502 34914
rect 17554 34862 17566 34914
rect 18722 34862 18734 34914
rect 18786 34862 18798 34914
rect 19058 34862 19070 34914
rect 19122 34862 19134 34914
rect 19842 34862 19854 34914
rect 19906 34862 19918 34914
rect 20514 34862 20526 34914
rect 20578 34862 20590 34914
rect 21298 34862 21310 34914
rect 21362 34862 21374 34914
rect 24658 34862 24670 34914
rect 24722 34862 24734 34914
rect 26226 34862 26238 34914
rect 26290 34862 26302 34914
rect 1934 34850 1986 34862
rect 1598 34802 1650 34814
rect 1598 34738 1650 34750
rect 2494 34802 2546 34814
rect 2494 34738 2546 34750
rect 2830 34802 2882 34814
rect 18286 34802 18338 34814
rect 9986 34750 9998 34802
rect 10050 34750 10062 34802
rect 2830 34738 2882 34750
rect 18286 34738 18338 34750
rect 25678 34802 25730 34814
rect 25678 34738 25730 34750
rect 8206 34690 8258 34702
rect 8206 34626 8258 34638
rect 27246 34690 27298 34702
rect 27246 34626 27298 34638
rect 672 34522 27888 34556
rect 672 34470 3806 34522
rect 3858 34470 3910 34522
rect 3962 34470 4014 34522
rect 4066 34470 23806 34522
rect 23858 34470 23910 34522
rect 23962 34470 24014 34522
rect 24066 34470 27888 34522
rect 672 34436 27888 34470
rect 18958 34354 19010 34366
rect 18958 34290 19010 34302
rect 25678 34242 25730 34254
rect 27122 34190 27134 34242
rect 27186 34190 27198 34242
rect 25678 34178 25730 34190
rect 2830 34130 2882 34142
rect 10222 34130 10274 34142
rect 19518 34130 19570 34142
rect 1474 34078 1486 34130
rect 1538 34078 1550 34130
rect 1922 34078 1934 34130
rect 1986 34078 1998 34130
rect 3378 34078 3390 34130
rect 3442 34078 3454 34130
rect 4274 34078 4286 34130
rect 4338 34078 4350 34130
rect 5170 34078 5182 34130
rect 5234 34078 5246 34130
rect 8194 34078 8206 34130
rect 8258 34078 8270 34130
rect 9090 34078 9102 34130
rect 9154 34078 9166 34130
rect 9650 34078 9662 34130
rect 9714 34078 9726 34130
rect 10770 34078 10782 34130
rect 10834 34078 10846 34130
rect 10994 34078 11006 34130
rect 11058 34078 11070 34130
rect 11778 34078 11790 34130
rect 11842 34078 11854 34130
rect 12674 34078 12686 34130
rect 12738 34078 12750 34130
rect 17378 34078 17390 34130
rect 17442 34078 17454 34130
rect 24882 34078 24894 34130
rect 24946 34078 24958 34130
rect 2830 34066 2882 34078
rect 10222 34066 10274 34078
rect 19518 34066 19570 34078
rect 1150 34018 1202 34030
rect 8766 34018 8818 34030
rect 20078 34018 20130 34030
rect 2146 33966 2158 34018
rect 2210 33966 2222 34018
rect 9762 33966 9774 34018
rect 9826 33966 9838 34018
rect 13570 33966 13582 34018
rect 13634 33966 13646 34018
rect 17826 33966 17838 34018
rect 17890 33966 17902 34018
rect 26226 33966 26238 34018
rect 26290 33966 26302 34018
rect 1150 33954 1202 33966
rect 8766 33954 8818 33966
rect 20078 33954 20130 33966
rect 5518 33906 5570 33918
rect 5518 33842 5570 33854
rect 6638 33906 6690 33918
rect 7746 33854 7758 33906
rect 7810 33854 7822 33906
rect 16258 33854 16270 33906
rect 16322 33854 16334 33906
rect 6638 33842 6690 33854
rect 672 33738 27888 33772
rect 672 33686 4466 33738
rect 4518 33686 4570 33738
rect 4622 33686 4674 33738
rect 4726 33686 24466 33738
rect 24518 33686 24570 33738
rect 24622 33686 24674 33738
rect 24726 33686 27888 33738
rect 672 33652 27888 33686
rect 2270 33458 2322 33470
rect 8878 33458 8930 33470
rect 3266 33406 3278 33458
rect 3330 33406 3342 33458
rect 7634 33406 7646 33458
rect 7698 33406 7710 33458
rect 10882 33406 10894 33458
rect 10946 33406 10958 33458
rect 18722 33406 18734 33458
rect 18786 33406 18798 33458
rect 2270 33394 2322 33406
rect 8878 33394 8930 33406
rect 1038 33346 1090 33358
rect 3726 33346 3778 33358
rect 2706 33294 2718 33346
rect 2770 33294 2782 33346
rect 3042 33294 3054 33346
rect 3106 33294 3118 33346
rect 4498 33294 4510 33346
rect 4562 33294 4574 33346
rect 5282 33294 5294 33346
rect 5346 33294 5358 33346
rect 8194 33294 8206 33346
rect 8258 33294 8270 33346
rect 10322 33294 10334 33346
rect 10386 33294 10398 33346
rect 12562 33294 12574 33346
rect 12626 33294 12638 33346
rect 24882 33294 24894 33346
rect 24946 33294 24958 33346
rect 26226 33294 26238 33346
rect 26290 33294 26302 33346
rect 1038 33282 1090 33294
rect 3726 33282 3778 33294
rect 1598 33234 1650 33246
rect 1598 33170 1650 33182
rect 9438 33234 9490 33246
rect 13234 33182 13246 33234
rect 13298 33182 13310 33234
rect 15586 33182 15598 33234
rect 15650 33182 15662 33234
rect 18386 33182 18398 33234
rect 18450 33182 18462 33234
rect 9438 33170 9490 33182
rect 6526 33122 6578 33134
rect 6526 33058 6578 33070
rect 12014 33122 12066 33134
rect 12014 33058 12066 33070
rect 19966 33122 20018 33134
rect 19966 33058 20018 33070
rect 25678 33122 25730 33134
rect 25678 33058 25730 33070
rect 27246 33122 27298 33134
rect 27246 33058 27298 33070
rect 672 32954 27888 32988
rect 672 32902 3806 32954
rect 3858 32902 3910 32954
rect 3962 32902 4014 32954
rect 4066 32902 23806 32954
rect 23858 32902 23910 32954
rect 23962 32902 24014 32954
rect 24066 32902 27888 32954
rect 672 32868 27888 32902
rect 2830 32786 2882 32798
rect 2830 32722 2882 32734
rect 3838 32674 3890 32686
rect 19742 32674 19794 32686
rect 22094 32674 22146 32686
rect 15586 32622 15598 32674
rect 15650 32622 15662 32674
rect 20738 32622 20750 32674
rect 20802 32622 20814 32674
rect 3838 32610 3890 32622
rect 19742 32610 19794 32622
rect 22094 32610 22146 32622
rect 21198 32562 21250 32574
rect 1138 32510 1150 32562
rect 1202 32510 1214 32562
rect 3378 32510 3390 32562
rect 3442 32510 3454 32562
rect 5058 32510 5070 32562
rect 5122 32510 5134 32562
rect 7186 32510 7198 32562
rect 7250 32510 7262 32562
rect 9874 32510 9886 32562
rect 9938 32510 9950 32562
rect 14802 32510 14814 32562
rect 14866 32510 14878 32562
rect 19282 32510 19294 32562
rect 19346 32510 19358 32562
rect 26450 32510 26462 32562
rect 26514 32510 26526 32562
rect 21198 32498 21250 32510
rect 1698 32398 1710 32450
rect 1762 32398 1774 32450
rect 4946 32398 4958 32450
rect 5010 32398 5022 32450
rect 7634 32398 7646 32450
rect 7698 32398 7710 32450
rect 27010 32398 27022 32450
rect 27074 32398 27086 32450
rect 5518 32338 5570 32350
rect 5518 32274 5570 32286
rect 8878 32338 8930 32350
rect 11454 32338 11506 32350
rect 10322 32286 10334 32338
rect 10386 32286 10398 32338
rect 8878 32274 8930 32286
rect 11454 32274 11506 32286
rect 21534 32338 21586 32350
rect 21534 32274 21586 32286
rect 672 32170 27888 32204
rect 672 32118 4466 32170
rect 4518 32118 4570 32170
rect 4622 32118 4674 32170
rect 4726 32118 24466 32170
rect 24518 32118 24570 32170
rect 24622 32118 24674 32170
rect 24726 32118 27888 32170
rect 672 32084 27888 32118
rect 21186 31950 21198 32002
rect 21250 31950 21262 32002
rect 9662 31890 9714 31902
rect 2034 31838 2046 31890
rect 2098 31838 2110 31890
rect 6066 31838 6078 31890
rect 6130 31838 6142 31890
rect 9662 31826 9714 31838
rect 11118 31890 11170 31902
rect 12910 31890 12962 31902
rect 12450 31838 12462 31890
rect 12514 31838 12526 31890
rect 11118 31826 11170 31838
rect 12910 31826 12962 31838
rect 17278 31890 17330 31902
rect 18498 31838 18510 31890
rect 18562 31838 18574 31890
rect 17278 31826 17330 31838
rect 3278 31778 3330 31790
rect 6526 31778 6578 31790
rect 10222 31778 10274 31790
rect 16718 31778 16770 31790
rect 1698 31726 1710 31778
rect 1762 31726 1774 31778
rect 5394 31726 5406 31778
rect 5458 31726 5470 31778
rect 5954 31726 5966 31778
rect 6018 31726 6030 31778
rect 7298 31726 7310 31778
rect 7362 31726 7374 31778
rect 8082 31726 8094 31778
rect 8146 31726 8158 31778
rect 11778 31726 11790 31778
rect 11842 31726 11854 31778
rect 12226 31726 12238 31778
rect 12290 31726 12302 31778
rect 13458 31726 13470 31778
rect 13522 31726 13534 31778
rect 14466 31726 14478 31778
rect 14530 31726 14542 31778
rect 18050 31726 18062 31778
rect 18114 31726 18126 31778
rect 20626 31726 20638 31778
rect 20690 31726 20702 31778
rect 20962 31726 20974 31778
rect 21026 31726 21038 31778
rect 21746 31726 21758 31778
rect 21810 31726 21822 31778
rect 22418 31726 22430 31778
rect 22482 31726 22494 31778
rect 23202 31726 23214 31778
rect 23266 31726 23278 31778
rect 24658 31726 24670 31778
rect 24722 31726 24734 31778
rect 26450 31726 26462 31778
rect 26514 31726 26526 31778
rect 3278 31714 3330 31726
rect 6526 31714 6578 31726
rect 10222 31714 10274 31726
rect 16718 31714 16770 31726
rect 5070 31666 5122 31678
rect 11454 31666 11506 31678
rect 10658 31614 10670 31666
rect 10722 31614 10734 31666
rect 5070 31602 5122 31614
rect 11454 31602 11506 31614
rect 20190 31666 20242 31678
rect 20190 31602 20242 31614
rect 25678 31666 25730 31678
rect 27122 31614 27134 31666
rect 27186 31614 27198 31666
rect 25678 31602 25730 31614
rect 19742 31554 19794 31566
rect 19742 31490 19794 31502
rect 672 31386 27888 31420
rect 672 31334 3806 31386
rect 3858 31334 3910 31386
rect 3962 31334 4014 31386
rect 4066 31334 23806 31386
rect 23858 31334 23910 31386
rect 23962 31334 24014 31386
rect 24066 31334 27888 31386
rect 672 31300 27888 31334
rect 4286 31218 4338 31230
rect 4286 31154 4338 31166
rect 1598 31106 1650 31118
rect 5518 31106 5570 31118
rect 2706 31054 2718 31106
rect 2770 31054 2782 31106
rect 1598 31042 1650 31054
rect 5518 31042 5570 31054
rect 6414 31106 6466 31118
rect 6414 31042 6466 31054
rect 12238 31106 12290 31118
rect 12238 31042 12290 31054
rect 10558 30994 10610 31006
rect 22094 30994 22146 31006
rect 5058 30942 5070 30994
rect 5122 30942 5134 30994
rect 5954 30942 5966 30994
rect 6018 30942 6030 30994
rect 6962 30942 6974 30994
rect 7026 30942 7038 30994
rect 9090 30942 9102 30994
rect 9154 30942 9166 30994
rect 9986 30942 9998 30994
rect 10050 30942 10062 30994
rect 11330 30942 11342 30994
rect 11394 30942 11406 30994
rect 11778 30942 11790 30994
rect 11842 30942 11854 30994
rect 13458 30942 13470 30994
rect 13522 30942 13534 30994
rect 15810 30942 15822 30994
rect 15874 30942 15886 30994
rect 16258 30942 16270 30994
rect 16322 30942 16334 30994
rect 17714 30942 17726 30994
rect 17778 30942 17790 30994
rect 18498 30942 18510 30994
rect 18562 30942 18574 30994
rect 20962 30942 20974 30994
rect 21026 30942 21038 30994
rect 21522 30942 21534 30994
rect 21586 30942 21598 30994
rect 22642 30942 22654 30994
rect 22706 30942 22718 30994
rect 23650 30942 23662 30994
rect 23714 30942 23726 30994
rect 24770 30942 24782 30994
rect 24834 30942 24846 30994
rect 10558 30930 10610 30942
rect 22094 30930 22146 30942
rect 15038 30882 15090 30894
rect 7298 30830 7310 30882
rect 7362 30830 7374 30882
rect 11218 30830 11230 30882
rect 11282 30830 11294 30882
rect 15038 30818 15090 30830
rect 15486 30882 15538 30894
rect 16942 30882 16994 30894
rect 16482 30830 16494 30882
rect 16546 30830 16558 30882
rect 15486 30818 15538 30830
rect 16942 30818 16994 30830
rect 20638 30882 20690 30894
rect 21634 30830 21646 30882
rect 21698 30830 21710 30882
rect 25442 30830 25454 30882
rect 25506 30830 25518 30882
rect 26226 30830 26238 30882
rect 26290 30830 26302 30882
rect 27010 30830 27022 30882
rect 27074 30830 27086 30882
rect 20638 30818 20690 30830
rect 1038 30770 1090 30782
rect 8542 30770 8594 30782
rect 3154 30718 3166 30770
rect 3218 30718 3230 30770
rect 13906 30718 13918 30770
rect 13970 30718 13982 30770
rect 1038 30706 1090 30718
rect 8542 30706 8594 30718
rect 672 30602 27888 30636
rect 672 30550 4466 30602
rect 4518 30550 4570 30602
rect 4622 30550 4674 30602
rect 4726 30550 24466 30602
rect 24518 30550 24570 30602
rect 24622 30550 24674 30602
rect 24726 30550 27888 30602
rect 672 30516 27888 30550
rect 20862 30434 20914 30446
rect 17490 30382 17502 30434
rect 17554 30382 17566 30434
rect 19730 30382 19742 30434
rect 19794 30382 19806 30434
rect 20862 30370 20914 30382
rect 4498 30270 4510 30322
rect 4562 30270 4574 30322
rect 10882 30270 10894 30322
rect 10946 30270 10958 30322
rect 13570 30270 13582 30322
rect 13634 30270 13646 30322
rect 21858 30270 21870 30322
rect 21922 30270 21934 30322
rect 2606 30210 2658 30222
rect 4958 30210 5010 30222
rect 8878 30210 8930 30222
rect 2258 30158 2270 30210
rect 2322 30158 2334 30210
rect 3826 30158 3838 30210
rect 3890 30158 3902 30210
rect 4274 30158 4286 30210
rect 4338 30158 4350 30210
rect 5506 30158 5518 30210
rect 5570 30158 5582 30210
rect 6514 30158 6526 30210
rect 6578 30158 6590 30210
rect 7298 30158 7310 30210
rect 7362 30158 7374 30210
rect 2606 30146 2658 30158
rect 4958 30146 5010 30158
rect 8878 30146 8930 30158
rect 12126 30210 12178 30222
rect 12126 30146 12178 30158
rect 12574 30210 12626 30222
rect 14030 30210 14082 30222
rect 23102 30210 23154 30222
rect 12898 30158 12910 30210
rect 12962 30158 12974 30210
rect 13346 30158 13358 30210
rect 13410 30158 13422 30210
rect 14578 30158 14590 30210
rect 14642 30158 14654 30210
rect 15698 30158 15710 30210
rect 15762 30158 15774 30210
rect 17042 30158 17054 30210
rect 17106 30158 17118 30210
rect 19282 30158 19294 30210
rect 19346 30158 19358 30210
rect 21410 30158 21422 30210
rect 21474 30158 21486 30210
rect 26226 30158 26238 30210
rect 26290 30158 26302 30210
rect 12574 30146 12626 30158
rect 14030 30146 14082 30158
rect 23102 30146 23154 30158
rect 3502 30098 3554 30110
rect 1474 30046 1486 30098
rect 1538 30046 1550 30098
rect 3042 30046 3054 30098
rect 3106 30046 3118 30098
rect 3502 30034 3554 30046
rect 9438 30098 9490 30110
rect 10546 30046 10558 30098
rect 10610 30046 10622 30098
rect 27122 30046 27134 30098
rect 27186 30046 27198 30098
rect 9438 30034 9490 30046
rect 8094 29986 8146 29998
rect 8094 29922 8146 29934
rect 18622 29986 18674 29998
rect 18622 29922 18674 29934
rect 672 29818 27888 29852
rect 672 29766 3806 29818
rect 3858 29766 3910 29818
rect 3962 29766 4014 29818
rect 4066 29766 23806 29818
rect 23858 29766 23910 29818
rect 23962 29766 24014 29818
rect 24066 29766 27888 29818
rect 672 29732 27888 29766
rect 4286 29650 4338 29662
rect 4286 29586 4338 29598
rect 7198 29650 7250 29662
rect 7198 29586 7250 29598
rect 10110 29650 10162 29662
rect 10110 29586 10162 29598
rect 1598 29538 1650 29550
rect 14030 29538 14082 29550
rect 8530 29486 8542 29538
rect 8594 29486 8606 29538
rect 1598 29474 1650 29486
rect 14030 29474 14082 29486
rect 16046 29426 16098 29438
rect 2594 29374 2606 29426
rect 2658 29374 2670 29426
rect 5618 29374 5630 29426
rect 5682 29374 5694 29426
rect 13570 29374 13582 29426
rect 13634 29374 13646 29426
rect 14690 29374 14702 29426
rect 14754 29374 14766 29426
rect 15138 29374 15150 29426
rect 15202 29374 15214 29426
rect 16370 29374 16382 29426
rect 16434 29374 16446 29426
rect 17490 29374 17502 29426
rect 17554 29374 17566 29426
rect 18050 29374 18062 29426
rect 18114 29374 18126 29426
rect 26226 29374 26238 29426
rect 26290 29374 26302 29426
rect 16046 29362 16098 29374
rect 11678 29314 11730 29326
rect 3154 29262 3166 29314
rect 3218 29262 3230 29314
rect 5954 29262 5966 29314
rect 6018 29262 6030 29314
rect 11678 29250 11730 29262
rect 14366 29314 14418 29326
rect 18498 29262 18510 29314
rect 18562 29262 18574 29314
rect 27010 29262 27022 29314
rect 27074 29262 27086 29314
rect 14366 29250 14418 29262
rect 1038 29202 1090 29214
rect 12238 29202 12290 29214
rect 19742 29202 19794 29214
rect 8978 29150 8990 29202
rect 9042 29150 9054 29202
rect 15362 29150 15374 29202
rect 15426 29150 15438 29202
rect 1038 29138 1090 29150
rect 12238 29138 12290 29150
rect 19742 29138 19794 29150
rect 672 29034 27888 29068
rect 672 28982 4466 29034
rect 4518 28982 4570 29034
rect 4622 28982 4674 29034
rect 4726 28982 24466 29034
rect 24518 28982 24570 29034
rect 24622 28982 24674 29034
rect 24726 28982 27888 29034
rect 672 28948 27888 28982
rect 3614 28866 3666 28878
rect 15486 28866 15538 28878
rect 12562 28814 12574 28866
rect 12626 28814 12638 28866
rect 17826 28814 17838 28866
rect 17890 28814 17902 28866
rect 3614 28802 3666 28814
rect 15486 28802 15538 28814
rect 11566 28754 11618 28766
rect 2370 28702 2382 28754
rect 2434 28702 2446 28754
rect 9874 28702 9886 28754
rect 9938 28702 9950 28754
rect 20402 28702 20414 28754
rect 20466 28702 20478 28754
rect 11566 28690 11618 28702
rect 5630 28642 5682 28654
rect 4162 28590 4174 28642
rect 4226 28590 4238 28642
rect 5630 28578 5682 28590
rect 6190 28642 6242 28654
rect 11118 28642 11170 28654
rect 13022 28642 13074 28654
rect 16046 28642 16098 28654
rect 21086 28642 21138 28654
rect 7298 28590 7310 28642
rect 7362 28590 7374 28642
rect 11890 28590 11902 28642
rect 11954 28590 11966 28642
rect 12338 28590 12350 28642
rect 12402 28590 12414 28642
rect 13570 28590 13582 28642
rect 13634 28590 13646 28642
rect 14690 28590 14702 28642
rect 14754 28590 14766 28642
rect 19842 28590 19854 28642
rect 19906 28590 19918 28642
rect 20290 28590 20302 28642
rect 20354 28590 20366 28642
rect 21410 28590 21422 28642
rect 21474 28590 21486 28642
rect 21634 28590 21646 28642
rect 21698 28590 21710 28642
rect 22418 28590 22430 28642
rect 22482 28590 22494 28642
rect 26226 28590 26238 28642
rect 26290 28590 26302 28642
rect 6190 28578 6242 28590
rect 11118 28578 11170 28590
rect 13022 28578 13074 28590
rect 16046 28578 16098 28590
rect 21086 28578 21138 28590
rect 19406 28530 19458 28542
rect 2034 28478 2046 28530
rect 2098 28478 2110 28530
rect 4946 28478 4958 28530
rect 5010 28478 5022 28530
rect 7970 28478 7982 28530
rect 8034 28478 8046 28530
rect 9538 28478 9550 28530
rect 9602 28478 9614 28530
rect 17378 28478 17390 28530
rect 17442 28478 17454 28530
rect 27122 28478 27134 28530
rect 27186 28478 27198 28530
rect 19406 28466 19458 28478
rect 18958 28418 19010 28430
rect 18958 28354 19010 28366
rect 672 28250 27888 28284
rect 672 28198 3806 28250
rect 3858 28198 3910 28250
rect 3962 28198 4014 28250
rect 4066 28198 23806 28250
rect 23858 28198 23910 28250
rect 23962 28198 24014 28250
rect 24066 28198 27888 28250
rect 672 28164 27888 28198
rect 7422 28082 7474 28094
rect 7422 28018 7474 28030
rect 12126 28082 12178 28094
rect 12126 28018 12178 28030
rect 1038 27970 1090 27982
rect 1038 27906 1090 27918
rect 13582 27970 13634 27982
rect 13582 27906 13634 27918
rect 21198 27970 21250 27982
rect 21198 27906 21250 27918
rect 25678 27970 25730 27982
rect 27122 27918 27134 27970
rect 27186 27918 27198 27970
rect 25678 27906 25730 27918
rect 15262 27858 15314 27870
rect 20638 27858 20690 27870
rect 1474 27806 1486 27858
rect 1538 27806 1550 27858
rect 2258 27806 2270 27858
rect 2322 27806 2334 27858
rect 6514 27806 6526 27858
rect 6578 27806 6590 27858
rect 8082 27806 8094 27858
rect 8146 27806 8158 27858
rect 10434 27806 10446 27858
rect 10498 27806 10510 27858
rect 13906 27806 13918 27858
rect 13970 27806 13982 27858
rect 14354 27806 14366 27858
rect 14418 27806 14430 27858
rect 15810 27806 15822 27858
rect 15874 27806 15886 27858
rect 16594 27806 16606 27858
rect 16658 27806 16670 27858
rect 18050 27806 18062 27858
rect 18114 27806 18126 27858
rect 24882 27806 24894 27858
rect 24946 27806 24958 27858
rect 15262 27794 15314 27806
rect 20638 27794 20690 27806
rect 5518 27746 5570 27758
rect 2706 27694 2718 27746
rect 2770 27694 2782 27746
rect 8642 27694 8654 27746
rect 8706 27694 8718 27746
rect 10994 27694 11006 27746
rect 11058 27694 11070 27746
rect 18498 27694 18510 27746
rect 18562 27694 18574 27746
rect 26226 27694 26238 27746
rect 26290 27694 26302 27746
rect 5518 27682 5570 27694
rect 3950 27634 4002 27646
rect 3950 27570 4002 27582
rect 4958 27634 5010 27646
rect 4958 27570 5010 27582
rect 9774 27634 9826 27646
rect 19742 27634 19794 27646
rect 14578 27582 14590 27634
rect 14642 27582 14654 27634
rect 9774 27570 9826 27582
rect 19742 27570 19794 27582
rect 672 27466 27888 27500
rect 672 27414 4466 27466
rect 4518 27414 4570 27466
rect 4622 27414 4674 27466
rect 4726 27414 24466 27466
rect 24518 27414 24570 27466
rect 24622 27414 24674 27466
rect 24726 27414 27888 27466
rect 672 27380 27888 27414
rect 13134 27298 13186 27310
rect 1698 27246 1710 27298
rect 1762 27246 1774 27298
rect 4274 27246 4286 27298
rect 4338 27246 4350 27298
rect 10098 27246 10110 27298
rect 10162 27246 10174 27298
rect 12002 27246 12014 27298
rect 12066 27246 12078 27298
rect 13134 27234 13186 27246
rect 15374 27298 15426 27310
rect 15374 27234 15426 27246
rect 8318 27186 8370 27198
rect 17390 27186 17442 27198
rect 14130 27134 14142 27186
rect 14194 27134 14206 27186
rect 18386 27134 18398 27186
rect 18450 27134 18462 27186
rect 27010 27134 27022 27186
rect 27074 27134 27086 27186
rect 8318 27122 8370 27134
rect 17390 27122 17442 27134
rect 4734 27074 4786 27086
rect 1250 27022 1262 27074
rect 1314 27022 1326 27074
rect 3602 27022 3614 27074
rect 3666 27022 3678 27074
rect 4050 27022 4062 27074
rect 4114 27022 4126 27074
rect 5282 27022 5294 27074
rect 5346 27022 5358 27074
rect 6290 27022 6302 27074
rect 6354 27022 6366 27074
rect 7858 27022 7870 27074
rect 7922 27022 7934 27074
rect 13794 27022 13806 27074
rect 13858 27022 13870 27074
rect 17714 27022 17726 27074
rect 17778 27022 17790 27074
rect 18162 27022 18174 27074
rect 18226 27022 18238 27074
rect 18946 27022 18958 27074
rect 19010 27022 19022 27074
rect 19394 27022 19406 27074
rect 19458 27022 19470 27074
rect 20514 27022 20526 27074
rect 20578 27022 20590 27074
rect 24658 27022 24670 27074
rect 24722 27022 24734 27074
rect 26226 27022 26238 27074
rect 26290 27022 26302 27074
rect 4734 27010 4786 27022
rect 3278 26962 3330 26974
rect 10546 26910 10558 26962
rect 10610 26910 10622 26962
rect 11554 26910 11566 26962
rect 11618 26910 11630 26962
rect 3278 26898 3330 26910
rect 2830 26850 2882 26862
rect 2830 26786 2882 26798
rect 8990 26850 9042 26862
rect 8990 26786 9042 26798
rect 25678 26850 25730 26862
rect 25678 26786 25730 26798
rect 672 26682 27888 26716
rect 672 26630 3806 26682
rect 3858 26630 3910 26682
rect 3962 26630 4014 26682
rect 4066 26630 23806 26682
rect 23858 26630 23910 26682
rect 23962 26630 24014 26682
rect 24066 26630 27888 26682
rect 672 26596 27888 26630
rect 3614 26514 3666 26526
rect 3614 26450 3666 26462
rect 19966 26514 20018 26526
rect 19966 26450 20018 26462
rect 27246 26514 27298 26526
rect 27246 26450 27298 26462
rect 5518 26402 5570 26414
rect 2034 26350 2046 26402
rect 2098 26350 2110 26402
rect 6402 26350 6414 26402
rect 6466 26350 6478 26402
rect 17714 26350 17726 26402
rect 17778 26350 17790 26402
rect 18386 26350 18398 26402
rect 18450 26350 18462 26402
rect 5518 26338 5570 26350
rect 10670 26290 10722 26302
rect 15262 26290 15314 26302
rect 9314 26238 9326 26290
rect 9378 26238 9390 26290
rect 9874 26238 9886 26290
rect 9938 26238 9950 26290
rect 11106 26238 11118 26290
rect 11170 26238 11182 26290
rect 12002 26238 12014 26290
rect 12066 26238 12078 26290
rect 13234 26238 13246 26290
rect 13298 26238 13310 26290
rect 20738 26238 20750 26290
rect 20802 26238 20814 26290
rect 10670 26226 10722 26238
rect 15262 26226 15314 26238
rect 8990 26178 9042 26190
rect 15822 26178 15874 26190
rect 2482 26126 2494 26178
rect 2546 26126 2558 26178
rect 6738 26126 6750 26178
rect 6802 26126 6814 26178
rect 13682 26126 13694 26178
rect 13746 26126 13758 26178
rect 18722 26126 18734 26178
rect 18786 26126 18798 26178
rect 26226 26126 26238 26178
rect 26290 26126 26302 26178
rect 8990 26114 9042 26126
rect 15822 26114 15874 26126
rect 4958 26066 5010 26078
rect 4958 26002 5010 26014
rect 7982 26066 8034 26078
rect 14814 26066 14866 26078
rect 9986 26014 9998 26066
rect 10050 26014 10062 26066
rect 7982 26002 8034 26014
rect 14814 26002 14866 26014
rect 17278 26066 17330 26078
rect 22430 26066 22482 26078
rect 21298 26014 21310 26066
rect 21362 26014 21374 26066
rect 17278 26002 17330 26014
rect 22430 26002 22482 26014
rect 672 25898 27888 25932
rect 672 25846 4466 25898
rect 4518 25846 4570 25898
rect 4622 25846 4674 25898
rect 4726 25846 24466 25898
rect 24518 25846 24570 25898
rect 24622 25846 24674 25898
rect 24726 25846 27888 25898
rect 672 25812 27888 25846
rect 10670 25730 10722 25742
rect 18622 25730 18674 25742
rect 3602 25678 3614 25730
rect 3666 25678 3678 25730
rect 9538 25678 9550 25730
rect 9602 25678 9614 25730
rect 14914 25678 14926 25730
rect 14978 25678 14990 25730
rect 10670 25666 10722 25678
rect 18622 25666 18674 25678
rect 21310 25730 21362 25742
rect 21310 25666 21362 25678
rect 19182 25618 19234 25630
rect 22318 25618 22370 25630
rect 7074 25566 7086 25618
rect 7138 25566 7150 25618
rect 11666 25566 11678 25618
rect 11730 25566 11742 25618
rect 20066 25566 20078 25618
rect 20130 25566 20142 25618
rect 26226 25566 26238 25618
rect 26290 25566 26302 25618
rect 19182 25554 19234 25566
rect 22318 25554 22370 25566
rect 4062 25506 4114 25518
rect 17278 25506 17330 25518
rect 2146 25454 2158 25506
rect 2210 25454 2222 25506
rect 2930 25454 2942 25506
rect 2994 25454 3006 25506
rect 3378 25454 3390 25506
rect 3442 25454 3454 25506
rect 4610 25454 4622 25506
rect 4674 25454 4686 25506
rect 5730 25454 5742 25506
rect 5794 25454 5806 25506
rect 6514 25454 6526 25506
rect 6578 25454 6590 25506
rect 8978 25454 8990 25506
rect 9042 25454 9054 25506
rect 11330 25454 11342 25506
rect 11394 25454 11406 25506
rect 16818 25454 16830 25506
rect 16882 25454 16894 25506
rect 4062 25442 4114 25454
rect 17278 25442 17330 25454
rect 21758 25506 21810 25518
rect 24658 25454 24670 25506
rect 24722 25454 24734 25506
rect 21758 25442 21810 25454
rect 1262 25394 1314 25406
rect 1262 25330 1314 25342
rect 2606 25394 2658 25406
rect 27246 25394 27298 25406
rect 14466 25342 14478 25394
rect 14530 25342 14542 25394
rect 19730 25342 19742 25394
rect 19794 25342 19806 25394
rect 2606 25330 2658 25342
rect 27246 25330 27298 25342
rect 8206 25282 8258 25294
rect 8206 25218 8258 25230
rect 12910 25282 12962 25294
rect 12910 25218 12962 25230
rect 16046 25282 16098 25294
rect 16046 25218 16098 25230
rect 25678 25282 25730 25294
rect 25678 25218 25730 25230
rect 672 25114 27888 25148
rect 672 25062 3806 25114
rect 3858 25062 3910 25114
rect 3962 25062 4014 25114
rect 4066 25062 23806 25114
rect 23858 25062 23910 25114
rect 23962 25062 24014 25114
rect 24066 25062 27888 25114
rect 672 25028 27888 25062
rect 3502 24946 3554 24958
rect 3502 24882 3554 24894
rect 5518 24946 5570 24958
rect 5518 24882 5570 24894
rect 11118 24834 11170 24846
rect 11118 24770 11170 24782
rect 18734 24834 18786 24846
rect 18734 24770 18786 24782
rect 20638 24834 20690 24846
rect 25554 24782 25566 24834
rect 25618 24782 25630 24834
rect 27122 24782 27134 24834
rect 27186 24782 27198 24834
rect 20638 24770 20690 24782
rect 8430 24722 8482 24734
rect 10558 24722 10610 24734
rect 16046 24722 16098 24734
rect 1810 24670 1822 24722
rect 1874 24670 1886 24722
rect 5058 24670 5070 24722
rect 5122 24670 5134 24722
rect 7410 24670 7422 24722
rect 7474 24670 7486 24722
rect 7746 24670 7758 24722
rect 7810 24670 7822 24722
rect 9202 24670 9214 24722
rect 9266 24670 9278 24722
rect 9986 24670 9998 24722
rect 10050 24670 10062 24722
rect 14914 24670 14926 24722
rect 14978 24670 14990 24722
rect 15362 24670 15374 24722
rect 15426 24670 15438 24722
rect 16594 24670 16606 24722
rect 16658 24670 16670 24722
rect 17502 24717 17554 24729
rect 22318 24722 22370 24734
rect 8430 24658 8482 24670
rect 10558 24658 10610 24670
rect 16046 24658 16098 24670
rect 21074 24670 21086 24722
rect 21138 24670 21150 24722
rect 21410 24670 21422 24722
rect 21474 24670 21486 24722
rect 22642 24670 22654 24722
rect 22706 24670 22718 24722
rect 23650 24670 23662 24722
rect 23714 24670 23726 24722
rect 24882 24670 24894 24722
rect 24946 24670 24958 24722
rect 26226 24670 26238 24722
rect 26290 24670 26302 24722
rect 17502 24653 17554 24665
rect 22318 24658 22370 24670
rect 6974 24610 7026 24622
rect 13358 24610 13410 24622
rect 2370 24558 2382 24610
rect 2434 24558 2446 24610
rect 7970 24558 7982 24610
rect 8034 24558 8046 24610
rect 6974 24546 7026 24558
rect 13358 24546 13410 24558
rect 14590 24610 14642 24622
rect 21634 24558 21646 24610
rect 21698 24558 21710 24610
rect 14590 24546 14642 24558
rect 12798 24498 12850 24510
rect 18174 24498 18226 24510
rect 15586 24446 15598 24498
rect 15650 24446 15662 24498
rect 12798 24434 12850 24446
rect 18174 24434 18226 24446
rect 672 24330 27888 24364
rect 672 24278 4466 24330
rect 4518 24278 4570 24330
rect 4622 24278 4674 24330
rect 4726 24278 24466 24330
rect 24518 24278 24570 24330
rect 24622 24278 24674 24330
rect 24726 24278 27888 24330
rect 672 24244 27888 24278
rect 1038 24162 1090 24174
rect 22094 24162 22146 24174
rect 12226 24110 12238 24162
rect 12290 24110 12302 24162
rect 17714 24110 17726 24162
rect 17778 24110 17790 24162
rect 1038 24098 1090 24110
rect 22094 24098 22146 24110
rect 1598 24050 1650 24062
rect 10334 24050 10386 24062
rect 3378 23998 3390 24050
rect 3442 23998 3454 24050
rect 6514 23998 6526 24050
rect 6578 23998 6590 24050
rect 1598 23986 1650 23998
rect 10334 23986 10386 23998
rect 16046 24050 16098 24062
rect 22542 24050 22594 24062
rect 20962 23998 20974 24050
rect 21026 23998 21038 24050
rect 16046 23986 16098 23998
rect 22542 23986 22594 23998
rect 23102 24050 23154 24062
rect 24658 23998 24670 24050
rect 24722 23998 24734 24050
rect 23102 23986 23154 23998
rect 2382 23938 2434 23950
rect 4062 23938 4114 23950
rect 10894 23938 10946 23950
rect 12910 23938 12962 23950
rect 15486 23938 15538 23950
rect 18174 23938 18226 23950
rect 2818 23886 2830 23938
rect 2882 23886 2894 23938
rect 3154 23886 3166 23938
rect 3218 23886 3230 23938
rect 4610 23886 4622 23938
rect 4674 23886 4686 23938
rect 5506 23886 5518 23938
rect 5570 23886 5582 23938
rect 6066 23886 6078 23938
rect 6130 23886 6142 23938
rect 11554 23886 11566 23938
rect 11618 23886 11630 23938
rect 12002 23886 12014 23938
rect 12066 23886 12078 23938
rect 13458 23886 13470 23938
rect 13522 23886 13534 23938
rect 14354 23886 14366 23938
rect 14418 23886 14430 23938
rect 17042 23886 17054 23938
rect 17106 23886 17118 23938
rect 17490 23886 17502 23938
rect 17554 23886 17566 23938
rect 18722 23886 18734 23938
rect 18786 23886 18798 23938
rect 18946 23886 18958 23938
rect 19010 23886 19022 23938
rect 19842 23886 19854 23938
rect 19906 23886 19918 23938
rect 20514 23886 20526 23938
rect 20578 23886 20590 23938
rect 26226 23886 26238 23938
rect 26290 23886 26302 23938
rect 2382 23874 2434 23886
rect 4062 23874 4114 23886
rect 10894 23874 10946 23886
rect 12910 23874 12962 23886
rect 15486 23874 15538 23886
rect 18174 23874 18226 23886
rect 11230 23826 11282 23838
rect 6178 23774 6190 23826
rect 6242 23774 6254 23826
rect 11230 23762 11282 23774
rect 16718 23826 16770 23838
rect 16718 23762 16770 23774
rect 27246 23826 27298 23838
rect 27246 23762 27298 23774
rect 7758 23714 7810 23726
rect 7758 23650 7810 23662
rect 25678 23714 25730 23726
rect 25678 23650 25730 23662
rect 672 23546 27888 23580
rect 672 23494 3806 23546
rect 3858 23494 3910 23546
rect 3962 23494 4014 23546
rect 4066 23494 23806 23546
rect 23858 23494 23910 23546
rect 23962 23494 24014 23546
rect 24066 23494 27888 23546
rect 672 23460 27888 23494
rect 3838 23378 3890 23390
rect 3838 23314 3890 23326
rect 16270 23378 16322 23390
rect 16270 23314 16322 23326
rect 13246 23266 13298 23278
rect 2258 23214 2270 23266
rect 2322 23214 2334 23266
rect 5282 23214 5294 23266
rect 5346 23214 5358 23266
rect 27122 23214 27134 23266
rect 27186 23214 27198 23266
rect 13246 23202 13298 23214
rect 19966 23154 20018 23166
rect 1586 23102 1598 23154
rect 1650 23102 1662 23154
rect 6290 23102 6302 23154
rect 6354 23102 6366 23154
rect 9314 23102 9326 23154
rect 9378 23102 9390 23154
rect 10322 23102 10334 23154
rect 10386 23102 10398 23154
rect 14690 23102 14702 23154
rect 14754 23102 14766 23154
rect 19966 23090 20018 23102
rect 1150 23042 1202 23054
rect 19630 23042 19682 23054
rect 2706 22990 2718 23042
rect 2770 22990 2782 23042
rect 6850 22990 6862 23042
rect 6914 22990 6926 23042
rect 8866 22990 8878 23042
rect 8930 22990 8942 23042
rect 15138 22990 15150 23042
rect 15202 22990 15214 23042
rect 26226 22990 26238 23042
rect 26290 22990 26302 23042
rect 1150 22978 1202 22990
rect 19630 22978 19682 22990
rect 5742 22930 5794 22942
rect 5742 22866 5794 22878
rect 7758 22930 7810 22942
rect 12014 22930 12066 22942
rect 10882 22878 10894 22930
rect 10946 22878 10958 22930
rect 7758 22866 7810 22878
rect 12014 22866 12066 22878
rect 13806 22930 13858 22942
rect 13806 22866 13858 22878
rect 19854 22930 19906 22942
rect 19854 22866 19906 22878
rect 20078 22930 20130 22942
rect 20078 22866 20130 22878
rect 672 22762 27888 22796
rect 672 22710 4466 22762
rect 4518 22710 4570 22762
rect 4622 22710 4674 22762
rect 4726 22710 24466 22762
rect 24518 22710 24570 22762
rect 24622 22710 24674 22762
rect 24726 22710 27888 22762
rect 672 22676 27888 22710
rect 2830 22594 2882 22606
rect 13358 22594 13410 22606
rect 12226 22542 12238 22594
rect 12290 22542 12302 22594
rect 2830 22530 2882 22542
rect 13358 22530 13410 22542
rect 23438 22482 23490 22494
rect 1586 22430 1598 22482
rect 1650 22430 1662 22482
rect 6066 22430 6078 22482
rect 6130 22430 6142 22482
rect 9986 22430 9998 22482
rect 10050 22430 10062 22482
rect 14802 22430 14814 22482
rect 14866 22430 14878 22482
rect 17938 22430 17950 22482
rect 18002 22430 18014 22482
rect 20290 22430 20302 22482
rect 20354 22430 20366 22482
rect 26226 22430 26238 22482
rect 26290 22430 26302 22482
rect 23438 22418 23490 22430
rect 20750 22370 20802 22382
rect 22878 22370 22930 22382
rect 4274 22318 4286 22370
rect 4338 22318 4350 22370
rect 9538 22318 9550 22370
rect 9602 22318 9614 22370
rect 14354 22318 14366 22370
rect 14418 22318 14430 22370
rect 18386 22318 18398 22370
rect 18450 22318 18462 22370
rect 19618 22318 19630 22370
rect 19682 22318 19694 22370
rect 20066 22318 20078 22370
rect 20130 22318 20142 22370
rect 21298 22318 21310 22370
rect 21362 22318 21374 22370
rect 22418 22318 22430 22370
rect 22482 22318 22494 22370
rect 24882 22318 24894 22370
rect 24946 22318 24958 22370
rect 20750 22306 20802 22318
rect 22878 22306 22930 22318
rect 3502 22258 3554 22270
rect 19294 22258 19346 22270
rect 1250 22206 1262 22258
rect 1314 22206 1326 22258
rect 5618 22206 5630 22258
rect 5682 22206 5694 22258
rect 11778 22206 11790 22258
rect 11842 22206 11854 22258
rect 3502 22194 3554 22206
rect 19294 22194 19346 22206
rect 27246 22258 27298 22270
rect 27246 22194 27298 22206
rect 7198 22146 7250 22158
rect 7198 22082 7250 22094
rect 11118 22146 11170 22158
rect 11118 22082 11170 22094
rect 16046 22146 16098 22158
rect 16046 22082 16098 22094
rect 16830 22146 16882 22158
rect 16830 22082 16882 22094
rect 25678 22146 25730 22158
rect 25678 22082 25730 22094
rect 672 21978 27888 22012
rect 672 21926 3806 21978
rect 3858 21926 3910 21978
rect 3962 21926 4014 21978
rect 4066 21926 23806 21978
rect 23858 21926 23910 21978
rect 23962 21926 24014 21978
rect 24066 21926 27888 21978
rect 672 21892 27888 21926
rect 14030 21698 14082 21710
rect 2706 21646 2718 21698
rect 2770 21646 2782 21698
rect 14030 21634 14082 21646
rect 14478 21698 14530 21710
rect 23998 21698 24050 21710
rect 18162 21646 18174 21698
rect 18226 21646 18238 21698
rect 27122 21646 27134 21698
rect 27186 21646 27198 21698
rect 14478 21634 14530 21646
rect 23998 21634 24050 21646
rect 7086 21586 7138 21598
rect 12126 21586 12178 21598
rect 16158 21586 16210 21598
rect 19294 21586 19346 21598
rect 20638 21586 20690 21598
rect 21982 21586 22034 21598
rect 5394 21534 5406 21586
rect 5458 21534 5470 21586
rect 6514 21534 6526 21586
rect 6578 21534 6590 21586
rect 7634 21534 7646 21586
rect 7698 21534 7710 21586
rect 8082 21534 8094 21586
rect 8146 21534 8158 21586
rect 10434 21534 10446 21586
rect 10498 21534 10510 21586
rect 14802 21534 14814 21586
rect 14866 21534 14878 21586
rect 15250 21534 15262 21586
rect 15314 21534 15326 21586
rect 16482 21534 16494 21586
rect 16546 21534 16558 21586
rect 17490 21534 17502 21586
rect 17554 21534 17566 21586
rect 19058 21534 19070 21586
rect 19122 21534 19134 21586
rect 19618 21534 19630 21586
rect 19682 21534 19694 21586
rect 20850 21534 20862 21586
rect 20914 21534 20926 21586
rect 21074 21534 21086 21586
rect 21138 21534 21150 21586
rect 22194 21534 22206 21586
rect 22258 21534 22270 21586
rect 23538 21534 23550 21586
rect 23602 21534 23614 21586
rect 26226 21534 26238 21586
rect 26290 21534 26302 21586
rect 7086 21522 7138 21534
rect 12126 21522 12178 21534
rect 16158 21522 16210 21534
rect 19294 21522 19346 21534
rect 20638 21522 20690 21534
rect 21982 21522 22034 21534
rect 8542 21474 8594 21486
rect 18510 21474 18562 21486
rect 3042 21422 3054 21474
rect 3106 21422 3118 21474
rect 7522 21422 7534 21474
rect 7586 21422 7598 21474
rect 15474 21422 15486 21474
rect 15538 21422 15550 21474
rect 8542 21410 8594 21422
rect 18510 21410 18562 21422
rect 18846 21474 18898 21486
rect 18846 21410 18898 21422
rect 20078 21474 20130 21486
rect 20078 21410 20130 21422
rect 21870 21474 21922 21486
rect 21870 21410 21922 21422
rect 25902 21474 25954 21486
rect 25902 21410 25954 21422
rect 4286 21362 4338 21374
rect 13470 21362 13522 21374
rect 10994 21310 11006 21362
rect 11058 21310 11070 21362
rect 4286 21298 4338 21310
rect 13470 21298 13522 21310
rect 18286 21362 18338 21374
rect 18286 21298 18338 21310
rect 19630 21362 19682 21374
rect 19630 21298 19682 21310
rect 19966 21362 20018 21374
rect 19966 21298 20018 21310
rect 25342 21362 25394 21374
rect 25342 21298 25394 21310
rect 672 21194 27888 21228
rect 672 21142 4466 21194
rect 4518 21142 4570 21194
rect 4622 21142 4674 21194
rect 4726 21142 24466 21194
rect 24518 21142 24570 21194
rect 24622 21142 24674 21194
rect 24726 21142 27888 21194
rect 672 21108 27888 21142
rect 17950 21026 18002 21038
rect 11330 20974 11342 21026
rect 11394 20974 11406 21026
rect 14914 20974 14926 21026
rect 14978 20974 14990 21026
rect 19730 20974 19742 21026
rect 19794 20974 19806 21026
rect 17950 20962 18002 20974
rect 1822 20914 1874 20926
rect 9438 20914 9490 20926
rect 3154 20862 3166 20914
rect 3218 20862 3230 20914
rect 6962 20862 6974 20914
rect 7026 20862 7038 20914
rect 1822 20850 1874 20862
rect 9438 20850 9490 20862
rect 10334 20914 10386 20926
rect 10334 20850 10386 20862
rect 16046 20914 16098 20926
rect 20190 20914 20242 20926
rect 16818 20862 16830 20914
rect 16882 20862 16894 20914
rect 17266 20862 17278 20914
rect 17330 20862 17342 20914
rect 16046 20850 16098 20862
rect 20190 20850 20242 20862
rect 25006 20914 25058 20926
rect 25006 20850 25058 20862
rect 26462 20914 26514 20926
rect 26462 20850 26514 20862
rect 27358 20914 27410 20926
rect 27358 20850 27410 20862
rect 3614 20802 3666 20814
rect 8878 20802 8930 20814
rect 12014 20802 12066 20814
rect 2594 20750 2606 20802
rect 2658 20750 2670 20802
rect 3042 20750 3054 20802
rect 3106 20750 3118 20802
rect 4386 20750 4398 20802
rect 4450 20750 4462 20802
rect 5282 20750 5294 20802
rect 5346 20750 5358 20802
rect 10770 20750 10782 20802
rect 10834 20750 10846 20802
rect 11106 20750 11118 20802
rect 11170 20750 11182 20802
rect 12338 20750 12350 20802
rect 12402 20750 12414 20802
rect 13346 20750 13358 20802
rect 13410 20750 13422 20802
rect 14354 20750 14366 20802
rect 14418 20750 14430 20802
rect 17154 20750 17166 20802
rect 17218 20750 17230 20802
rect 19058 20756 19070 20808
rect 19122 20756 19134 20808
rect 25566 20802 25618 20814
rect 19506 20750 19518 20802
rect 19570 20750 19582 20802
rect 20962 20750 20974 20802
rect 21026 20750 21038 20802
rect 21746 20750 21758 20802
rect 21810 20750 21822 20802
rect 3614 20738 3666 20750
rect 8878 20738 8930 20750
rect 12014 20738 12066 20750
rect 25566 20738 25618 20750
rect 25902 20802 25954 20814
rect 26898 20750 26910 20802
rect 26962 20750 26974 20802
rect 25902 20738 25954 20750
rect 2158 20690 2210 20702
rect 18734 20690 18786 20702
rect 1362 20638 1374 20690
rect 1426 20638 1438 20690
rect 7410 20638 7422 20690
rect 7474 20638 7486 20690
rect 2158 20626 2210 20638
rect 18734 20626 18786 20638
rect 5854 20578 5906 20590
rect 5854 20514 5906 20526
rect 17614 20578 17666 20590
rect 17614 20514 17666 20526
rect 672 20410 27888 20444
rect 672 20358 3806 20410
rect 3858 20358 3910 20410
rect 3962 20358 4014 20410
rect 4066 20358 23806 20410
rect 23858 20358 23910 20410
rect 23962 20358 24014 20410
rect 24066 20358 27888 20410
rect 672 20324 27888 20358
rect 5518 20242 5570 20254
rect 5518 20178 5570 20190
rect 11118 20242 11170 20254
rect 11118 20178 11170 20190
rect 3278 20130 3330 20142
rect 3278 20066 3330 20078
rect 6974 20130 7026 20142
rect 6974 20066 7026 20078
rect 19966 20130 20018 20142
rect 19966 20066 20018 20078
rect 20638 20130 20690 20142
rect 20962 20078 20974 20130
rect 21026 20078 21038 20130
rect 20638 20066 20690 20078
rect 8430 20018 8482 20030
rect 14478 20018 14530 20030
rect 26014 20018 26066 20030
rect 1698 19966 1710 20018
rect 1762 19966 1774 20018
rect 5170 19966 5182 20018
rect 5234 19966 5246 20018
rect 7298 19966 7310 20018
rect 7362 19966 7374 20018
rect 7858 19966 7870 20018
rect 7922 19966 7934 20018
rect 9090 19966 9102 20018
rect 9154 19966 9166 20018
rect 8430 19954 8482 19966
rect 9986 19961 9998 20013
rect 10050 19961 10062 20013
rect 10546 19966 10558 20018
rect 10610 19966 10622 20018
rect 13122 19966 13134 20018
rect 13186 19966 13198 20018
rect 13570 19966 13582 20018
rect 13634 19966 13646 20018
rect 14802 19966 14814 20018
rect 14866 19966 14878 20018
rect 15026 19966 15038 20018
rect 15090 19966 15102 20018
rect 15810 19966 15822 20018
rect 15874 19966 15886 20018
rect 16482 19966 16494 20018
rect 16546 19966 16558 20018
rect 19730 19966 19742 20018
rect 19794 19966 19806 20018
rect 14478 19954 14530 19966
rect 26014 19954 26066 19966
rect 26574 20018 26626 20030
rect 26574 19954 26626 19966
rect 27470 20018 27522 20030
rect 27470 19954 27522 19966
rect 12798 19906 12850 19918
rect 18622 19906 18674 19918
rect 7970 19854 7982 19906
rect 8034 19854 8046 19906
rect 13794 19854 13806 19906
rect 13858 19854 13870 19906
rect 17042 19854 17054 19906
rect 17106 19854 17118 19906
rect 12798 19842 12850 19854
rect 18622 19842 18674 19854
rect 20078 19906 20130 19918
rect 20078 19842 20130 19854
rect 20862 19906 20914 19918
rect 20862 19842 20914 19854
rect 26910 19906 26962 19918
rect 26910 19842 26962 19854
rect 18174 19794 18226 19806
rect 2146 19742 2158 19794
rect 2210 19742 2222 19794
rect 18174 19730 18226 19742
rect 18734 19794 18786 19806
rect 18734 19730 18786 19742
rect 18846 19794 18898 19806
rect 18846 19730 18898 19742
rect 672 19626 27888 19660
rect 672 19574 4466 19626
rect 4518 19574 4570 19626
rect 4622 19574 4674 19626
rect 4726 19574 24466 19626
rect 24518 19574 24570 19626
rect 24622 19574 24674 19626
rect 24726 19574 27888 19626
rect 672 19540 27888 19574
rect 27470 19458 27522 19470
rect 10882 19406 10894 19458
rect 10946 19406 10958 19458
rect 13458 19406 13470 19458
rect 13522 19406 13534 19458
rect 17378 19406 17390 19458
rect 17442 19406 17454 19458
rect 20290 19406 20302 19458
rect 20354 19406 20366 19458
rect 27470 19394 27522 19406
rect 6526 19346 6578 19358
rect 2258 19294 2270 19346
rect 2322 19294 2334 19346
rect 3378 19294 3390 19346
rect 3442 19294 3454 19346
rect 6066 19294 6078 19346
rect 6130 19294 6142 19346
rect 6526 19282 6578 19294
rect 9886 19346 9938 19358
rect 9886 19282 9938 19294
rect 12014 19346 12066 19358
rect 12014 19282 12066 19294
rect 19854 19346 19906 19358
rect 19854 19282 19906 19294
rect 25902 19346 25954 19358
rect 25902 19282 25954 19294
rect 26462 19346 26514 19358
rect 26462 19282 26514 19294
rect 4622 19234 4674 19246
rect 13918 19234 13970 19246
rect 16046 19234 16098 19246
rect 5394 19182 5406 19234
rect 5458 19182 5470 19234
rect 5842 19182 5854 19234
rect 5906 19182 5918 19234
rect 7074 19182 7086 19234
rect 7138 19182 7150 19234
rect 7298 19182 7310 19234
rect 7362 19182 7374 19234
rect 8194 19182 8206 19234
rect 8258 19182 8270 19234
rect 9426 19182 9438 19234
rect 9490 19182 9502 19234
rect 10322 19182 10334 19234
rect 10386 19182 10398 19234
rect 12786 19182 12798 19234
rect 12850 19182 12862 19234
rect 13234 19182 13246 19234
rect 13298 19182 13310 19234
rect 14466 19182 14478 19234
rect 14530 19182 14542 19234
rect 14690 19182 14702 19234
rect 14754 19182 14766 19234
rect 15474 19182 15486 19234
rect 15538 19182 15550 19234
rect 4622 19170 4674 19182
rect 13918 19170 13970 19182
rect 16046 19170 16098 19182
rect 16942 19234 16994 19246
rect 17390 19234 17442 19246
rect 17154 19182 17166 19234
rect 17218 19182 17230 19234
rect 17714 19182 17726 19234
rect 17778 19182 17790 19234
rect 18162 19182 18174 19234
rect 18226 19182 18238 19234
rect 19282 19182 19294 19234
rect 19346 19182 19358 19234
rect 20402 19182 20414 19234
rect 20466 19182 20478 19234
rect 20850 19182 20862 19234
rect 20914 19182 20926 19234
rect 16942 19170 16994 19182
rect 17390 19170 17442 19182
rect 1262 19122 1314 19134
rect 5070 19122 5122 19134
rect 3042 19070 3054 19122
rect 3106 19070 3118 19122
rect 1262 19058 1314 19070
rect 5070 19058 5122 19070
rect 12462 19122 12514 19134
rect 12462 19058 12514 19070
rect 21310 19122 21362 19134
rect 21310 19058 21362 19070
rect 26910 19122 26962 19134
rect 26910 19058 26962 19070
rect 16158 19010 16210 19022
rect 16158 18946 16210 18958
rect 672 18842 27888 18876
rect 672 18790 3806 18842
rect 3858 18790 3910 18842
rect 3962 18790 4014 18842
rect 4066 18790 23806 18842
rect 23858 18790 23910 18842
rect 23962 18790 24014 18842
rect 24066 18790 27888 18842
rect 672 18756 27888 18790
rect 12126 18674 12178 18686
rect 12126 18610 12178 18622
rect 14590 18674 14642 18686
rect 14590 18610 14642 18622
rect 2706 18510 2718 18562
rect 2770 18510 2782 18562
rect 5058 18510 5070 18562
rect 5122 18510 5134 18562
rect 6066 18510 6078 18562
rect 6130 18510 6142 18562
rect 8306 18510 8318 18562
rect 8370 18510 8382 18562
rect 10546 18510 10558 18562
rect 10610 18510 10622 18562
rect 13010 18510 13022 18562
rect 13074 18510 13086 18562
rect 1598 18450 1650 18462
rect 1598 18386 1650 18398
rect 2158 18450 2210 18462
rect 2158 18386 2210 18398
rect 5518 18450 5570 18462
rect 5518 18386 5570 18398
rect 7646 18450 7698 18462
rect 19070 18450 19122 18462
rect 26014 18450 26066 18462
rect 15810 18398 15822 18450
rect 15874 18398 15886 18450
rect 16594 18398 16606 18450
rect 16658 18398 16670 18450
rect 16818 18398 16830 18450
rect 16882 18398 16894 18450
rect 17938 18398 17950 18450
rect 18002 18398 18014 18450
rect 18498 18398 18510 18450
rect 18562 18398 18574 18450
rect 20962 18398 20974 18450
rect 21026 18398 21038 18450
rect 21410 18398 21422 18450
rect 21474 18398 21486 18450
rect 22642 18398 22654 18450
rect 22706 18398 22718 18450
rect 23650 18398 23662 18450
rect 23714 18398 23726 18450
rect 7646 18386 7698 18398
rect 19070 18386 19122 18398
rect 26014 18386 26066 18398
rect 26574 18450 26626 18462
rect 27346 18398 27358 18450
rect 27410 18398 27422 18450
rect 26574 18386 26626 18398
rect 17390 18338 17442 18350
rect 18846 18338 18898 18350
rect 8754 18286 8766 18338
rect 8818 18286 8830 18338
rect 13346 18286 13358 18338
rect 13410 18286 13422 18338
rect 17826 18286 17838 18338
rect 17890 18286 17902 18338
rect 17390 18274 17442 18286
rect 18846 18274 18898 18286
rect 20638 18338 20690 18350
rect 20638 18274 20690 18286
rect 22094 18338 22146 18350
rect 22094 18274 22146 18286
rect 26910 18338 26962 18350
rect 26910 18274 26962 18286
rect 4286 18226 4338 18238
rect 9886 18226 9938 18238
rect 19518 18226 19570 18238
rect 3154 18174 3166 18226
rect 3218 18174 3230 18226
rect 6514 18174 6526 18226
rect 6578 18174 6590 18226
rect 10994 18174 11006 18226
rect 11058 18174 11070 18226
rect 4286 18162 4338 18174
rect 9886 18162 9938 18174
rect 19518 18162 19570 18174
rect 19630 18226 19682 18238
rect 19630 18162 19682 18174
rect 19742 18226 19794 18238
rect 21634 18174 21646 18226
rect 21698 18174 21710 18226
rect 19742 18162 19794 18174
rect 672 18058 27888 18092
rect 672 18006 4466 18058
rect 4518 18006 4570 18058
rect 4622 18006 4674 18058
rect 4726 18006 24466 18058
rect 24518 18006 24570 18058
rect 24622 18006 24674 18058
rect 24726 18006 27888 18058
rect 672 17972 27888 18006
rect 13806 17890 13858 17902
rect 10434 17838 10446 17890
rect 10498 17838 10510 17890
rect 12674 17838 12686 17890
rect 12738 17838 12750 17890
rect 13806 17826 13858 17838
rect 16830 17890 16882 17902
rect 16830 17826 16882 17838
rect 21534 17890 21586 17902
rect 21534 17826 21586 17838
rect 27470 17890 27522 17902
rect 27470 17826 27522 17838
rect 5070 17778 5122 17790
rect 6526 17778 6578 17790
rect 3714 17726 3726 17778
rect 3778 17726 3790 17778
rect 6066 17726 6078 17778
rect 6130 17726 6142 17778
rect 5070 17714 5122 17726
rect 6526 17714 6578 17726
rect 8878 17778 8930 17790
rect 8878 17714 8930 17726
rect 9438 17778 9490 17790
rect 9438 17714 9490 17726
rect 17278 17778 17330 17790
rect 17278 17714 17330 17726
rect 17502 17778 17554 17790
rect 24558 17778 24610 17790
rect 18834 17726 18846 17778
rect 18898 17726 18910 17778
rect 22754 17726 22766 17778
rect 22818 17726 22830 17778
rect 17502 17714 17554 17726
rect 24558 17714 24610 17726
rect 26014 17778 26066 17790
rect 26014 17714 26066 17726
rect 26574 17778 26626 17790
rect 26574 17714 26626 17726
rect 26910 17778 26962 17790
rect 26910 17714 26962 17726
rect 1822 17671 1874 17683
rect 3278 17666 3330 17678
rect 15710 17666 15762 17678
rect 1822 17607 1874 17619
rect 2706 17614 2718 17666
rect 2770 17614 2782 17666
rect 3938 17614 3950 17666
rect 4002 17614 4014 17666
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 5394 17614 5406 17666
rect 5458 17614 5470 17666
rect 5954 17614 5966 17666
rect 6018 17614 6030 17666
rect 7298 17614 7310 17666
rect 7362 17614 7374 17666
rect 8194 17614 8206 17666
rect 8258 17614 8270 17666
rect 9986 17614 9998 17666
rect 10050 17614 10062 17666
rect 12114 17614 12126 17666
rect 12178 17614 12190 17666
rect 3278 17602 3330 17614
rect 15710 17602 15762 17614
rect 16718 17666 16770 17678
rect 19294 17666 19346 17678
rect 25118 17666 25170 17678
rect 18274 17614 18286 17666
rect 18338 17614 18350 17666
rect 18610 17614 18622 17666
rect 18674 17614 18686 17666
rect 20066 17614 20078 17666
rect 20130 17614 20142 17666
rect 20850 17614 20862 17666
rect 20914 17614 20926 17666
rect 16718 17602 16770 17614
rect 19294 17602 19346 17614
rect 25118 17602 25170 17614
rect 4734 17554 4786 17566
rect 17390 17554 17442 17566
rect 15250 17502 15262 17554
rect 15314 17502 15326 17554
rect 4734 17490 4786 17502
rect 17390 17490 17442 17502
rect 17838 17554 17890 17566
rect 23090 17502 23102 17554
rect 23154 17502 23166 17554
rect 17838 17490 17890 17502
rect 11566 17442 11618 17454
rect 11566 17378 11618 17390
rect 672 17274 27888 17308
rect 672 17222 3806 17274
rect 3858 17222 3910 17274
rect 3962 17222 4014 17274
rect 4066 17222 23806 17274
rect 23858 17222 23910 17274
rect 23962 17222 24014 17274
rect 24066 17222 27888 17274
rect 672 17188 27888 17222
rect 2830 17106 2882 17118
rect 2830 17042 2882 17054
rect 5966 17106 6018 17118
rect 5966 17042 6018 17054
rect 18286 17106 18338 17118
rect 18286 17042 18338 17054
rect 18510 17106 18562 17118
rect 18510 17042 18562 17054
rect 19966 17106 20018 17118
rect 19966 17042 20018 17054
rect 3838 16994 3890 17006
rect 26014 16994 26066 17006
rect 1250 16942 1262 16994
rect 1314 16942 1326 16994
rect 19618 16942 19630 16994
rect 19682 16942 19694 16994
rect 27010 16942 27022 16994
rect 27074 16942 27086 16994
rect 3838 16930 3890 16942
rect 26014 16930 26066 16942
rect 16158 16882 16210 16894
rect 18734 16882 18786 16894
rect 3378 16830 3390 16882
rect 3442 16830 3454 16882
rect 5058 16830 5070 16882
rect 5122 16830 5134 16882
rect 8418 16830 8430 16882
rect 8482 16830 8494 16882
rect 9314 16830 9326 16882
rect 9378 16830 9390 16882
rect 9874 16830 9886 16882
rect 9938 16830 9950 16882
rect 10546 16830 10558 16882
rect 10610 16830 10622 16882
rect 11218 16830 11230 16882
rect 11282 16830 11294 16882
rect 12002 16830 12014 16882
rect 12066 16830 12078 16882
rect 15026 16830 15038 16882
rect 15090 16830 15102 16882
rect 15474 16830 15486 16882
rect 15538 16830 15550 16882
rect 16930 16830 16942 16882
rect 16994 16830 17006 16882
rect 17714 16830 17726 16882
rect 17778 16830 17790 16882
rect 16158 16818 16210 16830
rect 18734 16818 18786 16830
rect 19182 16882 19234 16894
rect 19182 16818 19234 16830
rect 20974 16882 21026 16894
rect 26574 16882 26626 16894
rect 23874 16830 23886 16882
rect 23938 16830 23950 16882
rect 27346 16830 27358 16882
rect 27410 16830 27422 16882
rect 20974 16818 21026 16830
rect 26574 16818 26626 16830
rect 8990 16770 9042 16782
rect 1586 16718 1598 16770
rect 1650 16718 1662 16770
rect 8082 16718 8094 16770
rect 8146 16718 8158 16770
rect 8990 16706 9042 16718
rect 14702 16770 14754 16782
rect 18958 16770 19010 16782
rect 15698 16718 15710 16770
rect 15762 16718 15774 16770
rect 14702 16706 14754 16718
rect 18958 16706 19010 16718
rect 19070 16770 19122 16782
rect 19070 16706 19122 16718
rect 19742 16770 19794 16782
rect 19742 16706 19794 16718
rect 6862 16658 6914 16670
rect 20750 16658 20802 16670
rect 9986 16606 9998 16658
rect 10050 16606 10062 16658
rect 6862 16594 6914 16606
rect 20750 16594 20802 16606
rect 20862 16658 20914 16670
rect 20862 16594 20914 16606
rect 22206 16658 22258 16670
rect 23314 16606 23326 16658
rect 23378 16606 23390 16658
rect 22206 16594 22258 16606
rect 672 16490 27888 16524
rect 672 16438 4466 16490
rect 4518 16438 4570 16490
rect 4622 16438 4674 16490
rect 4726 16438 24466 16490
rect 24518 16438 24570 16490
rect 24622 16438 24674 16490
rect 24726 16438 27888 16490
rect 672 16404 27888 16438
rect 2942 16322 2994 16334
rect 5182 16322 5234 16334
rect 4050 16270 4062 16322
rect 4114 16270 4126 16322
rect 2942 16258 2994 16270
rect 5182 16258 5234 16270
rect 8206 16322 8258 16334
rect 12798 16322 12850 16334
rect 17950 16322 18002 16334
rect 27470 16322 27522 16334
rect 11666 16270 11678 16322
rect 11730 16270 11742 16322
rect 17042 16270 17054 16322
rect 17106 16270 17118 16322
rect 19954 16270 19966 16322
rect 20018 16270 20030 16322
rect 8206 16258 8258 16270
rect 12798 16258 12850 16270
rect 17950 16258 18002 16270
rect 27470 16258 27522 16270
rect 5966 16210 6018 16222
rect 10446 16210 10498 16222
rect 16046 16210 16098 16222
rect 1810 16158 1822 16210
rect 1874 16158 1886 16210
rect 6962 16158 6974 16210
rect 7026 16158 7038 16210
rect 13794 16158 13806 16210
rect 13858 16158 13870 16210
rect 5966 16146 6018 16158
rect 10446 16146 10498 16158
rect 16046 16146 16098 16158
rect 26014 16210 26066 16222
rect 26014 16146 26066 16158
rect 26910 16210 26962 16222
rect 26910 16146 26962 16158
rect 5854 16098 5906 16110
rect 1362 16046 1374 16098
rect 1426 16046 1438 16098
rect 3602 16046 3614 16098
rect 3666 16046 3678 16098
rect 5854 16034 5906 16046
rect 6190 16098 6242 16110
rect 16718 16098 16770 16110
rect 17838 16098 17890 16110
rect 9202 16046 9214 16098
rect 9266 16046 9278 16098
rect 9986 16046 9998 16098
rect 10050 16046 10062 16098
rect 11106 16046 11118 16098
rect 11170 16046 11182 16098
rect 13458 16046 13470 16098
rect 13522 16046 13534 16098
rect 15586 16046 15598 16098
rect 15650 16046 15662 16098
rect 16930 16046 16942 16098
rect 16994 16046 17006 16098
rect 17266 16046 17278 16098
rect 17330 16046 17342 16098
rect 6190 16034 6242 16046
rect 16718 16034 16770 16046
rect 17838 16034 17890 16046
rect 18174 16098 18226 16110
rect 18174 16034 18226 16046
rect 18286 16098 18338 16110
rect 18958 16098 19010 16110
rect 26574 16098 26626 16110
rect 18610 16046 18622 16098
rect 18674 16046 18686 16098
rect 19394 16046 19406 16098
rect 19458 16046 19470 16098
rect 19730 16046 19742 16098
rect 19794 16046 19806 16098
rect 20514 16046 20526 16098
rect 20578 16046 20590 16098
rect 21186 16046 21198 16098
rect 21250 16046 21262 16098
rect 22082 16046 22094 16098
rect 22146 16046 22158 16098
rect 18286 16034 18338 16046
rect 18958 16034 19010 16046
rect 26574 16034 26626 16046
rect 6626 15934 6638 15986
rect 6690 15934 6702 15986
rect 8878 15874 8930 15886
rect 8878 15810 8930 15822
rect 9214 15874 9266 15886
rect 9214 15810 9266 15822
rect 15038 15874 15090 15886
rect 17266 15822 17278 15874
rect 17330 15822 17342 15874
rect 15038 15810 15090 15822
rect 672 15706 27888 15740
rect 672 15654 3806 15706
rect 3858 15654 3910 15706
rect 3962 15654 4014 15706
rect 4066 15654 23806 15706
rect 23858 15654 23910 15706
rect 23962 15654 24014 15706
rect 24066 15654 27888 15706
rect 672 15620 27888 15654
rect 6750 15538 6802 15550
rect 6750 15474 6802 15486
rect 9886 15538 9938 15550
rect 9886 15474 9938 15486
rect 12126 15538 12178 15550
rect 18610 15486 18622 15538
rect 18674 15486 18686 15538
rect 12126 15474 12178 15486
rect 2158 15426 2210 15438
rect 20638 15426 20690 15438
rect 4162 15374 4174 15426
rect 4226 15374 4238 15426
rect 5170 15374 5182 15426
rect 5234 15374 5246 15426
rect 10546 15374 10558 15426
rect 10610 15374 10622 15426
rect 2158 15362 2210 15374
rect 20638 15362 20690 15374
rect 26014 15426 26066 15438
rect 26014 15362 26066 15374
rect 26910 15426 26962 15438
rect 26910 15362 26962 15374
rect 2606 15314 2658 15326
rect 1698 15262 1710 15314
rect 1762 15262 1774 15314
rect 2606 15250 2658 15262
rect 7086 15314 7138 15326
rect 7086 15250 7138 15262
rect 7534 15314 7586 15326
rect 7534 15250 7586 15262
rect 7758 15314 7810 15326
rect 14366 15314 14418 15326
rect 16158 15314 16210 15326
rect 18846 15314 18898 15326
rect 22094 15314 22146 15326
rect 8306 15262 8318 15314
rect 8370 15262 8382 15314
rect 15138 15262 15150 15314
rect 15202 15262 15214 15314
rect 15474 15262 15486 15314
rect 15538 15262 15550 15314
rect 16706 15262 16718 15314
rect 16770 15262 16782 15314
rect 16930 15262 16942 15314
rect 16994 15262 17006 15314
rect 17714 15262 17726 15314
rect 17778 15262 17790 15314
rect 18386 15262 18398 15314
rect 18450 15262 18462 15314
rect 19730 15262 19742 15314
rect 19794 15262 19806 15314
rect 20962 15262 20974 15314
rect 21026 15262 21038 15314
rect 21410 15262 21422 15314
rect 21474 15262 21486 15314
rect 22754 15262 22766 15314
rect 22818 15262 22830 15314
rect 23762 15262 23774 15314
rect 23826 15262 23838 15314
rect 27346 15262 27358 15314
rect 27410 15262 27422 15314
rect 7758 15250 7810 15262
rect 14366 15250 14418 15262
rect 16158 15250 16210 15262
rect 18846 15250 18898 15262
rect 22094 15250 22146 15262
rect 7310 15202 7362 15214
rect 3714 15150 3726 15202
rect 3778 15150 3790 15202
rect 5618 15150 5630 15202
rect 5682 15150 5694 15202
rect 7310 15138 7362 15150
rect 7646 15202 7698 15214
rect 14702 15202 14754 15214
rect 19182 15202 19234 15214
rect 8754 15150 8766 15202
rect 8818 15150 8830 15202
rect 10882 15150 10894 15202
rect 10946 15150 10958 15202
rect 15698 15150 15710 15202
rect 15762 15150 15774 15202
rect 7646 15138 7698 15150
rect 14702 15138 14754 15150
rect 19182 15138 19234 15150
rect 20078 15202 20130 15214
rect 20078 15138 20130 15150
rect 14030 15090 14082 15102
rect 14030 15026 14082 15038
rect 18398 15090 18450 15102
rect 18398 15026 18450 15038
rect 19966 15090 20018 15102
rect 26574 15090 26626 15102
rect 21634 15038 21646 15090
rect 21698 15038 21710 15090
rect 19966 15026 20018 15038
rect 26574 15026 26626 15038
rect 672 14922 27888 14956
rect 672 14870 4466 14922
rect 4518 14870 4570 14922
rect 4622 14870 4674 14922
rect 4726 14870 24466 14922
rect 24518 14870 24570 14922
rect 24622 14870 24674 14922
rect 24726 14870 27888 14922
rect 672 14836 27888 14870
rect 3278 14754 3330 14766
rect 9102 14754 9154 14766
rect 2146 14702 2158 14754
rect 2210 14702 2222 14754
rect 5730 14702 5742 14754
rect 5794 14702 5806 14754
rect 3278 14690 3330 14702
rect 9102 14690 9154 14702
rect 12462 14754 12514 14766
rect 16830 14754 16882 14766
rect 13570 14702 13582 14754
rect 13634 14702 13646 14754
rect 12462 14690 12514 14702
rect 16830 14690 16882 14702
rect 16942 14754 16994 14766
rect 27470 14754 27522 14766
rect 22530 14702 22542 14754
rect 22594 14702 22606 14754
rect 16942 14690 16994 14702
rect 27470 14690 27522 14702
rect 4174 14642 4226 14654
rect 4174 14578 4226 14590
rect 6862 14642 6914 14654
rect 6862 14578 6914 14590
rect 8878 14642 8930 14654
rect 8878 14578 8930 14590
rect 9326 14642 9378 14654
rect 14702 14642 14754 14654
rect 11330 14590 11342 14642
rect 11394 14590 11406 14642
rect 9326 14578 9378 14590
rect 14702 14578 14754 14590
rect 15710 14642 15762 14654
rect 15710 14578 15762 14590
rect 17726 14642 17778 14654
rect 26910 14642 26962 14654
rect 18722 14590 18734 14642
rect 18786 14590 18798 14642
rect 22642 14590 22654 14642
rect 22706 14590 22718 14642
rect 25106 14590 25118 14642
rect 25170 14590 25182 14642
rect 17726 14578 17778 14590
rect 26910 14578 26962 14590
rect 4286 14530 4338 14542
rect 7758 14530 7810 14542
rect 1698 14478 1710 14530
rect 1762 14478 1774 14530
rect 3938 14478 3950 14530
rect 4002 14478 4014 14530
rect 5170 14478 5182 14530
rect 5234 14478 5246 14530
rect 4286 14466 4338 14478
rect 7758 14466 7810 14478
rect 7982 14530 8034 14542
rect 7982 14466 8034 14478
rect 8206 14530 8258 14542
rect 8206 14466 8258 14478
rect 8766 14530 8818 14542
rect 15150 14530 15202 14542
rect 9874 14478 9886 14530
rect 9938 14478 9950 14530
rect 10770 14478 10782 14530
rect 10834 14478 10846 14530
rect 8766 14466 8818 14478
rect 15150 14466 15202 14478
rect 16046 14530 16098 14542
rect 16046 14466 16098 14478
rect 16718 14530 16770 14542
rect 18050 14478 18062 14530
rect 18114 14478 18126 14530
rect 18498 14478 18510 14530
rect 18562 14478 18574 14530
rect 19282 14478 19294 14530
rect 19346 14478 19358 14530
rect 19730 14478 19742 14530
rect 19794 14478 19806 14530
rect 20738 14478 20750 14530
rect 20802 14478 20814 14530
rect 16718 14466 16770 14478
rect 8082 14366 8094 14418
rect 8146 14366 8158 14418
rect 10210 14366 10222 14418
rect 10274 14366 10286 14418
rect 13122 14366 13134 14418
rect 13186 14366 13198 14418
rect 22978 14366 22990 14418
rect 23042 14366 23054 14418
rect 24770 14366 24782 14418
rect 24834 14366 24846 14418
rect 7310 14306 7362 14318
rect 4722 14254 4734 14306
rect 4786 14254 4798 14306
rect 7310 14242 7362 14254
rect 7534 14306 7586 14318
rect 7534 14242 7586 14254
rect 16158 14306 16210 14318
rect 16158 14242 16210 14254
rect 21422 14306 21474 14318
rect 21422 14242 21474 14254
rect 26350 14306 26402 14318
rect 26350 14242 26402 14254
rect 672 14138 27888 14172
rect 672 14086 3806 14138
rect 3858 14086 3910 14138
rect 3962 14086 4014 14138
rect 4066 14086 23806 14138
rect 23858 14086 23910 14138
rect 23962 14086 24014 14138
rect 24066 14086 27888 14138
rect 672 14052 27888 14086
rect 5518 13970 5570 13982
rect 5518 13906 5570 13918
rect 17390 13970 17442 13982
rect 17390 13906 17442 13918
rect 19070 13970 19122 13982
rect 19070 13906 19122 13918
rect 19294 13970 19346 13982
rect 19294 13906 19346 13918
rect 4398 13858 4450 13870
rect 8542 13858 8594 13870
rect 26014 13858 26066 13870
rect 6962 13806 6974 13858
rect 7026 13806 7038 13858
rect 12786 13806 12798 13858
rect 12850 13806 12862 13858
rect 19730 13806 19742 13858
rect 19794 13806 19806 13858
rect 27010 13806 27022 13858
rect 27074 13806 27086 13858
rect 4398 13794 4450 13806
rect 8542 13794 8594 13806
rect 26014 13794 26066 13806
rect 10670 13746 10722 13758
rect 17726 13746 17778 13758
rect 19518 13746 19570 13758
rect 1810 13694 1822 13746
rect 1874 13694 1886 13746
rect 3938 13694 3950 13746
rect 4002 13694 4014 13746
rect 9314 13694 9326 13746
rect 9378 13694 9390 13746
rect 9762 13694 9774 13746
rect 9826 13694 9838 13746
rect 10994 13694 11006 13746
rect 11058 13694 11070 13746
rect 11218 13694 11230 13746
rect 11282 13694 11294 13746
rect 12002 13694 12014 13746
rect 12066 13694 12078 13746
rect 14130 13694 14142 13746
rect 14194 13694 14206 13746
rect 14578 13694 14590 13746
rect 14642 13694 14654 13746
rect 15698 13694 15710 13746
rect 15762 13694 15774 13746
rect 16706 13694 16718 13746
rect 16770 13694 16782 13746
rect 18386 13694 18398 13746
rect 18450 13694 18462 13746
rect 10670 13682 10722 13694
rect 17726 13682 17778 13694
rect 19518 13682 19570 13694
rect 21422 13746 21474 13758
rect 26574 13746 26626 13758
rect 22978 13694 22990 13746
rect 23042 13694 23054 13746
rect 25218 13694 25230 13746
rect 25282 13694 25294 13746
rect 27346 13694 27358 13746
rect 27410 13694 27422 13746
rect 21422 13682 21474 13694
rect 26574 13682 26626 13694
rect 3390 13634 3442 13646
rect 8990 13634 9042 13646
rect 12910 13634 12962 13646
rect 4946 13582 4958 13634
rect 5010 13582 5022 13634
rect 7410 13582 7422 13634
rect 7474 13582 7486 13634
rect 9986 13582 9998 13634
rect 10050 13582 10062 13634
rect 3390 13570 3442 13582
rect 8990 13570 9042 13582
rect 12910 13570 12962 13582
rect 13134 13634 13186 13646
rect 13134 13570 13186 13582
rect 13694 13634 13746 13646
rect 15150 13634 15202 13646
rect 19966 13634 20018 13646
rect 14690 13582 14702 13634
rect 14754 13582 14766 13634
rect 18274 13582 18286 13634
rect 18338 13582 18350 13634
rect 13694 13570 13746 13582
rect 15150 13570 15202 13582
rect 19966 13570 20018 13582
rect 20638 13634 20690 13646
rect 20638 13570 20690 13582
rect 20862 13634 20914 13646
rect 24770 13582 24782 13634
rect 24834 13582 24846 13634
rect 20862 13570 20914 13582
rect 19742 13522 19794 13534
rect 2258 13470 2270 13522
rect 2322 13470 2334 13522
rect 19742 13458 19794 13470
rect 20750 13522 20802 13534
rect 23662 13522 23714 13534
rect 22530 13470 22542 13522
rect 22594 13470 22606 13522
rect 20750 13458 20802 13470
rect 23662 13458 23714 13470
rect 672 13354 27888 13388
rect 672 13302 4466 13354
rect 4518 13302 4570 13354
rect 4622 13302 4674 13354
rect 4726 13302 24466 13354
rect 24518 13302 24570 13354
rect 24622 13302 24674 13354
rect 24726 13302 27888 13354
rect 672 13268 27888 13302
rect 3614 13186 3666 13198
rect 3614 13122 3666 13134
rect 5742 13186 5794 13198
rect 5742 13122 5794 13134
rect 7870 13186 7922 13198
rect 7870 13122 7922 13134
rect 13806 13186 13858 13198
rect 13806 13122 13858 13134
rect 16046 13186 16098 13198
rect 16046 13122 16098 13134
rect 25118 13186 25170 13198
rect 25118 13122 25170 13134
rect 27470 13186 27522 13198
rect 27470 13122 27522 13134
rect 3166 13074 3218 13086
rect 1474 13022 1486 13074
rect 1538 13022 1550 13074
rect 3166 13010 3218 13022
rect 3502 13074 3554 13086
rect 18734 13074 18786 13086
rect 4610 13022 4622 13074
rect 4674 13022 4686 13074
rect 10322 13022 10334 13074
rect 10386 13022 10398 13074
rect 12674 13022 12686 13074
rect 12738 13022 12750 13074
rect 14914 13022 14926 13074
rect 14978 13022 14990 13074
rect 17826 13022 17838 13074
rect 17890 13022 17902 13074
rect 3502 13010 3554 13022
rect 18734 13010 18786 13022
rect 19182 13074 19234 13086
rect 24558 13074 24610 13086
rect 20178 13022 20190 13074
rect 20242 13022 20254 13074
rect 19182 13010 19234 13022
rect 24558 13010 24610 13022
rect 2606 12962 2658 12974
rect 7982 12962 8034 12974
rect 20862 12962 20914 12974
rect 26574 12962 26626 12974
rect 2034 12910 2046 12962
rect 2098 12910 2110 12962
rect 4162 12910 4174 12962
rect 4226 12910 4238 12962
rect 7410 12910 7422 12962
rect 7474 12910 7486 12962
rect 8866 12910 8878 12962
rect 8930 12910 8942 12962
rect 14354 12910 14366 12962
rect 14418 12910 14430 12962
rect 17938 12910 17950 12962
rect 18002 12910 18014 12962
rect 18386 12910 18398 12962
rect 18450 12910 18462 12962
rect 19618 12910 19630 12962
rect 19682 12910 19694 12962
rect 19954 12910 19966 12962
rect 20018 12910 20030 12962
rect 21410 12910 21422 12962
rect 21474 12910 21486 12962
rect 22194 12910 22206 12962
rect 22258 12910 22270 12962
rect 24994 12910 25006 12962
rect 25058 12910 25070 12962
rect 2606 12898 2658 12910
rect 7982 12898 8034 12910
rect 20862 12898 20914 12910
rect 26574 12898 26626 12910
rect 6414 12850 6466 12862
rect 26014 12850 26066 12862
rect 9986 12798 9998 12850
rect 10050 12798 10062 12850
rect 12226 12798 12238 12850
rect 12290 12798 12302 12850
rect 27010 12798 27022 12850
rect 27074 12798 27086 12850
rect 6414 12786 6466 12798
rect 26014 12786 26066 12798
rect 7870 12738 7922 12750
rect 7870 12674 7922 12686
rect 8206 12738 8258 12750
rect 8206 12674 8258 12686
rect 8878 12738 8930 12750
rect 8878 12674 8930 12686
rect 9214 12738 9266 12750
rect 9214 12674 9266 12686
rect 11566 12738 11618 12750
rect 11566 12674 11618 12686
rect 16830 12738 16882 12750
rect 16830 12674 16882 12686
rect 17166 12738 17218 12750
rect 17166 12674 17218 12686
rect 18398 12738 18450 12750
rect 18398 12674 18450 12686
rect 672 12570 27888 12604
rect 672 12518 3806 12570
rect 3858 12518 3910 12570
rect 3962 12518 4014 12570
rect 4066 12518 23806 12570
rect 23858 12518 23910 12570
rect 23962 12518 24014 12570
rect 24066 12518 27888 12570
rect 672 12484 27888 12518
rect 3614 12402 3666 12414
rect 3614 12338 3666 12350
rect 13022 12402 13074 12414
rect 18286 12402 18338 12414
rect 17490 12350 17502 12402
rect 17554 12350 17566 12402
rect 13022 12338 13074 12350
rect 18286 12338 18338 12350
rect 21534 12402 21586 12414
rect 21534 12338 21586 12350
rect 11006 12290 11058 12302
rect 5282 12238 5294 12290
rect 5346 12238 5358 12290
rect 9426 12238 9438 12290
rect 9490 12238 9502 12290
rect 11006 12226 11058 12238
rect 12014 12290 12066 12302
rect 12014 12226 12066 12238
rect 20750 12290 20802 12302
rect 20750 12226 20802 12238
rect 8766 12178 8818 12190
rect 16494 12178 16546 12190
rect 2034 12126 2046 12178
rect 2098 12126 2110 12178
rect 6066 12126 6078 12178
rect 6130 12126 6142 12178
rect 11554 12126 11566 12178
rect 11618 12126 11630 12178
rect 14018 12126 14030 12178
rect 14082 12126 14094 12178
rect 14802 12126 14814 12178
rect 14866 12126 14878 12178
rect 8766 12114 8818 12126
rect 16494 12114 16546 12126
rect 16942 12178 16994 12190
rect 18062 12178 18114 12190
rect 17154 12126 17166 12178
rect 17218 12126 17230 12178
rect 17602 12126 17614 12178
rect 17666 12126 17678 12178
rect 16942 12114 16994 12126
rect 18062 12114 18114 12126
rect 18510 12178 18562 12190
rect 18510 12114 18562 12126
rect 18958 12178 19010 12190
rect 18958 12114 19010 12126
rect 19518 12178 19570 12190
rect 19518 12114 19570 12126
rect 19630 12178 19682 12190
rect 20862 12178 20914 12190
rect 19954 12126 19966 12178
rect 20018 12126 20030 12178
rect 19630 12114 19682 12126
rect 20862 12114 20914 12126
rect 21646 12178 21698 12190
rect 26014 12178 26066 12190
rect 24210 12126 24222 12178
rect 24274 12126 24286 12178
rect 27346 12126 27358 12178
rect 27410 12126 27422 12178
rect 21646 12114 21698 12126
rect 26014 12114 26066 12126
rect 8542 12066 8594 12078
rect 2482 12014 2494 12066
rect 2546 12014 2558 12066
rect 6514 12014 6526 12066
rect 6578 12014 6590 12066
rect 7298 12014 7310 12066
rect 7362 12014 7374 12066
rect 8542 12002 8594 12014
rect 8654 12066 8706 12078
rect 26910 12066 26962 12078
rect 9762 12014 9774 12066
rect 9826 12014 9838 12066
rect 15250 12014 15262 12066
rect 15314 12014 15326 12066
rect 8654 12002 8706 12014
rect 26910 12002 26962 12014
rect 17726 11954 17778 11966
rect 8082 11902 8094 11954
rect 8146 11902 8158 11954
rect 17726 11890 17778 11902
rect 18734 11954 18786 11966
rect 18734 11890 18786 11902
rect 18846 11954 18898 11966
rect 18846 11890 18898 11902
rect 19406 11954 19458 11966
rect 19406 11890 19458 11902
rect 20638 11954 20690 11966
rect 20638 11890 20690 11902
rect 21086 11954 21138 11966
rect 21086 11890 21138 11902
rect 22542 11954 22594 11966
rect 26574 11954 26626 11966
rect 23650 11902 23662 11954
rect 23714 11902 23726 11954
rect 22542 11890 22594 11902
rect 26574 11890 26626 11902
rect 672 11786 27888 11820
rect 672 11734 4466 11786
rect 4518 11734 4570 11786
rect 4622 11734 4674 11786
rect 4726 11734 24466 11786
rect 24518 11734 24570 11786
rect 24622 11734 24674 11786
rect 24726 11734 27888 11786
rect 672 11700 27888 11734
rect 1598 11618 1650 11630
rect 8318 11618 8370 11630
rect 2706 11566 2718 11618
rect 2770 11566 2782 11618
rect 7522 11566 7534 11618
rect 7586 11566 7598 11618
rect 1598 11554 1650 11566
rect 8318 11554 8370 11566
rect 9774 11618 9826 11630
rect 9774 11554 9826 11566
rect 11454 11618 11506 11630
rect 11454 11554 11506 11566
rect 14142 11618 14194 11630
rect 14142 11554 14194 11566
rect 15598 11618 15650 11630
rect 23214 11618 23266 11630
rect 18722 11566 18734 11618
rect 18786 11566 18798 11618
rect 15598 11554 15650 11566
rect 23214 11554 23266 11566
rect 27470 11618 27522 11630
rect 27470 11554 27522 11566
rect 6638 11506 6690 11518
rect 5394 11454 5406 11506
rect 5458 11454 5470 11506
rect 6638 11442 6690 11454
rect 7086 11506 7138 11518
rect 7086 11442 7138 11454
rect 8206 11506 8258 11518
rect 8206 11442 8258 11454
rect 9886 11506 9938 11518
rect 9886 11442 9938 11454
rect 11006 11506 11058 11518
rect 11006 11442 11058 11454
rect 11118 11506 11170 11518
rect 16718 11506 16770 11518
rect 13010 11454 13022 11506
rect 13074 11454 13086 11506
rect 11118 11442 11170 11454
rect 16718 11442 16770 11454
rect 17054 11506 17106 11518
rect 17054 11442 17106 11454
rect 19182 11506 19234 11518
rect 19182 11442 19234 11454
rect 23774 11506 23826 11518
rect 23774 11442 23826 11454
rect 26014 11506 26066 11518
rect 26014 11442 26066 11454
rect 26910 11506 26962 11518
rect 26910 11442 26962 11454
rect 8990 11394 9042 11406
rect 3154 11342 3166 11394
rect 3218 11342 3230 11394
rect 3826 11342 3838 11394
rect 3890 11342 3902 11394
rect 7298 11342 7310 11394
rect 7362 11342 7374 11394
rect 7746 11342 7758 11394
rect 7810 11342 7822 11394
rect 8990 11330 9042 11342
rect 9102 11394 9154 11406
rect 9102 11330 9154 11342
rect 9326 11394 9378 11406
rect 9326 11330 9378 11342
rect 10782 11394 10834 11406
rect 10782 11330 10834 11342
rect 11678 11394 11730 11406
rect 26574 11394 26626 11406
rect 12002 11342 12014 11394
rect 12066 11342 12078 11394
rect 12450 11342 12462 11394
rect 12514 11342 12526 11394
rect 18050 11342 18062 11394
rect 18114 11342 18126 11394
rect 18498 11342 18510 11394
rect 18562 11342 18574 11394
rect 19842 11342 19854 11394
rect 19906 11342 19918 11394
rect 20850 11342 20862 11394
rect 20914 11342 20926 11394
rect 11678 11330 11730 11342
rect 26574 11330 26626 11342
rect 4286 11282 4338 11294
rect 11566 11282 11618 11294
rect 5058 11230 5070 11282
rect 5122 11230 5134 11282
rect 4286 11218 4338 11230
rect 11566 11218 11618 11230
rect 17726 11282 17778 11294
rect 17726 11218 17778 11230
rect 9438 11170 9490 11182
rect 7634 11118 7646 11170
rect 7698 11118 7710 11170
rect 9438 11106 9490 11118
rect 15374 11170 15426 11182
rect 15374 11106 15426 11118
rect 15710 11170 15762 11182
rect 15710 11106 15762 11118
rect 672 11002 27888 11036
rect 672 10950 3806 11002
rect 3858 10950 3910 11002
rect 3962 10950 4014 11002
rect 4066 10950 23806 11002
rect 23858 10950 23910 11002
rect 23962 10950 24014 11002
rect 24066 10950 27888 11002
rect 672 10916 27888 10950
rect 3614 10834 3666 10846
rect 3614 10770 3666 10782
rect 7198 10834 7250 10846
rect 18286 10834 18338 10846
rect 12002 10782 12014 10834
rect 12066 10782 12078 10834
rect 7198 10770 7250 10782
rect 18286 10770 18338 10782
rect 13246 10722 13298 10734
rect 17726 10722 17778 10734
rect 5170 10670 5182 10722
rect 5234 10670 5246 10722
rect 7970 10670 7982 10722
rect 8034 10670 8046 10722
rect 14690 10670 14702 10722
rect 14754 10670 14766 10722
rect 13246 10658 13298 10670
rect 17726 10658 17778 10670
rect 26014 10722 26066 10734
rect 27010 10670 27022 10722
rect 27074 10670 27086 10722
rect 26014 10658 26066 10670
rect 7422 10610 7474 10622
rect 7870 10610 7922 10622
rect 2034 10558 2046 10610
rect 2098 10558 2110 10610
rect 7746 10558 7758 10610
rect 7810 10558 7822 10610
rect 7422 10546 7474 10558
rect 7870 10546 7922 10558
rect 8766 10610 8818 10622
rect 11454 10610 11506 10622
rect 10882 10558 10894 10610
rect 10946 10558 10958 10610
rect 8766 10546 8818 10558
rect 11454 10546 11506 10558
rect 11902 10610 11954 10622
rect 12798 10610 12850 10622
rect 12114 10558 12126 10610
rect 12178 10558 12190 10610
rect 11902 10546 11954 10558
rect 12798 10546 12850 10558
rect 13022 10610 13074 10622
rect 13022 10546 13074 10558
rect 13470 10610 13522 10622
rect 13470 10546 13522 10558
rect 16606 10610 16658 10622
rect 17490 10558 17502 10610
rect 17554 10558 17566 10610
rect 19842 10558 19854 10610
rect 19906 10558 19918 10610
rect 27346 10558 27358 10610
rect 27410 10558 27422 10610
rect 16606 10546 16658 10558
rect 6750 10498 6802 10510
rect 5618 10446 5630 10498
rect 5682 10446 5694 10498
rect 6750 10434 6802 10446
rect 9326 10498 9378 10510
rect 9326 10434 9378 10446
rect 9662 10498 9714 10510
rect 9662 10434 9714 10446
rect 10110 10498 10162 10510
rect 10110 10434 10162 10446
rect 10670 10498 10722 10510
rect 10670 10434 10722 10446
rect 11118 10498 11170 10510
rect 17838 10498 17890 10510
rect 11666 10446 11678 10498
rect 11730 10446 11742 10498
rect 15026 10446 15038 10498
rect 15090 10446 15102 10498
rect 19394 10446 19406 10498
rect 19458 10446 19470 10498
rect 11118 10434 11170 10446
rect 17838 10434 17890 10446
rect 8094 10386 8146 10398
rect 2482 10334 2494 10386
rect 2546 10334 2558 10386
rect 8094 10322 8146 10334
rect 9550 10386 9602 10398
rect 9550 10322 9602 10334
rect 9886 10386 9938 10398
rect 9886 10322 9938 10334
rect 11230 10386 11282 10398
rect 11230 10322 11282 10334
rect 12238 10386 12290 10398
rect 12238 10322 12290 10334
rect 13582 10386 13634 10398
rect 13582 10322 13634 10334
rect 13694 10386 13746 10398
rect 13694 10322 13746 10334
rect 16270 10386 16322 10398
rect 16270 10322 16322 10334
rect 16942 10386 16994 10398
rect 16942 10322 16994 10334
rect 17166 10386 17218 10398
rect 17166 10322 17218 10334
rect 17278 10386 17330 10398
rect 17278 10322 17330 10334
rect 26574 10386 26626 10398
rect 26574 10322 26626 10334
rect 672 10218 27888 10252
rect 672 10166 4466 10218
rect 4518 10166 4570 10218
rect 4622 10166 4674 10218
rect 4726 10166 24466 10218
rect 24518 10166 24570 10218
rect 24622 10166 24674 10218
rect 24726 10166 27888 10218
rect 672 10132 27888 10166
rect 6526 10050 6578 10062
rect 13918 10050 13970 10062
rect 16046 10050 16098 10062
rect 27470 10050 27522 10062
rect 7410 9998 7422 10050
rect 7474 9998 7486 10050
rect 12674 9998 12686 10050
rect 12738 9998 12750 10050
rect 15250 9998 15262 10050
rect 15314 9998 15326 10050
rect 18946 9998 18958 10050
rect 19010 9998 19022 10050
rect 6526 9986 6578 9998
rect 13918 9986 13970 9998
rect 16046 9986 16098 9998
rect 27470 9986 27522 9998
rect 7086 9938 7138 9950
rect 2258 9886 2270 9938
rect 2322 9886 2334 9938
rect 5282 9886 5294 9938
rect 5346 9886 5358 9938
rect 7086 9874 7138 9886
rect 9102 9938 9154 9950
rect 13134 9938 13186 9950
rect 17166 9938 17218 9950
rect 10098 9886 10110 9938
rect 10162 9886 10174 9938
rect 15138 9886 15150 9938
rect 15202 9886 15214 9938
rect 9102 9874 9154 9886
rect 13134 9874 13186 9886
rect 17166 9874 17218 9886
rect 19406 9938 19458 9950
rect 19406 9874 19458 9886
rect 26910 9938 26962 9950
rect 26910 9874 26962 9886
rect 7534 9826 7586 9838
rect 10782 9826 10834 9838
rect 13246 9826 13298 9838
rect 14926 9826 14978 9838
rect 16158 9826 16210 9838
rect 3826 9774 3838 9826
rect 3890 9774 3902 9826
rect 4946 9774 4958 9826
rect 5010 9774 5022 9826
rect 7298 9774 7310 9826
rect 7362 9774 7374 9826
rect 7858 9774 7870 9826
rect 7922 9774 7934 9826
rect 9538 9774 9550 9826
rect 9602 9774 9614 9826
rect 9986 9774 9998 9826
rect 10050 9774 10062 9826
rect 11330 9774 11342 9826
rect 11394 9774 11406 9826
rect 12226 9774 12238 9826
rect 12290 9774 12302 9826
rect 13458 9774 13470 9826
rect 13522 9774 13534 9826
rect 13794 9774 13806 9826
rect 13858 9774 13870 9826
rect 15698 9774 15710 9826
rect 15762 9774 15774 9826
rect 7534 9762 7586 9774
rect 10782 9762 10834 9774
rect 13246 9762 13298 9774
rect 14926 9762 14978 9774
rect 16158 9762 16210 9774
rect 16606 9826 16658 9838
rect 16606 9762 16658 9774
rect 17054 9826 17106 9838
rect 17054 9762 17106 9774
rect 17278 9826 17330 9838
rect 25678 9826 25730 9838
rect 18386 9774 18398 9826
rect 18450 9774 18462 9826
rect 18834 9774 18846 9826
rect 18898 9774 18910 9826
rect 20066 9774 20078 9826
rect 20130 9774 20142 9826
rect 21074 9774 21086 9826
rect 21138 9774 21150 9826
rect 17278 9762 17330 9774
rect 25678 9762 25730 9774
rect 26574 9826 26626 9838
rect 26574 9762 26626 9774
rect 1262 9714 1314 9726
rect 1262 9650 1314 9662
rect 2830 9714 2882 9726
rect 2830 9650 2882 9662
rect 17950 9714 18002 9726
rect 17950 9650 18002 9662
rect 25118 9714 25170 9726
rect 25118 9650 25170 9662
rect 26014 9714 26066 9726
rect 26014 9650 26066 9662
rect 14030 9602 14082 9614
rect 14030 9538 14082 9550
rect 14254 9602 14306 9614
rect 15474 9550 15486 9602
rect 15538 9550 15550 9602
rect 14254 9538 14306 9550
rect 672 9434 27888 9468
rect 672 9382 3806 9434
rect 3858 9382 3910 9434
rect 3962 9382 4014 9434
rect 4066 9382 23806 9434
rect 23858 9382 23910 9434
rect 23962 9382 24014 9434
rect 24066 9382 27888 9434
rect 672 9348 27888 9382
rect 1262 9266 1314 9278
rect 1262 9202 1314 9214
rect 9662 9266 9714 9278
rect 9662 9202 9714 9214
rect 13806 9266 13858 9278
rect 13806 9202 13858 9214
rect 16494 9266 16546 9278
rect 16494 9202 16546 9214
rect 17054 9266 17106 9278
rect 17054 9202 17106 9214
rect 26462 9266 26514 9278
rect 26462 9202 26514 9214
rect 5518 9154 5570 9166
rect 3042 9102 3054 9154
rect 3106 9102 3118 9154
rect 5518 9090 5570 9102
rect 6414 9154 6466 9166
rect 6414 9090 6466 9102
rect 7422 9154 7474 9166
rect 25342 9154 25394 9166
rect 18610 9102 18622 9154
rect 18674 9102 18686 9154
rect 7422 9090 7474 9102
rect 25342 9090 25394 9102
rect 5854 9042 5906 9054
rect 7310 9042 7362 9054
rect 2258 8990 2270 9042
rect 2322 8990 2334 9042
rect 3826 8990 3838 9042
rect 3890 8990 3902 9042
rect 5058 8990 5070 9042
rect 5122 8990 5134 9042
rect 6962 8990 6974 9042
rect 7026 8990 7038 9042
rect 5854 8978 5906 8990
rect 7310 8978 7362 8990
rect 7534 9042 7586 9054
rect 8082 8990 8094 9042
rect 8146 8990 8158 9042
rect 10434 8990 10446 9042
rect 10498 8990 10510 9042
rect 12786 8990 12798 9042
rect 12850 8990 12862 9042
rect 14802 8990 14814 9042
rect 14866 8990 14878 9042
rect 27234 8990 27246 9042
rect 27298 8990 27310 9042
rect 7534 8978 7586 8990
rect 12126 8930 12178 8942
rect 10882 8878 10894 8930
rect 10946 8878 10958 8930
rect 18162 8878 18174 8930
rect 18226 8878 18238 8930
rect 12126 8866 12178 8878
rect 25902 8818 25954 8830
rect 8530 8766 8542 8818
rect 8594 8766 8606 8818
rect 15362 8766 15374 8818
rect 15426 8766 15438 8818
rect 25902 8754 25954 8766
rect 672 8650 27888 8684
rect 672 8598 4466 8650
rect 4518 8598 4570 8650
rect 4622 8598 4674 8650
rect 4726 8598 24466 8650
rect 24518 8598 24570 8650
rect 24622 8598 24674 8650
rect 24726 8598 27888 8650
rect 672 8564 27888 8598
rect 12238 8482 12290 8494
rect 12238 8418 12290 8430
rect 7198 8370 7250 8382
rect 3042 8318 3054 8370
rect 3106 8318 3118 8370
rect 6178 8318 6190 8370
rect 6242 8318 6254 8370
rect 7198 8306 7250 8318
rect 8094 8370 8146 8382
rect 8094 8306 8146 8318
rect 8206 8370 8258 8382
rect 14926 8370 14978 8382
rect 11106 8318 11118 8370
rect 11170 8318 11182 8370
rect 13234 8318 13246 8370
rect 13298 8318 13310 8370
rect 8206 8306 8258 8318
rect 14926 8306 14978 8318
rect 15598 8370 15650 8382
rect 15598 8306 15650 8318
rect 15710 8370 15762 8382
rect 15710 8306 15762 8318
rect 17614 8370 17666 8382
rect 17614 8306 17666 8318
rect 19518 8370 19570 8382
rect 20514 8318 20526 8370
rect 20578 8318 20590 8370
rect 19518 8306 19570 8318
rect 16942 8258 16994 8270
rect 17390 8258 17442 8270
rect 20974 8258 21026 8270
rect 2258 8206 2270 8258
rect 2322 8206 2334 8258
rect 3602 8206 3614 8258
rect 3666 8206 3678 8258
rect 6626 8206 6638 8258
rect 6690 8206 6702 8258
rect 10546 8206 10558 8258
rect 10610 8206 10622 8258
rect 15362 8206 15374 8258
rect 15426 8206 15438 8258
rect 17266 8206 17278 8258
rect 17330 8206 17342 8258
rect 19954 8206 19966 8258
rect 20018 8206 20030 8258
rect 20290 8206 20302 8258
rect 20354 8206 20366 8258
rect 21634 8206 21646 8258
rect 21698 8206 21710 8258
rect 22530 8206 22542 8258
rect 22594 8206 22606 8258
rect 27346 8206 27358 8258
rect 27410 8206 27422 8258
rect 16942 8194 16994 8206
rect 17390 8194 17442 8206
rect 20974 8194 21026 8206
rect 7758 8146 7810 8158
rect 26462 8146 26514 8158
rect 12898 8094 12910 8146
rect 12962 8094 12974 8146
rect 17490 8094 17502 8146
rect 17554 8094 17566 8146
rect 7758 8082 7810 8094
rect 26462 8082 26514 8094
rect 1262 8034 1314 8046
rect 1262 7970 1314 7982
rect 5070 8034 5122 8046
rect 5070 7970 5122 7982
rect 8206 8034 8258 8046
rect 8206 7970 8258 7982
rect 14478 8034 14530 8046
rect 14478 7970 14530 7982
rect 15038 8034 15090 8046
rect 16718 8034 16770 8046
rect 16146 7982 16158 8034
rect 16210 7982 16222 8034
rect 15038 7970 15090 7982
rect 16718 7970 16770 7982
rect 672 7866 27888 7900
rect 672 7814 3806 7866
rect 3858 7814 3910 7866
rect 3962 7814 4014 7866
rect 4066 7814 23806 7866
rect 23858 7814 23910 7866
rect 23962 7814 24014 7866
rect 24066 7814 27888 7866
rect 672 7780 27888 7814
rect 10894 7698 10946 7710
rect 10894 7634 10946 7646
rect 12238 7698 12290 7710
rect 12238 7634 12290 7646
rect 16606 7698 16658 7710
rect 16606 7634 16658 7646
rect 16718 7698 16770 7710
rect 16718 7634 16770 7646
rect 5518 7586 5570 7598
rect 1474 7534 1486 7586
rect 1538 7534 1550 7586
rect 2930 7534 2942 7586
rect 2994 7534 3006 7586
rect 5518 7522 5570 7534
rect 7310 7586 7362 7598
rect 26014 7586 26066 7598
rect 9314 7534 9326 7586
rect 9378 7534 9390 7586
rect 17042 7534 17054 7586
rect 17106 7534 17118 7586
rect 27010 7534 27022 7586
rect 27074 7534 27086 7586
rect 7310 7522 7362 7534
rect 26014 7522 26066 7534
rect 12126 7474 12178 7486
rect 14590 7474 14642 7486
rect 2258 7422 2270 7474
rect 2322 7422 2334 7474
rect 3826 7422 3838 7474
rect 3890 7422 3902 7474
rect 5058 7422 5070 7474
rect 5122 7422 5134 7474
rect 6850 7422 6862 7474
rect 6914 7422 6926 7474
rect 12898 7422 12910 7474
rect 12962 7422 12974 7474
rect 12126 7410 12178 7422
rect 14590 7410 14642 7422
rect 15934 7474 15986 7486
rect 16382 7474 16434 7486
rect 16146 7422 16158 7474
rect 16210 7422 16222 7474
rect 15934 7410 15986 7422
rect 16382 7410 16434 7422
rect 17390 7474 17442 7486
rect 17390 7410 17442 7422
rect 15598 7362 15650 7374
rect 9762 7310 9774 7362
rect 9826 7310 9838 7362
rect 13346 7310 13358 7362
rect 13410 7310 13422 7362
rect 15598 7298 15650 7310
rect 27470 7362 27522 7374
rect 27470 7298 27522 7310
rect 15710 7250 15762 7262
rect 15710 7186 15762 7198
rect 26574 7250 26626 7262
rect 26574 7186 26626 7198
rect 672 7082 27888 7116
rect 672 7030 4466 7082
rect 4518 7030 4570 7082
rect 4622 7030 4674 7082
rect 4726 7030 24466 7082
rect 24518 7030 24570 7082
rect 24622 7030 24674 7082
rect 24726 7030 27888 7082
rect 672 6996 27888 7030
rect 13918 6914 13970 6926
rect 13918 6850 13970 6862
rect 27470 6914 27522 6926
rect 27470 6850 27522 6862
rect 26014 6802 26066 6814
rect 12674 6750 12686 6802
rect 12738 6750 12750 6802
rect 26014 6738 26066 6750
rect 26910 6802 26962 6814
rect 26910 6738 26962 6750
rect 9662 6690 9714 6702
rect 11006 6690 11058 6702
rect 2034 6638 2046 6690
rect 2098 6638 2110 6690
rect 3826 6638 3838 6690
rect 3890 6638 3902 6690
rect 10098 6638 10110 6690
rect 10162 6638 10174 6690
rect 9662 6626 9714 6638
rect 11006 6626 11058 6638
rect 11566 6690 11618 6702
rect 26574 6690 26626 6702
rect 12338 6638 12350 6690
rect 12402 6638 12414 6690
rect 11566 6626 11618 6638
rect 26574 6626 26626 6638
rect 1362 6526 1374 6578
rect 1426 6526 1438 6578
rect 2830 6466 2882 6478
rect 2830 6402 2882 6414
rect 672 6298 27888 6332
rect 672 6246 3806 6298
rect 3858 6246 3910 6298
rect 3962 6246 4014 6298
rect 4066 6246 23806 6298
rect 23858 6246 23910 6298
rect 23962 6246 24014 6298
rect 24066 6246 27888 6298
rect 672 6212 27888 6246
rect 7758 6130 7810 6142
rect 7758 6066 7810 6078
rect 26462 6130 26514 6142
rect 26462 6066 26514 6078
rect 13806 6018 13858 6030
rect 1586 5966 1598 6018
rect 1650 5966 1662 6018
rect 9314 5966 9326 6018
rect 9378 5966 9390 6018
rect 12002 5966 12014 6018
rect 12066 5966 12078 6018
rect 13806 5954 13858 5966
rect 25342 6018 25394 6030
rect 25342 5954 25394 5966
rect 2606 5906 2658 5918
rect 2146 5854 2158 5906
rect 2210 5854 2222 5906
rect 14242 5854 14254 5906
rect 14306 5854 14318 5906
rect 14690 5854 14702 5906
rect 14754 5854 14766 5906
rect 16034 5854 16046 5906
rect 16098 5854 16110 5906
rect 16930 5854 16942 5906
rect 16994 5854 17006 5906
rect 27346 5854 27358 5906
rect 27410 5854 27422 5906
rect 2606 5842 2658 5854
rect 3166 5794 3218 5806
rect 3166 5730 3218 5742
rect 15262 5794 15314 5806
rect 15262 5730 15314 5742
rect 11566 5682 11618 5694
rect 25902 5682 25954 5694
rect 8866 5630 8878 5682
rect 8930 5630 8942 5682
rect 14802 5630 14814 5682
rect 14866 5630 14878 5682
rect 11566 5618 11618 5630
rect 25902 5618 25954 5630
rect 672 5514 27888 5548
rect 672 5462 4466 5514
rect 4518 5462 4570 5514
rect 4622 5462 4674 5514
rect 4726 5462 24466 5514
rect 24518 5462 24570 5514
rect 24622 5462 24674 5514
rect 24726 5462 27888 5514
rect 672 5428 27888 5462
rect 2606 5346 2658 5358
rect 2606 5282 2658 5294
rect 7758 5346 7810 5358
rect 14926 5346 14978 5358
rect 13794 5294 13806 5346
rect 13858 5294 13870 5346
rect 7758 5282 7810 5294
rect 14926 5282 14978 5294
rect 15374 5346 15426 5358
rect 15374 5282 15426 5294
rect 3166 5234 3218 5246
rect 1474 5182 1486 5234
rect 1538 5182 1550 5234
rect 3166 5170 3218 5182
rect 3502 5234 3554 5246
rect 3502 5170 3554 5182
rect 8318 5234 8370 5246
rect 8318 5170 8370 5182
rect 12798 5234 12850 5246
rect 12798 5170 12850 5182
rect 15934 5234 15986 5246
rect 26674 5182 26686 5234
rect 26738 5182 26750 5234
rect 15934 5170 15986 5182
rect 4062 5122 4114 5134
rect 2034 5070 2046 5122
rect 2098 5070 2110 5122
rect 12338 5070 12350 5122
rect 12402 5070 12414 5122
rect 13346 5070 13358 5122
rect 13410 5070 13422 5122
rect 27458 5070 27470 5122
rect 27522 5070 27534 5122
rect 4062 5058 4114 5070
rect 672 4730 27888 4764
rect 672 4678 3806 4730
rect 3858 4678 3910 4730
rect 3962 4678 4014 4730
rect 4066 4678 23806 4730
rect 23858 4678 23910 4730
rect 23962 4678 24014 4730
rect 24066 4678 27888 4730
rect 672 4644 27888 4678
rect 27470 4338 27522 4350
rect 27470 4274 27522 4286
rect 26910 4226 26962 4238
rect 1474 4174 1486 4226
rect 1538 4174 1550 4226
rect 2258 4174 2270 4226
rect 2322 4174 2334 4226
rect 26910 4162 26962 4174
rect 672 3946 27888 3980
rect 672 3894 4466 3946
rect 4518 3894 4570 3946
rect 4622 3894 4674 3946
rect 4726 3894 24466 3946
rect 24518 3894 24570 3946
rect 24622 3894 24674 3946
rect 24726 3894 27888 3946
rect 672 3860 27888 3894
rect 27470 3778 27522 3790
rect 27470 3714 27522 3726
rect 26910 3666 26962 3678
rect 26910 3602 26962 3614
rect 26574 3554 26626 3566
rect 2258 3502 2270 3554
rect 2322 3502 2334 3554
rect 26574 3490 26626 3502
rect 26114 3390 26126 3442
rect 26178 3390 26190 3442
rect 1262 3330 1314 3342
rect 1262 3266 1314 3278
rect 672 3162 27888 3196
rect 672 3110 3806 3162
rect 3858 3110 3910 3162
rect 3962 3110 4014 3162
rect 4066 3110 23806 3162
rect 23858 3110 23910 3162
rect 23962 3110 24014 3162
rect 24066 3110 27888 3162
rect 672 3076 27888 3110
rect 1474 2830 1486 2882
rect 1538 2830 1550 2882
rect 25218 2830 25230 2882
rect 25282 2830 25294 2882
rect 26114 2830 26126 2882
rect 26178 2830 26190 2882
rect 27010 2830 27022 2882
rect 27074 2830 27086 2882
rect 1038 2770 1090 2782
rect 1038 2706 1090 2718
rect 27470 2770 27522 2782
rect 27470 2706 27522 2718
rect 25678 2546 25730 2558
rect 25678 2482 25730 2494
rect 26574 2546 26626 2558
rect 26574 2482 26626 2494
rect 672 2378 27888 2412
rect 672 2326 4466 2378
rect 4518 2326 4570 2378
rect 4622 2326 4674 2378
rect 4726 2326 24466 2378
rect 24518 2326 24570 2378
rect 24622 2326 24674 2378
rect 24726 2326 27888 2378
rect 672 2292 27888 2326
rect 1038 2210 1090 2222
rect 1038 2146 1090 2158
rect 1598 2098 1650 2110
rect 1598 2034 1650 2046
rect 11454 2098 11506 2110
rect 11454 2034 11506 2046
rect 13246 2098 13298 2110
rect 13246 2034 13298 2046
rect 27470 2098 27522 2110
rect 27470 2034 27522 2046
rect 12014 1986 12066 1998
rect 12014 1922 12066 1934
rect 13806 1986 13858 1998
rect 26014 1986 26066 1998
rect 25554 1934 25566 1986
rect 25618 1934 25630 1986
rect 13806 1922 13858 1934
rect 26014 1922 26066 1934
rect 26910 1986 26962 1998
rect 26910 1922 26962 1934
rect 25218 1822 25230 1874
rect 25282 1822 25294 1874
rect 26450 1822 26462 1874
rect 26514 1822 26526 1874
rect 672 1594 27888 1628
rect 672 1542 3806 1594
rect 3858 1542 3910 1594
rect 3962 1542 4014 1594
rect 4066 1542 23806 1594
rect 23858 1542 23910 1594
rect 23962 1542 24014 1594
rect 24066 1542 27888 1594
rect 672 1508 27888 1542
rect 25678 1314 25730 1326
rect 7970 1262 7982 1314
rect 8034 1262 8046 1314
rect 24882 1262 24894 1314
rect 24946 1262 24958 1314
rect 25678 1250 25730 1262
rect 26574 1314 26626 1326
rect 26574 1250 26626 1262
rect 27134 1202 27186 1214
rect 27134 1138 27186 1150
rect 7534 978 7586 990
rect 7534 914 7586 926
rect 25342 978 25394 990
rect 25342 914 25394 926
rect 26238 978 26290 990
rect 26238 914 26290 926
rect 672 810 27888 844
rect 672 758 4466 810
rect 4518 758 4570 810
rect 4622 758 4674 810
rect 4726 758 24466 810
rect 24518 758 24570 810
rect 24622 758 24674 810
rect 24726 758 27888 810
rect 672 724 27888 758
<< via1 >>
rect 3806 56422 3858 56474
rect 3910 56422 3962 56474
rect 4014 56422 4066 56474
rect 23806 56422 23858 56474
rect 23910 56422 23962 56474
rect 24014 56422 24066 56474
rect 3614 56254 3666 56306
rect 5182 56254 5234 56306
rect 8990 56254 9042 56306
rect 10558 56254 10610 56306
rect 13022 56254 13074 56306
rect 14590 56254 14642 56306
rect 16494 56254 16546 56306
rect 18510 56254 18562 56306
rect 20302 56254 20354 56306
rect 22206 56254 22258 56306
rect 24446 56254 24498 56306
rect 26014 56254 26066 56306
rect 7422 56142 7474 56194
rect 21758 56030 21810 56082
rect 1038 55918 1090 55970
rect 3054 55918 3106 55970
rect 6190 55918 6242 55970
rect 8094 55918 8146 55970
rect 9998 55918 10050 55970
rect 11566 55918 11618 55970
rect 14030 55918 14082 55970
rect 15598 55918 15650 55970
rect 17502 55918 17554 55970
rect 19518 55918 19570 55970
rect 21310 55918 21362 55970
rect 23886 55918 23938 55970
rect 25454 55918 25506 55970
rect 1374 55806 1426 55858
rect 4466 55638 4518 55690
rect 4570 55638 4622 55690
rect 4674 55638 4726 55690
rect 24466 55638 24518 55690
rect 24570 55638 24622 55690
rect 24674 55638 24726 55690
rect 22990 55470 23042 55522
rect 21646 55358 21698 55410
rect 1038 55246 1090 55298
rect 3502 55246 3554 55298
rect 6302 55246 6354 55298
rect 12798 55246 12850 55298
rect 18286 55246 18338 55298
rect 19966 55246 20018 55298
rect 20526 55246 20578 55298
rect 20862 55246 20914 55298
rect 22430 55246 22482 55298
rect 24894 55246 24946 55298
rect 26238 55246 26290 55298
rect 1486 55134 1538 55186
rect 2494 55134 2546 55186
rect 6862 55134 6914 55186
rect 11902 55134 11954 55186
rect 17278 55134 17330 55186
rect 25678 55022 25730 55074
rect 27246 55022 27298 55074
rect 3806 54854 3858 54906
rect 3910 54854 3962 54906
rect 4014 54854 4066 54906
rect 23806 54854 23858 54906
rect 23910 54854 23962 54906
rect 24014 54854 24066 54906
rect 22542 54686 22594 54738
rect 23774 54686 23826 54738
rect 1486 54574 1538 54626
rect 19630 54574 19682 54626
rect 25566 54574 25618 54626
rect 21198 54462 21250 54514
rect 24110 54462 24162 54514
rect 24894 54462 24946 54514
rect 26350 54462 26402 54514
rect 21534 54350 21586 54402
rect 27022 54350 27074 54402
rect 1038 54238 1090 54290
rect 19070 54238 19122 54290
rect 20638 54238 20690 54290
rect 4466 54070 4518 54122
rect 4570 54070 4622 54122
rect 4674 54070 4726 54122
rect 24466 54070 24518 54122
rect 24570 54070 24622 54122
rect 24674 54070 24726 54122
rect 1038 53678 1090 53730
rect 22430 53678 22482 53730
rect 22766 53678 22818 53730
rect 23550 53678 23602 53730
rect 24670 53678 24722 53730
rect 26238 53678 26290 53730
rect 1598 53566 1650 53618
rect 21982 53566 22034 53618
rect 25678 53566 25730 53618
rect 27246 53454 27298 53506
rect 3806 53286 3858 53338
rect 3910 53286 3962 53338
rect 4014 53286 4066 53338
rect 23806 53286 23858 53338
rect 23910 53286 23962 53338
rect 24014 53286 24066 53338
rect 27134 53006 27186 53058
rect 23214 52894 23266 52946
rect 26462 52894 26514 52946
rect 1598 52782 1650 52834
rect 24670 52782 24722 52834
rect 25454 52782 25506 52834
rect 1038 52670 1090 52722
rect 23662 52670 23714 52722
rect 4466 52502 4518 52554
rect 4570 52502 4622 52554
rect 4674 52502 4726 52554
rect 24466 52502 24518 52554
rect 24570 52502 24622 52554
rect 24674 52502 24726 52554
rect 21982 52222 22034 52274
rect 26238 52222 26290 52274
rect 1038 52110 1090 52162
rect 1598 52110 1650 52162
rect 21422 52110 21474 52162
rect 22766 52110 22818 52162
rect 24894 52110 24946 52162
rect 23774 51998 23826 52050
rect 25678 51886 25730 51938
rect 27246 51886 27298 51938
rect 3806 51718 3858 51770
rect 3910 51718 3962 51770
rect 4014 51718 4066 51770
rect 23806 51718 23858 51770
rect 23910 51718 23962 51770
rect 24014 51718 24066 51770
rect 25678 51550 25730 51602
rect 1598 51214 1650 51266
rect 24670 51214 24722 51266
rect 26238 51214 26290 51266
rect 27022 51214 27074 51266
rect 1038 51102 1090 51154
rect 4466 50934 4518 50986
rect 4570 50934 4622 50986
rect 4674 50934 4726 50986
rect 24466 50934 24518 50986
rect 24570 50934 24622 50986
rect 24674 50934 24726 50986
rect 26238 50654 26290 50706
rect 1038 50542 1090 50594
rect 23886 50542 23938 50594
rect 24670 50542 24722 50594
rect 1598 50430 1650 50482
rect 23550 50430 23602 50482
rect 25678 50430 25730 50482
rect 27246 50318 27298 50370
rect 3806 50150 3858 50202
rect 3910 50150 3962 50202
rect 4014 50150 4066 50202
rect 23806 50150 23858 50202
rect 23910 50150 23962 50202
rect 24014 50150 24066 50202
rect 25678 49870 25730 49922
rect 27134 49870 27186 49922
rect 24670 49646 24722 49698
rect 26238 49646 26290 49698
rect 4466 49366 4518 49418
rect 4570 49366 4622 49418
rect 4674 49366 4726 49418
rect 24466 49366 24518 49418
rect 24570 49366 24622 49418
rect 24674 49366 24726 49418
rect 1038 48974 1090 49026
rect 24670 48974 24722 49026
rect 26238 48974 26290 49026
rect 1598 48862 1650 48914
rect 25678 48750 25730 48802
rect 27246 48750 27298 48802
rect 3806 48582 3858 48634
rect 3910 48582 3962 48634
rect 4014 48582 4066 48634
rect 23806 48582 23858 48634
rect 23910 48582 23962 48634
rect 24014 48582 24066 48634
rect 26462 48190 26514 48242
rect 1598 48078 1650 48130
rect 27022 48078 27074 48130
rect 1038 47966 1090 48018
rect 4466 47798 4518 47850
rect 4570 47798 4622 47850
rect 4674 47798 4726 47850
rect 24466 47798 24518 47850
rect 24570 47798 24622 47850
rect 24674 47798 24726 47850
rect 1038 47406 1090 47458
rect 24670 47406 24722 47458
rect 26238 47406 26290 47458
rect 25678 47294 25730 47346
rect 2046 47182 2098 47234
rect 27246 47182 27298 47234
rect 3806 47014 3858 47066
rect 3910 47014 3962 47066
rect 4014 47014 4066 47066
rect 23806 47014 23858 47066
rect 23910 47014 23962 47066
rect 24014 47014 24066 47066
rect 25678 46734 25730 46786
rect 27134 46734 27186 46786
rect 1598 46510 1650 46562
rect 2494 46510 2546 46562
rect 24670 46510 24722 46562
rect 26238 46510 26290 46562
rect 1038 46398 1090 46450
rect 1934 46398 1986 46450
rect 4466 46230 4518 46282
rect 4570 46230 4622 46282
rect 4674 46230 4726 46282
rect 24466 46230 24518 46282
rect 24570 46230 24622 46282
rect 24674 46230 24726 46282
rect 1150 45838 1202 45890
rect 24670 45838 24722 45890
rect 26238 45838 26290 45890
rect 1598 45726 1650 45778
rect 25678 45614 25730 45666
rect 27246 45614 27298 45666
rect 3806 45446 3858 45498
rect 3910 45446 3962 45498
rect 4014 45446 4066 45498
rect 23806 45446 23858 45498
rect 23910 45446 23962 45498
rect 24014 45446 24066 45498
rect 1598 44942 1650 44994
rect 26238 44942 26290 44994
rect 27022 44942 27074 44994
rect 1038 44830 1090 44882
rect 4466 44662 4518 44714
rect 4570 44662 4622 44714
rect 4674 44662 4726 44714
rect 24466 44662 24518 44714
rect 24570 44662 24622 44714
rect 24674 44662 24726 44714
rect 1038 44270 1090 44322
rect 24670 44270 24722 44322
rect 26238 44270 26290 44322
rect 1598 44158 1650 44210
rect 25678 44158 25730 44210
rect 27246 44046 27298 44098
rect 3806 43878 3858 43930
rect 3910 43878 3962 43930
rect 4014 43878 4066 43930
rect 23806 43878 23858 43930
rect 23910 43878 23962 43930
rect 24014 43878 24066 43930
rect 25678 43598 25730 43650
rect 26910 43598 26962 43650
rect 24894 43486 24946 43538
rect 1598 43374 1650 43426
rect 26238 43374 26290 43426
rect 1038 43262 1090 43314
rect 4466 43094 4518 43146
rect 4570 43094 4622 43146
rect 4674 43094 4726 43146
rect 24466 43094 24518 43146
rect 24570 43094 24622 43146
rect 24674 43094 24726 43146
rect 1038 42702 1090 42754
rect 1934 42702 1986 42754
rect 24670 42702 24722 42754
rect 26238 42702 26290 42754
rect 1598 42590 1650 42642
rect 2382 42590 2434 42642
rect 25678 42478 25730 42530
rect 27246 42478 27298 42530
rect 3806 42310 3858 42362
rect 3910 42310 3962 42362
rect 4014 42310 4066 42362
rect 23806 42310 23858 42362
rect 23910 42310 23962 42362
rect 24014 42310 24066 42362
rect 14142 41918 14194 41970
rect 1598 41806 1650 41858
rect 2494 41806 2546 41858
rect 14590 41806 14642 41858
rect 26238 41806 26290 41858
rect 27022 41806 27074 41858
rect 1038 41694 1090 41746
rect 1934 41694 1986 41746
rect 15822 41694 15874 41746
rect 4466 41526 4518 41578
rect 4570 41526 4622 41578
rect 4674 41526 4726 41578
rect 24466 41526 24518 41578
rect 24570 41526 24622 41578
rect 24674 41526 24726 41578
rect 10110 41246 10162 41298
rect 14366 41246 14418 41298
rect 1038 41134 1090 41186
rect 2046 41134 2098 41186
rect 10670 41134 10722 41186
rect 11790 41134 11842 41186
rect 24782 41134 24834 41186
rect 26462 41134 26514 41186
rect 1598 41022 1650 41074
rect 2494 41022 2546 41074
rect 12126 41022 12178 41074
rect 13918 41022 13970 41074
rect 25678 41022 25730 41074
rect 8990 40910 9042 40962
rect 15486 40910 15538 40962
rect 27246 40910 27298 40962
rect 3806 40742 3858 40794
rect 3910 40742 3962 40794
rect 4014 40742 4066 40794
rect 23806 40742 23858 40794
rect 23910 40742 23962 40794
rect 24014 40742 24066 40794
rect 2494 40462 2546 40514
rect 3278 40462 3330 40514
rect 25678 40462 25730 40514
rect 1150 40350 1202 40402
rect 1934 40350 1986 40402
rect 6078 40350 6130 40402
rect 6414 40350 6466 40402
rect 6862 40350 6914 40402
rect 8206 40350 8258 40402
rect 9214 40350 9266 40402
rect 10446 40350 10498 40402
rect 14366 40350 14418 40402
rect 26238 40350 26290 40402
rect 1598 40238 1650 40290
rect 7534 40238 7586 40290
rect 10894 40238 10946 40290
rect 12798 40238 12850 40290
rect 24670 40238 24722 40290
rect 27022 40238 27074 40290
rect 2830 40126 2882 40178
rect 7086 40126 7138 40178
rect 12126 40126 12178 40178
rect 13358 40126 13410 40178
rect 14926 40126 14978 40178
rect 16046 40126 16098 40178
rect 4466 39958 4518 40010
rect 4570 39958 4622 40010
rect 4674 39958 4726 40010
rect 24466 39958 24518 40010
rect 24570 39958 24622 40010
rect 24674 39958 24726 40010
rect 2494 39790 2546 39842
rect 6974 39790 7026 39842
rect 7870 39790 7922 39842
rect 2158 39678 2210 39730
rect 3054 39678 3106 39730
rect 7310 39678 7362 39730
rect 9550 39678 9602 39730
rect 1710 39566 1762 39618
rect 3950 39566 4002 39618
rect 8990 39566 9042 39618
rect 14030 39566 14082 39618
rect 24670 39566 24722 39618
rect 26238 39566 26290 39618
rect 3502 39454 3554 39506
rect 6526 39454 6578 39506
rect 10558 39454 10610 39506
rect 25678 39342 25730 39394
rect 27246 39342 27298 39394
rect 3806 39174 3858 39226
rect 3910 39174 3962 39226
rect 4014 39174 4066 39226
rect 23806 39174 23858 39226
rect 23910 39174 23962 39226
rect 24014 39174 24066 39226
rect 6974 39006 7026 39058
rect 1598 38894 1650 38946
rect 5406 38894 5458 38946
rect 12238 38894 12290 38946
rect 16942 38894 16994 38946
rect 2158 38782 2210 38834
rect 8318 38782 8370 38834
rect 8766 38782 8818 38834
rect 9438 38782 9490 38834
rect 10110 38782 10162 38834
rect 11006 38782 11058 38834
rect 11790 38782 11842 38834
rect 13134 38782 13186 38834
rect 13582 38782 13634 38834
rect 14254 38782 14306 38834
rect 14814 38782 14866 38834
rect 15822 38782 15874 38834
rect 5854 38670 5906 38722
rect 7982 38670 8034 38722
rect 8990 38670 9042 38722
rect 12798 38670 12850 38722
rect 13806 38670 13858 38722
rect 26238 38670 26290 38722
rect 27022 38670 27074 38722
rect 1038 38558 1090 38610
rect 2718 38558 2770 38610
rect 3838 38558 3890 38610
rect 16382 38558 16434 38610
rect 4466 38390 4518 38442
rect 4570 38390 4622 38442
rect 4674 38390 4726 38442
rect 24466 38390 24518 38442
rect 24570 38390 24622 38442
rect 24674 38390 24726 38442
rect 5966 38222 6018 38274
rect 8206 38222 8258 38274
rect 15150 38222 15202 38274
rect 1822 38110 1874 38162
rect 4734 38110 4786 38162
rect 6974 38110 7026 38162
rect 15710 38110 15762 38162
rect 6638 37998 6690 38050
rect 14702 37998 14754 38050
rect 24894 37998 24946 38050
rect 26238 37998 26290 38050
rect 1374 37886 1426 37938
rect 4398 37886 4450 37938
rect 9662 37886 9714 37938
rect 25678 37886 25730 37938
rect 26910 37886 26962 37938
rect 2942 37774 2994 37826
rect 3806 37606 3858 37658
rect 3910 37606 3962 37658
rect 4014 37606 4066 37658
rect 23806 37606 23858 37658
rect 23910 37606 23962 37658
rect 24014 37606 24066 37658
rect 8094 37438 8146 37490
rect 1710 37326 1762 37378
rect 2718 37326 2770 37378
rect 6526 37326 6578 37378
rect 12014 37326 12066 37378
rect 27134 37326 27186 37378
rect 2046 37214 2098 37266
rect 8654 37214 8706 37266
rect 13134 37214 13186 37266
rect 15486 37214 15538 37266
rect 15934 37214 15986 37266
rect 16606 37214 16658 37266
rect 17166 37214 17218 37266
rect 18174 37214 18226 37266
rect 9326 37102 9378 37154
rect 13582 37102 13634 37154
rect 15150 37102 15202 37154
rect 24670 37102 24722 37154
rect 25454 37102 25506 37154
rect 26238 37102 26290 37154
rect 3166 36990 3218 37042
rect 4286 36990 4338 37042
rect 6974 36990 7026 37042
rect 14702 36990 14754 37042
rect 16158 36990 16210 37042
rect 4466 36822 4518 36874
rect 4570 36822 4622 36874
rect 4674 36822 4726 36874
rect 24466 36822 24518 36874
rect 24570 36822 24622 36874
rect 24674 36822 24726 36874
rect 4174 36654 4226 36706
rect 7982 36654 8034 36706
rect 10222 36654 10274 36706
rect 10558 36654 10610 36706
rect 16718 36654 16770 36706
rect 6414 36542 6466 36594
rect 18286 36542 18338 36594
rect 19854 36542 19906 36594
rect 24670 36542 24722 36594
rect 2606 36430 2658 36482
rect 4734 36430 4786 36482
rect 6862 36430 6914 36482
rect 10894 36430 10946 36482
rect 17726 36430 17778 36482
rect 20414 36430 20466 36482
rect 26238 36430 26290 36482
rect 2158 36318 2210 36370
rect 7422 36318 7474 36370
rect 13582 36318 13634 36370
rect 17278 36318 17330 36370
rect 3054 36206 3106 36258
rect 5294 36206 5346 36258
rect 19406 36206 19458 36258
rect 25678 36206 25730 36258
rect 27246 36206 27298 36258
rect 3806 36038 3858 36090
rect 3910 36038 3962 36090
rect 4014 36038 4066 36090
rect 23806 36038 23858 36090
rect 23910 36038 23962 36090
rect 24014 36038 24066 36090
rect 2718 35758 2770 35810
rect 5518 35758 5570 35810
rect 6526 35758 6578 35810
rect 11790 35758 11842 35810
rect 3950 35646 4002 35698
rect 4398 35646 4450 35698
rect 8654 35646 8706 35698
rect 13582 35646 13634 35698
rect 2270 35534 2322 35586
rect 6862 35534 6914 35586
rect 9326 35534 9378 35586
rect 14814 35534 14866 35586
rect 26238 35534 26290 35586
rect 27022 35534 27074 35586
rect 1150 35422 1202 35474
rect 5966 35422 6018 35474
rect 8094 35422 8146 35474
rect 4466 35254 4518 35306
rect 4570 35254 4622 35306
rect 4674 35254 4726 35306
rect 24466 35254 24518 35306
rect 24570 35254 24622 35306
rect 24674 35254 24726 35306
rect 3838 35086 3890 35138
rect 4286 34974 4338 35026
rect 6974 34974 7026 35026
rect 14030 34974 14082 35026
rect 17950 34974 18002 35026
rect 19294 34974 19346 35026
rect 1038 34862 1090 34914
rect 1934 34862 1986 34914
rect 3166 34862 3218 34914
rect 3614 34862 3666 34914
rect 4846 34862 4898 34914
rect 5854 34862 5906 34914
rect 6526 34862 6578 34914
rect 9662 34862 9714 34914
rect 10894 34862 10946 34914
rect 17502 34862 17554 34914
rect 18734 34862 18786 34914
rect 19070 34862 19122 34914
rect 19854 34862 19906 34914
rect 20526 34862 20578 34914
rect 21310 34862 21362 34914
rect 24670 34862 24722 34914
rect 26238 34862 26290 34914
rect 1598 34750 1650 34802
rect 2494 34750 2546 34802
rect 2830 34750 2882 34802
rect 9998 34750 10050 34802
rect 18286 34750 18338 34802
rect 25678 34750 25730 34802
rect 8206 34638 8258 34690
rect 27246 34638 27298 34690
rect 3806 34470 3858 34522
rect 3910 34470 3962 34522
rect 4014 34470 4066 34522
rect 23806 34470 23858 34522
rect 23910 34470 23962 34522
rect 24014 34470 24066 34522
rect 18958 34302 19010 34354
rect 25678 34190 25730 34242
rect 27134 34190 27186 34242
rect 1486 34078 1538 34130
rect 1934 34078 1986 34130
rect 2830 34078 2882 34130
rect 3390 34078 3442 34130
rect 4286 34078 4338 34130
rect 5182 34078 5234 34130
rect 8206 34078 8258 34130
rect 9102 34078 9154 34130
rect 9662 34078 9714 34130
rect 10222 34078 10274 34130
rect 10782 34078 10834 34130
rect 11006 34078 11058 34130
rect 11790 34078 11842 34130
rect 12686 34078 12738 34130
rect 17390 34078 17442 34130
rect 19518 34078 19570 34130
rect 24894 34078 24946 34130
rect 1150 33966 1202 34018
rect 2158 33966 2210 34018
rect 8766 33966 8818 34018
rect 9774 33966 9826 34018
rect 13582 33966 13634 34018
rect 17838 33966 17890 34018
rect 20078 33966 20130 34018
rect 26238 33966 26290 34018
rect 5518 33854 5570 33906
rect 6638 33854 6690 33906
rect 7758 33854 7810 33906
rect 16270 33854 16322 33906
rect 4466 33686 4518 33738
rect 4570 33686 4622 33738
rect 4674 33686 4726 33738
rect 24466 33686 24518 33738
rect 24570 33686 24622 33738
rect 24674 33686 24726 33738
rect 2270 33406 2322 33458
rect 3278 33406 3330 33458
rect 7646 33406 7698 33458
rect 8878 33406 8930 33458
rect 10894 33406 10946 33458
rect 18734 33406 18786 33458
rect 1038 33294 1090 33346
rect 2718 33294 2770 33346
rect 3054 33294 3106 33346
rect 3726 33294 3778 33346
rect 4510 33294 4562 33346
rect 5294 33294 5346 33346
rect 8206 33294 8258 33346
rect 10334 33294 10386 33346
rect 12574 33294 12626 33346
rect 24894 33294 24946 33346
rect 26238 33294 26290 33346
rect 1598 33182 1650 33234
rect 9438 33182 9490 33234
rect 13246 33182 13298 33234
rect 15598 33182 15650 33234
rect 18398 33182 18450 33234
rect 6526 33070 6578 33122
rect 12014 33070 12066 33122
rect 19966 33070 20018 33122
rect 25678 33070 25730 33122
rect 27246 33070 27298 33122
rect 3806 32902 3858 32954
rect 3910 32902 3962 32954
rect 4014 32902 4066 32954
rect 23806 32902 23858 32954
rect 23910 32902 23962 32954
rect 24014 32902 24066 32954
rect 2830 32734 2882 32786
rect 3838 32622 3890 32674
rect 15598 32622 15650 32674
rect 19742 32622 19794 32674
rect 20750 32622 20802 32674
rect 22094 32622 22146 32674
rect 1150 32510 1202 32562
rect 3390 32510 3442 32562
rect 5070 32510 5122 32562
rect 7198 32510 7250 32562
rect 9886 32510 9938 32562
rect 14814 32510 14866 32562
rect 19294 32510 19346 32562
rect 21198 32510 21250 32562
rect 26462 32510 26514 32562
rect 1710 32398 1762 32450
rect 4958 32398 5010 32450
rect 7646 32398 7698 32450
rect 27022 32398 27074 32450
rect 5518 32286 5570 32338
rect 8878 32286 8930 32338
rect 10334 32286 10386 32338
rect 11454 32286 11506 32338
rect 21534 32286 21586 32338
rect 4466 32118 4518 32170
rect 4570 32118 4622 32170
rect 4674 32118 4726 32170
rect 24466 32118 24518 32170
rect 24570 32118 24622 32170
rect 24674 32118 24726 32170
rect 21198 31950 21250 32002
rect 2046 31838 2098 31890
rect 6078 31838 6130 31890
rect 9662 31838 9714 31890
rect 11118 31838 11170 31890
rect 12462 31838 12514 31890
rect 12910 31838 12962 31890
rect 17278 31838 17330 31890
rect 18510 31838 18562 31890
rect 1710 31726 1762 31778
rect 3278 31726 3330 31778
rect 5406 31726 5458 31778
rect 5966 31726 6018 31778
rect 6526 31726 6578 31778
rect 7310 31726 7362 31778
rect 8094 31726 8146 31778
rect 10222 31726 10274 31778
rect 11790 31726 11842 31778
rect 12238 31726 12290 31778
rect 13470 31726 13522 31778
rect 14478 31726 14530 31778
rect 16718 31726 16770 31778
rect 18062 31726 18114 31778
rect 20638 31726 20690 31778
rect 20974 31726 21026 31778
rect 21758 31726 21810 31778
rect 22430 31726 22482 31778
rect 23214 31726 23266 31778
rect 24670 31726 24722 31778
rect 26462 31726 26514 31778
rect 5070 31614 5122 31666
rect 10670 31614 10722 31666
rect 11454 31614 11506 31666
rect 20190 31614 20242 31666
rect 25678 31614 25730 31666
rect 27134 31614 27186 31666
rect 19742 31502 19794 31554
rect 3806 31334 3858 31386
rect 3910 31334 3962 31386
rect 4014 31334 4066 31386
rect 23806 31334 23858 31386
rect 23910 31334 23962 31386
rect 24014 31334 24066 31386
rect 4286 31166 4338 31218
rect 1598 31054 1650 31106
rect 2718 31054 2770 31106
rect 5518 31054 5570 31106
rect 6414 31054 6466 31106
rect 12238 31054 12290 31106
rect 5070 30942 5122 30994
rect 5966 30942 6018 30994
rect 6974 30942 7026 30994
rect 9102 30942 9154 30994
rect 9998 30942 10050 30994
rect 10558 30942 10610 30994
rect 11342 30942 11394 30994
rect 11790 30942 11842 30994
rect 13470 30942 13522 30994
rect 15822 30942 15874 30994
rect 16270 30942 16322 30994
rect 17726 30942 17778 30994
rect 18510 30942 18562 30994
rect 20974 30942 21026 30994
rect 21534 30942 21586 30994
rect 22094 30942 22146 30994
rect 22654 30942 22706 30994
rect 23662 30942 23714 30994
rect 24782 30942 24834 30994
rect 7310 30830 7362 30882
rect 11230 30830 11282 30882
rect 15038 30830 15090 30882
rect 15486 30830 15538 30882
rect 16494 30830 16546 30882
rect 16942 30830 16994 30882
rect 20638 30830 20690 30882
rect 21646 30830 21698 30882
rect 25454 30830 25506 30882
rect 26238 30830 26290 30882
rect 27022 30830 27074 30882
rect 1038 30718 1090 30770
rect 3166 30718 3218 30770
rect 8542 30718 8594 30770
rect 13918 30718 13970 30770
rect 4466 30550 4518 30602
rect 4570 30550 4622 30602
rect 4674 30550 4726 30602
rect 24466 30550 24518 30602
rect 24570 30550 24622 30602
rect 24674 30550 24726 30602
rect 17502 30382 17554 30434
rect 19742 30382 19794 30434
rect 20862 30382 20914 30434
rect 4510 30270 4562 30322
rect 10894 30270 10946 30322
rect 13582 30270 13634 30322
rect 21870 30270 21922 30322
rect 2270 30158 2322 30210
rect 2606 30158 2658 30210
rect 3838 30158 3890 30210
rect 4286 30158 4338 30210
rect 4958 30158 5010 30210
rect 5518 30158 5570 30210
rect 6526 30158 6578 30210
rect 7310 30158 7362 30210
rect 8878 30158 8930 30210
rect 12126 30158 12178 30210
rect 12574 30158 12626 30210
rect 12910 30158 12962 30210
rect 13358 30158 13410 30210
rect 14030 30158 14082 30210
rect 14590 30158 14642 30210
rect 15710 30158 15762 30210
rect 17054 30158 17106 30210
rect 19294 30158 19346 30210
rect 21422 30158 21474 30210
rect 23102 30158 23154 30210
rect 26238 30158 26290 30210
rect 1486 30046 1538 30098
rect 3054 30046 3106 30098
rect 3502 30046 3554 30098
rect 9438 30046 9490 30098
rect 10558 30046 10610 30098
rect 27134 30046 27186 30098
rect 8094 29934 8146 29986
rect 18622 29934 18674 29986
rect 3806 29766 3858 29818
rect 3910 29766 3962 29818
rect 4014 29766 4066 29818
rect 23806 29766 23858 29818
rect 23910 29766 23962 29818
rect 24014 29766 24066 29818
rect 4286 29598 4338 29650
rect 7198 29598 7250 29650
rect 10110 29598 10162 29650
rect 1598 29486 1650 29538
rect 8542 29486 8594 29538
rect 14030 29486 14082 29538
rect 2606 29374 2658 29426
rect 5630 29374 5682 29426
rect 13582 29374 13634 29426
rect 14702 29374 14754 29426
rect 15150 29374 15202 29426
rect 16046 29374 16098 29426
rect 16382 29374 16434 29426
rect 17502 29374 17554 29426
rect 18062 29374 18114 29426
rect 26238 29374 26290 29426
rect 3166 29262 3218 29314
rect 5966 29262 6018 29314
rect 11678 29262 11730 29314
rect 14366 29262 14418 29314
rect 18510 29262 18562 29314
rect 27022 29262 27074 29314
rect 1038 29150 1090 29202
rect 8990 29150 9042 29202
rect 12238 29150 12290 29202
rect 15374 29150 15426 29202
rect 19742 29150 19794 29202
rect 4466 28982 4518 29034
rect 4570 28982 4622 29034
rect 4674 28982 4726 29034
rect 24466 28982 24518 29034
rect 24570 28982 24622 29034
rect 24674 28982 24726 29034
rect 3614 28814 3666 28866
rect 12574 28814 12626 28866
rect 15486 28814 15538 28866
rect 17838 28814 17890 28866
rect 2382 28702 2434 28754
rect 9886 28702 9938 28754
rect 11566 28702 11618 28754
rect 20414 28702 20466 28754
rect 4174 28590 4226 28642
rect 5630 28590 5682 28642
rect 6190 28590 6242 28642
rect 7310 28590 7362 28642
rect 11118 28590 11170 28642
rect 11902 28590 11954 28642
rect 12350 28590 12402 28642
rect 13022 28590 13074 28642
rect 13582 28590 13634 28642
rect 14702 28590 14754 28642
rect 16046 28590 16098 28642
rect 19854 28590 19906 28642
rect 20302 28590 20354 28642
rect 21086 28590 21138 28642
rect 21422 28590 21474 28642
rect 21646 28590 21698 28642
rect 22430 28590 22482 28642
rect 26238 28590 26290 28642
rect 2046 28478 2098 28530
rect 4958 28478 5010 28530
rect 7982 28478 8034 28530
rect 9550 28478 9602 28530
rect 17390 28478 17442 28530
rect 19406 28478 19458 28530
rect 27134 28478 27186 28530
rect 18958 28366 19010 28418
rect 3806 28198 3858 28250
rect 3910 28198 3962 28250
rect 4014 28198 4066 28250
rect 23806 28198 23858 28250
rect 23910 28198 23962 28250
rect 24014 28198 24066 28250
rect 7422 28030 7474 28082
rect 12126 28030 12178 28082
rect 1038 27918 1090 27970
rect 13582 27918 13634 27970
rect 21198 27918 21250 27970
rect 25678 27918 25730 27970
rect 27134 27918 27186 27970
rect 1486 27806 1538 27858
rect 2270 27806 2322 27858
rect 6526 27806 6578 27858
rect 8094 27806 8146 27858
rect 10446 27806 10498 27858
rect 13918 27806 13970 27858
rect 14366 27806 14418 27858
rect 15262 27806 15314 27858
rect 15822 27806 15874 27858
rect 16606 27806 16658 27858
rect 18062 27806 18114 27858
rect 20638 27806 20690 27858
rect 24894 27806 24946 27858
rect 2718 27694 2770 27746
rect 5518 27694 5570 27746
rect 8654 27694 8706 27746
rect 11006 27694 11058 27746
rect 18510 27694 18562 27746
rect 26238 27694 26290 27746
rect 3950 27582 4002 27634
rect 4958 27582 5010 27634
rect 9774 27582 9826 27634
rect 14590 27582 14642 27634
rect 19742 27582 19794 27634
rect 4466 27414 4518 27466
rect 4570 27414 4622 27466
rect 4674 27414 4726 27466
rect 24466 27414 24518 27466
rect 24570 27414 24622 27466
rect 24674 27414 24726 27466
rect 1710 27246 1762 27298
rect 4286 27246 4338 27298
rect 10110 27246 10162 27298
rect 12014 27246 12066 27298
rect 13134 27246 13186 27298
rect 15374 27246 15426 27298
rect 8318 27134 8370 27186
rect 14142 27134 14194 27186
rect 17390 27134 17442 27186
rect 18398 27134 18450 27186
rect 27022 27134 27074 27186
rect 1262 27022 1314 27074
rect 3614 27022 3666 27074
rect 4062 27022 4114 27074
rect 4734 27022 4786 27074
rect 5294 27022 5346 27074
rect 6302 27022 6354 27074
rect 7870 27022 7922 27074
rect 13806 27022 13858 27074
rect 17726 27022 17778 27074
rect 18174 27022 18226 27074
rect 18958 27022 19010 27074
rect 19406 27022 19458 27074
rect 20526 27022 20578 27074
rect 24670 27022 24722 27074
rect 26238 27022 26290 27074
rect 3278 26910 3330 26962
rect 10558 26910 10610 26962
rect 11566 26910 11618 26962
rect 2830 26798 2882 26850
rect 8990 26798 9042 26850
rect 25678 26798 25730 26850
rect 3806 26630 3858 26682
rect 3910 26630 3962 26682
rect 4014 26630 4066 26682
rect 23806 26630 23858 26682
rect 23910 26630 23962 26682
rect 24014 26630 24066 26682
rect 3614 26462 3666 26514
rect 19966 26462 20018 26514
rect 27246 26462 27298 26514
rect 2046 26350 2098 26402
rect 5518 26350 5570 26402
rect 6414 26350 6466 26402
rect 17726 26350 17778 26402
rect 18398 26350 18450 26402
rect 9326 26238 9378 26290
rect 9886 26238 9938 26290
rect 10670 26238 10722 26290
rect 11118 26238 11170 26290
rect 12014 26238 12066 26290
rect 13246 26238 13298 26290
rect 15262 26238 15314 26290
rect 20750 26238 20802 26290
rect 2494 26126 2546 26178
rect 6750 26126 6802 26178
rect 8990 26126 9042 26178
rect 13694 26126 13746 26178
rect 15822 26126 15874 26178
rect 18734 26126 18786 26178
rect 26238 26126 26290 26178
rect 4958 26014 5010 26066
rect 7982 26014 8034 26066
rect 9998 26014 10050 26066
rect 14814 26014 14866 26066
rect 17278 26014 17330 26066
rect 21310 26014 21362 26066
rect 22430 26014 22482 26066
rect 4466 25846 4518 25898
rect 4570 25846 4622 25898
rect 4674 25846 4726 25898
rect 24466 25846 24518 25898
rect 24570 25846 24622 25898
rect 24674 25846 24726 25898
rect 3614 25678 3666 25730
rect 9550 25678 9602 25730
rect 10670 25678 10722 25730
rect 14926 25678 14978 25730
rect 18622 25678 18674 25730
rect 21310 25678 21362 25730
rect 7086 25566 7138 25618
rect 11678 25566 11730 25618
rect 19182 25566 19234 25618
rect 20078 25566 20130 25618
rect 22318 25566 22370 25618
rect 26238 25566 26290 25618
rect 2158 25454 2210 25506
rect 2942 25454 2994 25506
rect 3390 25454 3442 25506
rect 4062 25454 4114 25506
rect 4622 25454 4674 25506
rect 5742 25454 5794 25506
rect 6526 25454 6578 25506
rect 8990 25454 9042 25506
rect 11342 25454 11394 25506
rect 16830 25454 16882 25506
rect 17278 25454 17330 25506
rect 21758 25454 21810 25506
rect 24670 25454 24722 25506
rect 1262 25342 1314 25394
rect 2606 25342 2658 25394
rect 14478 25342 14530 25394
rect 19742 25342 19794 25394
rect 27246 25342 27298 25394
rect 8206 25230 8258 25282
rect 12910 25230 12962 25282
rect 16046 25230 16098 25282
rect 25678 25230 25730 25282
rect 3806 25062 3858 25114
rect 3910 25062 3962 25114
rect 4014 25062 4066 25114
rect 23806 25062 23858 25114
rect 23910 25062 23962 25114
rect 24014 25062 24066 25114
rect 3502 24894 3554 24946
rect 5518 24894 5570 24946
rect 11118 24782 11170 24834
rect 18734 24782 18786 24834
rect 20638 24782 20690 24834
rect 25566 24782 25618 24834
rect 27134 24782 27186 24834
rect 1822 24670 1874 24722
rect 5070 24670 5122 24722
rect 7422 24670 7474 24722
rect 7758 24670 7810 24722
rect 8430 24670 8482 24722
rect 9214 24670 9266 24722
rect 9998 24670 10050 24722
rect 10558 24670 10610 24722
rect 14926 24670 14978 24722
rect 15374 24670 15426 24722
rect 16046 24670 16098 24722
rect 16606 24670 16658 24722
rect 17502 24665 17554 24717
rect 21086 24670 21138 24722
rect 21422 24670 21474 24722
rect 22318 24670 22370 24722
rect 22654 24670 22706 24722
rect 23662 24670 23714 24722
rect 24894 24670 24946 24722
rect 26238 24670 26290 24722
rect 2382 24558 2434 24610
rect 6974 24558 7026 24610
rect 7982 24558 8034 24610
rect 13358 24558 13410 24610
rect 14590 24558 14642 24610
rect 21646 24558 21698 24610
rect 12798 24446 12850 24498
rect 15598 24446 15650 24498
rect 18174 24446 18226 24498
rect 4466 24278 4518 24330
rect 4570 24278 4622 24330
rect 4674 24278 4726 24330
rect 24466 24278 24518 24330
rect 24570 24278 24622 24330
rect 24674 24278 24726 24330
rect 1038 24110 1090 24162
rect 12238 24110 12290 24162
rect 17726 24110 17778 24162
rect 22094 24110 22146 24162
rect 1598 23998 1650 24050
rect 3390 23998 3442 24050
rect 6526 23998 6578 24050
rect 10334 23998 10386 24050
rect 16046 23998 16098 24050
rect 20974 23998 21026 24050
rect 22542 23998 22594 24050
rect 23102 23998 23154 24050
rect 24670 23998 24722 24050
rect 2382 23886 2434 23938
rect 2830 23886 2882 23938
rect 3166 23886 3218 23938
rect 4062 23886 4114 23938
rect 4622 23886 4674 23938
rect 5518 23886 5570 23938
rect 6078 23886 6130 23938
rect 10894 23886 10946 23938
rect 11566 23886 11618 23938
rect 12014 23886 12066 23938
rect 12910 23886 12962 23938
rect 13470 23886 13522 23938
rect 14366 23886 14418 23938
rect 15486 23886 15538 23938
rect 17054 23886 17106 23938
rect 17502 23886 17554 23938
rect 18174 23886 18226 23938
rect 18734 23886 18786 23938
rect 18958 23886 19010 23938
rect 19854 23886 19906 23938
rect 20526 23886 20578 23938
rect 26238 23886 26290 23938
rect 6190 23774 6242 23826
rect 11230 23774 11282 23826
rect 16718 23774 16770 23826
rect 27246 23774 27298 23826
rect 7758 23662 7810 23714
rect 25678 23662 25730 23714
rect 3806 23494 3858 23546
rect 3910 23494 3962 23546
rect 4014 23494 4066 23546
rect 23806 23494 23858 23546
rect 23910 23494 23962 23546
rect 24014 23494 24066 23546
rect 3838 23326 3890 23378
rect 16270 23326 16322 23378
rect 2270 23214 2322 23266
rect 5294 23214 5346 23266
rect 13246 23214 13298 23266
rect 27134 23214 27186 23266
rect 1598 23102 1650 23154
rect 6302 23102 6354 23154
rect 9326 23102 9378 23154
rect 10334 23102 10386 23154
rect 14702 23102 14754 23154
rect 19966 23102 20018 23154
rect 1150 22990 1202 23042
rect 2718 22990 2770 23042
rect 6862 22990 6914 23042
rect 8878 22990 8930 23042
rect 15150 22990 15202 23042
rect 19630 22990 19682 23042
rect 26238 22990 26290 23042
rect 5742 22878 5794 22930
rect 7758 22878 7810 22930
rect 10894 22878 10946 22930
rect 12014 22878 12066 22930
rect 13806 22878 13858 22930
rect 19854 22878 19906 22930
rect 20078 22878 20130 22930
rect 4466 22710 4518 22762
rect 4570 22710 4622 22762
rect 4674 22710 4726 22762
rect 24466 22710 24518 22762
rect 24570 22710 24622 22762
rect 24674 22710 24726 22762
rect 2830 22542 2882 22594
rect 12238 22542 12290 22594
rect 13358 22542 13410 22594
rect 1598 22430 1650 22482
rect 6078 22430 6130 22482
rect 9998 22430 10050 22482
rect 14814 22430 14866 22482
rect 17950 22430 18002 22482
rect 20302 22430 20354 22482
rect 23438 22430 23490 22482
rect 26238 22430 26290 22482
rect 4286 22318 4338 22370
rect 9550 22318 9602 22370
rect 14366 22318 14418 22370
rect 18398 22318 18450 22370
rect 19630 22318 19682 22370
rect 20078 22318 20130 22370
rect 20750 22318 20802 22370
rect 21310 22318 21362 22370
rect 22430 22318 22482 22370
rect 22878 22318 22930 22370
rect 24894 22318 24946 22370
rect 1262 22206 1314 22258
rect 3502 22206 3554 22258
rect 5630 22206 5682 22258
rect 11790 22206 11842 22258
rect 19294 22206 19346 22258
rect 27246 22206 27298 22258
rect 7198 22094 7250 22146
rect 11118 22094 11170 22146
rect 16046 22094 16098 22146
rect 16830 22094 16882 22146
rect 25678 22094 25730 22146
rect 3806 21926 3858 21978
rect 3910 21926 3962 21978
rect 4014 21926 4066 21978
rect 23806 21926 23858 21978
rect 23910 21926 23962 21978
rect 24014 21926 24066 21978
rect 2718 21646 2770 21698
rect 14030 21646 14082 21698
rect 14478 21646 14530 21698
rect 18174 21646 18226 21698
rect 23998 21646 24050 21698
rect 27134 21646 27186 21698
rect 5406 21534 5458 21586
rect 6526 21534 6578 21586
rect 7086 21534 7138 21586
rect 7646 21534 7698 21586
rect 8094 21534 8146 21586
rect 10446 21534 10498 21586
rect 12126 21534 12178 21586
rect 14814 21534 14866 21586
rect 15262 21534 15314 21586
rect 16158 21534 16210 21586
rect 16494 21534 16546 21586
rect 17502 21534 17554 21586
rect 19070 21534 19122 21586
rect 19294 21534 19346 21586
rect 19630 21534 19682 21586
rect 20638 21534 20690 21586
rect 20862 21534 20914 21586
rect 21086 21534 21138 21586
rect 21982 21534 22034 21586
rect 22206 21534 22258 21586
rect 23550 21534 23602 21586
rect 26238 21534 26290 21586
rect 3054 21422 3106 21474
rect 7534 21422 7586 21474
rect 8542 21422 8594 21474
rect 15486 21422 15538 21474
rect 18510 21422 18562 21474
rect 18846 21422 18898 21474
rect 20078 21422 20130 21474
rect 21870 21422 21922 21474
rect 25902 21422 25954 21474
rect 4286 21310 4338 21362
rect 11006 21310 11058 21362
rect 13470 21310 13522 21362
rect 18286 21310 18338 21362
rect 19630 21310 19682 21362
rect 19966 21310 20018 21362
rect 25342 21310 25394 21362
rect 4466 21142 4518 21194
rect 4570 21142 4622 21194
rect 4674 21142 4726 21194
rect 24466 21142 24518 21194
rect 24570 21142 24622 21194
rect 24674 21142 24726 21194
rect 11342 20974 11394 21026
rect 14926 20974 14978 21026
rect 17950 20974 18002 21026
rect 19742 20974 19794 21026
rect 1822 20862 1874 20914
rect 3166 20862 3218 20914
rect 6974 20862 7026 20914
rect 9438 20862 9490 20914
rect 10334 20862 10386 20914
rect 16046 20862 16098 20914
rect 16830 20862 16882 20914
rect 17278 20862 17330 20914
rect 20190 20862 20242 20914
rect 25006 20862 25058 20914
rect 26462 20862 26514 20914
rect 27358 20862 27410 20914
rect 2606 20750 2658 20802
rect 3054 20750 3106 20802
rect 3614 20750 3666 20802
rect 4398 20750 4450 20802
rect 5294 20750 5346 20802
rect 8878 20750 8930 20802
rect 10782 20750 10834 20802
rect 11118 20750 11170 20802
rect 12014 20750 12066 20802
rect 12350 20750 12402 20802
rect 13358 20750 13410 20802
rect 14366 20750 14418 20802
rect 17166 20750 17218 20802
rect 19070 20756 19122 20808
rect 19518 20750 19570 20802
rect 20974 20750 21026 20802
rect 21758 20750 21810 20802
rect 25566 20750 25618 20802
rect 25902 20750 25954 20802
rect 26910 20750 26962 20802
rect 1374 20638 1426 20690
rect 2158 20638 2210 20690
rect 7422 20638 7474 20690
rect 18734 20638 18786 20690
rect 5854 20526 5906 20578
rect 17614 20526 17666 20578
rect 3806 20358 3858 20410
rect 3910 20358 3962 20410
rect 4014 20358 4066 20410
rect 23806 20358 23858 20410
rect 23910 20358 23962 20410
rect 24014 20358 24066 20410
rect 5518 20190 5570 20242
rect 11118 20190 11170 20242
rect 3278 20078 3330 20130
rect 6974 20078 7026 20130
rect 19966 20078 20018 20130
rect 20638 20078 20690 20130
rect 20974 20078 21026 20130
rect 1710 19966 1762 20018
rect 5182 19966 5234 20018
rect 7310 19966 7362 20018
rect 7870 19966 7922 20018
rect 8430 19966 8482 20018
rect 9102 19966 9154 20018
rect 9998 19961 10050 20013
rect 10558 19966 10610 20018
rect 13134 19966 13186 20018
rect 13582 19966 13634 20018
rect 14478 19966 14530 20018
rect 14814 19966 14866 20018
rect 15038 19966 15090 20018
rect 15822 19966 15874 20018
rect 16494 19966 16546 20018
rect 19742 19966 19794 20018
rect 26014 19966 26066 20018
rect 26574 19966 26626 20018
rect 27470 19966 27522 20018
rect 7982 19854 8034 19906
rect 12798 19854 12850 19906
rect 13806 19854 13858 19906
rect 17054 19854 17106 19906
rect 18622 19854 18674 19906
rect 20078 19854 20130 19906
rect 20862 19854 20914 19906
rect 26910 19854 26962 19906
rect 2158 19742 2210 19794
rect 18174 19742 18226 19794
rect 18734 19742 18786 19794
rect 18846 19742 18898 19794
rect 4466 19574 4518 19626
rect 4570 19574 4622 19626
rect 4674 19574 4726 19626
rect 24466 19574 24518 19626
rect 24570 19574 24622 19626
rect 24674 19574 24726 19626
rect 10894 19406 10946 19458
rect 13470 19406 13522 19458
rect 17390 19406 17442 19458
rect 20302 19406 20354 19458
rect 27470 19406 27522 19458
rect 2270 19294 2322 19346
rect 3390 19294 3442 19346
rect 6078 19294 6130 19346
rect 6526 19294 6578 19346
rect 9886 19294 9938 19346
rect 12014 19294 12066 19346
rect 19854 19294 19906 19346
rect 25902 19294 25954 19346
rect 26462 19294 26514 19346
rect 4622 19182 4674 19234
rect 5406 19182 5458 19234
rect 5854 19182 5906 19234
rect 7086 19182 7138 19234
rect 7310 19182 7362 19234
rect 8206 19182 8258 19234
rect 9438 19182 9490 19234
rect 10334 19182 10386 19234
rect 12798 19182 12850 19234
rect 13246 19182 13298 19234
rect 13918 19182 13970 19234
rect 14478 19182 14530 19234
rect 14702 19182 14754 19234
rect 15486 19182 15538 19234
rect 16046 19182 16098 19234
rect 16942 19182 16994 19234
rect 17166 19182 17218 19234
rect 17390 19182 17442 19234
rect 17726 19182 17778 19234
rect 18174 19182 18226 19234
rect 19294 19182 19346 19234
rect 20414 19182 20466 19234
rect 20862 19182 20914 19234
rect 1262 19070 1314 19122
rect 3054 19070 3106 19122
rect 5070 19070 5122 19122
rect 12462 19070 12514 19122
rect 21310 19070 21362 19122
rect 26910 19070 26962 19122
rect 16158 18958 16210 19010
rect 3806 18790 3858 18842
rect 3910 18790 3962 18842
rect 4014 18790 4066 18842
rect 23806 18790 23858 18842
rect 23910 18790 23962 18842
rect 24014 18790 24066 18842
rect 12126 18622 12178 18674
rect 14590 18622 14642 18674
rect 2718 18510 2770 18562
rect 5070 18510 5122 18562
rect 6078 18510 6130 18562
rect 8318 18510 8370 18562
rect 10558 18510 10610 18562
rect 13022 18510 13074 18562
rect 1598 18398 1650 18450
rect 2158 18398 2210 18450
rect 5518 18398 5570 18450
rect 7646 18398 7698 18450
rect 15822 18398 15874 18450
rect 16606 18398 16658 18450
rect 16830 18398 16882 18450
rect 17950 18398 18002 18450
rect 18510 18398 18562 18450
rect 19070 18398 19122 18450
rect 20974 18398 21026 18450
rect 21422 18398 21474 18450
rect 22654 18398 22706 18450
rect 23662 18398 23714 18450
rect 26014 18398 26066 18450
rect 26574 18398 26626 18450
rect 27358 18398 27410 18450
rect 8766 18286 8818 18338
rect 13358 18286 13410 18338
rect 17390 18286 17442 18338
rect 17838 18286 17890 18338
rect 18846 18286 18898 18338
rect 20638 18286 20690 18338
rect 22094 18286 22146 18338
rect 26910 18286 26962 18338
rect 3166 18174 3218 18226
rect 4286 18174 4338 18226
rect 6526 18174 6578 18226
rect 9886 18174 9938 18226
rect 11006 18174 11058 18226
rect 19518 18174 19570 18226
rect 19630 18174 19682 18226
rect 19742 18174 19794 18226
rect 21646 18174 21698 18226
rect 4466 18006 4518 18058
rect 4570 18006 4622 18058
rect 4674 18006 4726 18058
rect 24466 18006 24518 18058
rect 24570 18006 24622 18058
rect 24674 18006 24726 18058
rect 10446 17838 10498 17890
rect 12686 17838 12738 17890
rect 13806 17838 13858 17890
rect 16830 17838 16882 17890
rect 21534 17838 21586 17890
rect 27470 17838 27522 17890
rect 3726 17726 3778 17778
rect 5070 17726 5122 17778
rect 6078 17726 6130 17778
rect 6526 17726 6578 17778
rect 8878 17726 8930 17778
rect 9438 17726 9490 17778
rect 17278 17726 17330 17778
rect 17502 17726 17554 17778
rect 18846 17726 18898 17778
rect 22766 17726 22818 17778
rect 24558 17726 24610 17778
rect 26014 17726 26066 17778
rect 26574 17726 26626 17778
rect 26910 17726 26962 17778
rect 1822 17619 1874 17671
rect 2718 17614 2770 17666
rect 3278 17614 3330 17666
rect 3950 17614 4002 17666
rect 4286 17614 4338 17666
rect 5406 17614 5458 17666
rect 5966 17614 6018 17666
rect 7310 17614 7362 17666
rect 8206 17614 8258 17666
rect 9998 17614 10050 17666
rect 12126 17614 12178 17666
rect 15710 17614 15762 17666
rect 16718 17614 16770 17666
rect 18286 17614 18338 17666
rect 18622 17614 18674 17666
rect 19294 17614 19346 17666
rect 20078 17614 20130 17666
rect 20862 17614 20914 17666
rect 25118 17614 25170 17666
rect 4734 17502 4786 17554
rect 15262 17502 15314 17554
rect 17390 17502 17442 17554
rect 17838 17502 17890 17554
rect 23102 17502 23154 17554
rect 11566 17390 11618 17442
rect 3806 17222 3858 17274
rect 3910 17222 3962 17274
rect 4014 17222 4066 17274
rect 23806 17222 23858 17274
rect 23910 17222 23962 17274
rect 24014 17222 24066 17274
rect 2830 17054 2882 17106
rect 5966 17054 6018 17106
rect 18286 17054 18338 17106
rect 18510 17054 18562 17106
rect 19966 17054 20018 17106
rect 1262 16942 1314 16994
rect 3838 16942 3890 16994
rect 19630 16942 19682 16994
rect 26014 16942 26066 16994
rect 27022 16942 27074 16994
rect 3390 16830 3442 16882
rect 5070 16830 5122 16882
rect 8430 16830 8482 16882
rect 9326 16830 9378 16882
rect 9886 16830 9938 16882
rect 10558 16830 10610 16882
rect 11230 16830 11282 16882
rect 12014 16830 12066 16882
rect 15038 16830 15090 16882
rect 15486 16830 15538 16882
rect 16158 16830 16210 16882
rect 16942 16830 16994 16882
rect 17726 16830 17778 16882
rect 18734 16830 18786 16882
rect 19182 16830 19234 16882
rect 20974 16830 21026 16882
rect 23886 16830 23938 16882
rect 26574 16830 26626 16882
rect 27358 16830 27410 16882
rect 1598 16718 1650 16770
rect 8094 16718 8146 16770
rect 8990 16718 9042 16770
rect 14702 16718 14754 16770
rect 15710 16718 15762 16770
rect 18958 16718 19010 16770
rect 19070 16718 19122 16770
rect 19742 16718 19794 16770
rect 6862 16606 6914 16658
rect 9998 16606 10050 16658
rect 20750 16606 20802 16658
rect 20862 16606 20914 16658
rect 22206 16606 22258 16658
rect 23326 16606 23378 16658
rect 4466 16438 4518 16490
rect 4570 16438 4622 16490
rect 4674 16438 4726 16490
rect 24466 16438 24518 16490
rect 24570 16438 24622 16490
rect 24674 16438 24726 16490
rect 2942 16270 2994 16322
rect 4062 16270 4114 16322
rect 5182 16270 5234 16322
rect 8206 16270 8258 16322
rect 11678 16270 11730 16322
rect 12798 16270 12850 16322
rect 17054 16270 17106 16322
rect 17950 16270 18002 16322
rect 19966 16270 20018 16322
rect 27470 16270 27522 16322
rect 1822 16158 1874 16210
rect 5966 16158 6018 16210
rect 6974 16158 7026 16210
rect 10446 16158 10498 16210
rect 13806 16158 13858 16210
rect 16046 16158 16098 16210
rect 26014 16158 26066 16210
rect 26910 16158 26962 16210
rect 1374 16046 1426 16098
rect 3614 16046 3666 16098
rect 5854 16046 5906 16098
rect 6190 16046 6242 16098
rect 9214 16046 9266 16098
rect 9998 16046 10050 16098
rect 11118 16046 11170 16098
rect 13470 16046 13522 16098
rect 15598 16046 15650 16098
rect 16718 16046 16770 16098
rect 16942 16046 16994 16098
rect 17278 16046 17330 16098
rect 17838 16046 17890 16098
rect 18174 16046 18226 16098
rect 18286 16046 18338 16098
rect 18622 16046 18674 16098
rect 18958 16046 19010 16098
rect 19406 16046 19458 16098
rect 19742 16046 19794 16098
rect 20526 16046 20578 16098
rect 21198 16046 21250 16098
rect 22094 16046 22146 16098
rect 26574 16046 26626 16098
rect 6638 15934 6690 15986
rect 8878 15822 8930 15874
rect 9214 15822 9266 15874
rect 15038 15822 15090 15874
rect 17278 15822 17330 15874
rect 3806 15654 3858 15706
rect 3910 15654 3962 15706
rect 4014 15654 4066 15706
rect 23806 15654 23858 15706
rect 23910 15654 23962 15706
rect 24014 15654 24066 15706
rect 6750 15486 6802 15538
rect 9886 15486 9938 15538
rect 12126 15486 12178 15538
rect 18622 15486 18674 15538
rect 2158 15374 2210 15426
rect 4174 15374 4226 15426
rect 5182 15374 5234 15426
rect 10558 15374 10610 15426
rect 20638 15374 20690 15426
rect 26014 15374 26066 15426
rect 26910 15374 26962 15426
rect 1710 15262 1762 15314
rect 2606 15262 2658 15314
rect 7086 15262 7138 15314
rect 7534 15262 7586 15314
rect 7758 15262 7810 15314
rect 8318 15262 8370 15314
rect 14366 15262 14418 15314
rect 15150 15262 15202 15314
rect 15486 15262 15538 15314
rect 16158 15262 16210 15314
rect 16718 15262 16770 15314
rect 16942 15262 16994 15314
rect 17726 15262 17778 15314
rect 18398 15262 18450 15314
rect 18846 15262 18898 15314
rect 19742 15262 19794 15314
rect 20974 15262 21026 15314
rect 21422 15262 21474 15314
rect 22094 15262 22146 15314
rect 22766 15262 22818 15314
rect 23774 15262 23826 15314
rect 27358 15262 27410 15314
rect 3726 15150 3778 15202
rect 5630 15150 5682 15202
rect 7310 15150 7362 15202
rect 7646 15150 7698 15202
rect 8766 15150 8818 15202
rect 10894 15150 10946 15202
rect 14702 15150 14754 15202
rect 15710 15150 15762 15202
rect 19182 15150 19234 15202
rect 20078 15150 20130 15202
rect 14030 15038 14082 15090
rect 18398 15038 18450 15090
rect 19966 15038 20018 15090
rect 21646 15038 21698 15090
rect 26574 15038 26626 15090
rect 4466 14870 4518 14922
rect 4570 14870 4622 14922
rect 4674 14870 4726 14922
rect 24466 14870 24518 14922
rect 24570 14870 24622 14922
rect 24674 14870 24726 14922
rect 2158 14702 2210 14754
rect 3278 14702 3330 14754
rect 5742 14702 5794 14754
rect 9102 14702 9154 14754
rect 12462 14702 12514 14754
rect 13582 14702 13634 14754
rect 16830 14702 16882 14754
rect 16942 14702 16994 14754
rect 22542 14702 22594 14754
rect 27470 14702 27522 14754
rect 4174 14590 4226 14642
rect 6862 14590 6914 14642
rect 8878 14590 8930 14642
rect 9326 14590 9378 14642
rect 11342 14590 11394 14642
rect 14702 14590 14754 14642
rect 15710 14590 15762 14642
rect 17726 14590 17778 14642
rect 18734 14590 18786 14642
rect 22654 14590 22706 14642
rect 25118 14590 25170 14642
rect 26910 14590 26962 14642
rect 1710 14478 1762 14530
rect 3950 14478 4002 14530
rect 4286 14478 4338 14530
rect 5182 14478 5234 14530
rect 7758 14478 7810 14530
rect 7982 14478 8034 14530
rect 8206 14478 8258 14530
rect 8766 14478 8818 14530
rect 9886 14478 9938 14530
rect 10782 14478 10834 14530
rect 15150 14478 15202 14530
rect 16046 14478 16098 14530
rect 16718 14478 16770 14530
rect 18062 14478 18114 14530
rect 18510 14478 18562 14530
rect 19294 14478 19346 14530
rect 19742 14478 19794 14530
rect 20750 14478 20802 14530
rect 8094 14366 8146 14418
rect 10222 14366 10274 14418
rect 13134 14366 13186 14418
rect 22990 14366 23042 14418
rect 24782 14366 24834 14418
rect 4734 14254 4786 14306
rect 7310 14254 7362 14306
rect 7534 14254 7586 14306
rect 16158 14254 16210 14306
rect 21422 14254 21474 14306
rect 26350 14254 26402 14306
rect 3806 14086 3858 14138
rect 3910 14086 3962 14138
rect 4014 14086 4066 14138
rect 23806 14086 23858 14138
rect 23910 14086 23962 14138
rect 24014 14086 24066 14138
rect 5518 13918 5570 13970
rect 17390 13918 17442 13970
rect 19070 13918 19122 13970
rect 19294 13918 19346 13970
rect 4398 13806 4450 13858
rect 6974 13806 7026 13858
rect 8542 13806 8594 13858
rect 12798 13806 12850 13858
rect 19742 13806 19794 13858
rect 26014 13806 26066 13858
rect 27022 13806 27074 13858
rect 1822 13694 1874 13746
rect 3950 13694 4002 13746
rect 9326 13694 9378 13746
rect 9774 13694 9826 13746
rect 10670 13694 10722 13746
rect 11006 13694 11058 13746
rect 11230 13694 11282 13746
rect 12014 13694 12066 13746
rect 14142 13694 14194 13746
rect 14590 13694 14642 13746
rect 15710 13694 15762 13746
rect 16718 13694 16770 13746
rect 17726 13694 17778 13746
rect 18398 13694 18450 13746
rect 19518 13694 19570 13746
rect 21422 13694 21474 13746
rect 22990 13694 23042 13746
rect 25230 13694 25282 13746
rect 26574 13694 26626 13746
rect 27358 13694 27410 13746
rect 3390 13582 3442 13634
rect 4958 13582 5010 13634
rect 7422 13582 7474 13634
rect 8990 13582 9042 13634
rect 9998 13582 10050 13634
rect 12910 13582 12962 13634
rect 13134 13582 13186 13634
rect 13694 13582 13746 13634
rect 14702 13582 14754 13634
rect 15150 13582 15202 13634
rect 18286 13582 18338 13634
rect 19966 13582 20018 13634
rect 20638 13582 20690 13634
rect 20862 13582 20914 13634
rect 24782 13582 24834 13634
rect 2270 13470 2322 13522
rect 19742 13470 19794 13522
rect 20750 13470 20802 13522
rect 22542 13470 22594 13522
rect 23662 13470 23714 13522
rect 4466 13302 4518 13354
rect 4570 13302 4622 13354
rect 4674 13302 4726 13354
rect 24466 13302 24518 13354
rect 24570 13302 24622 13354
rect 24674 13302 24726 13354
rect 3614 13134 3666 13186
rect 5742 13134 5794 13186
rect 7870 13134 7922 13186
rect 13806 13134 13858 13186
rect 16046 13134 16098 13186
rect 25118 13134 25170 13186
rect 27470 13134 27522 13186
rect 1486 13022 1538 13074
rect 3166 13022 3218 13074
rect 3502 13022 3554 13074
rect 4622 13022 4674 13074
rect 10334 13022 10386 13074
rect 12686 13022 12738 13074
rect 14926 13022 14978 13074
rect 17838 13022 17890 13074
rect 18734 13022 18786 13074
rect 19182 13022 19234 13074
rect 20190 13022 20242 13074
rect 24558 13022 24610 13074
rect 2046 12910 2098 12962
rect 2606 12910 2658 12962
rect 4174 12910 4226 12962
rect 7422 12910 7474 12962
rect 7982 12910 8034 12962
rect 8878 12910 8930 12962
rect 14366 12910 14418 12962
rect 17950 12910 18002 12962
rect 18398 12910 18450 12962
rect 19630 12910 19682 12962
rect 19966 12910 20018 12962
rect 20862 12910 20914 12962
rect 21422 12910 21474 12962
rect 22206 12910 22258 12962
rect 25006 12910 25058 12962
rect 26574 12910 26626 12962
rect 6414 12798 6466 12850
rect 9998 12798 10050 12850
rect 12238 12798 12290 12850
rect 26014 12798 26066 12850
rect 27022 12798 27074 12850
rect 7870 12686 7922 12738
rect 8206 12686 8258 12738
rect 8878 12686 8930 12738
rect 9214 12686 9266 12738
rect 11566 12686 11618 12738
rect 16830 12686 16882 12738
rect 17166 12686 17218 12738
rect 18398 12686 18450 12738
rect 3806 12518 3858 12570
rect 3910 12518 3962 12570
rect 4014 12518 4066 12570
rect 23806 12518 23858 12570
rect 23910 12518 23962 12570
rect 24014 12518 24066 12570
rect 3614 12350 3666 12402
rect 13022 12350 13074 12402
rect 17502 12350 17554 12402
rect 18286 12350 18338 12402
rect 21534 12350 21586 12402
rect 5294 12238 5346 12290
rect 9438 12238 9490 12290
rect 11006 12238 11058 12290
rect 12014 12238 12066 12290
rect 20750 12238 20802 12290
rect 2046 12126 2098 12178
rect 6078 12126 6130 12178
rect 8766 12126 8818 12178
rect 11566 12126 11618 12178
rect 14030 12126 14082 12178
rect 14814 12126 14866 12178
rect 16494 12126 16546 12178
rect 16942 12126 16994 12178
rect 17166 12126 17218 12178
rect 17614 12126 17666 12178
rect 18062 12126 18114 12178
rect 18510 12126 18562 12178
rect 18958 12126 19010 12178
rect 19518 12126 19570 12178
rect 19630 12126 19682 12178
rect 19966 12126 20018 12178
rect 20862 12126 20914 12178
rect 21646 12126 21698 12178
rect 24222 12126 24274 12178
rect 26014 12126 26066 12178
rect 27358 12126 27410 12178
rect 2494 12014 2546 12066
rect 6526 12014 6578 12066
rect 7310 12014 7362 12066
rect 8542 12014 8594 12066
rect 8654 12014 8706 12066
rect 9774 12014 9826 12066
rect 15262 12014 15314 12066
rect 26910 12014 26962 12066
rect 8094 11902 8146 11954
rect 17726 11902 17778 11954
rect 18734 11902 18786 11954
rect 18846 11902 18898 11954
rect 19406 11902 19458 11954
rect 20638 11902 20690 11954
rect 21086 11902 21138 11954
rect 22542 11902 22594 11954
rect 23662 11902 23714 11954
rect 26574 11902 26626 11954
rect 4466 11734 4518 11786
rect 4570 11734 4622 11786
rect 4674 11734 4726 11786
rect 24466 11734 24518 11786
rect 24570 11734 24622 11786
rect 24674 11734 24726 11786
rect 1598 11566 1650 11618
rect 2718 11566 2770 11618
rect 7534 11566 7586 11618
rect 8318 11566 8370 11618
rect 9774 11566 9826 11618
rect 11454 11566 11506 11618
rect 14142 11566 14194 11618
rect 15598 11566 15650 11618
rect 18734 11566 18786 11618
rect 23214 11566 23266 11618
rect 27470 11566 27522 11618
rect 5406 11454 5458 11506
rect 6638 11454 6690 11506
rect 7086 11454 7138 11506
rect 8206 11454 8258 11506
rect 9886 11454 9938 11506
rect 11006 11454 11058 11506
rect 11118 11454 11170 11506
rect 13022 11454 13074 11506
rect 16718 11454 16770 11506
rect 17054 11454 17106 11506
rect 19182 11454 19234 11506
rect 23774 11454 23826 11506
rect 26014 11454 26066 11506
rect 26910 11454 26962 11506
rect 3166 11342 3218 11394
rect 3838 11342 3890 11394
rect 7310 11342 7362 11394
rect 7758 11342 7810 11394
rect 8990 11342 9042 11394
rect 9102 11342 9154 11394
rect 9326 11342 9378 11394
rect 10782 11342 10834 11394
rect 11678 11342 11730 11394
rect 12014 11342 12066 11394
rect 12462 11342 12514 11394
rect 18062 11342 18114 11394
rect 18510 11342 18562 11394
rect 19854 11342 19906 11394
rect 20862 11342 20914 11394
rect 26574 11342 26626 11394
rect 4286 11230 4338 11282
rect 5070 11230 5122 11282
rect 11566 11230 11618 11282
rect 17726 11230 17778 11282
rect 7646 11118 7698 11170
rect 9438 11118 9490 11170
rect 15374 11118 15426 11170
rect 15710 11118 15762 11170
rect 3806 10950 3858 11002
rect 3910 10950 3962 11002
rect 4014 10950 4066 11002
rect 23806 10950 23858 11002
rect 23910 10950 23962 11002
rect 24014 10950 24066 11002
rect 3614 10782 3666 10834
rect 7198 10782 7250 10834
rect 12014 10782 12066 10834
rect 18286 10782 18338 10834
rect 5182 10670 5234 10722
rect 7982 10670 8034 10722
rect 13246 10670 13298 10722
rect 14702 10670 14754 10722
rect 17726 10670 17778 10722
rect 26014 10670 26066 10722
rect 27022 10670 27074 10722
rect 2046 10558 2098 10610
rect 7422 10558 7474 10610
rect 7758 10558 7810 10610
rect 7870 10558 7922 10610
rect 8766 10558 8818 10610
rect 10894 10558 10946 10610
rect 11454 10558 11506 10610
rect 11902 10558 11954 10610
rect 12126 10558 12178 10610
rect 12798 10558 12850 10610
rect 13022 10558 13074 10610
rect 13470 10558 13522 10610
rect 16606 10558 16658 10610
rect 17502 10558 17554 10610
rect 19854 10558 19906 10610
rect 27358 10558 27410 10610
rect 5630 10446 5682 10498
rect 6750 10446 6802 10498
rect 9326 10446 9378 10498
rect 9662 10446 9714 10498
rect 10110 10446 10162 10498
rect 10670 10446 10722 10498
rect 11118 10446 11170 10498
rect 11678 10446 11730 10498
rect 15038 10446 15090 10498
rect 17838 10446 17890 10498
rect 19406 10446 19458 10498
rect 2494 10334 2546 10386
rect 8094 10334 8146 10386
rect 9550 10334 9602 10386
rect 9886 10334 9938 10386
rect 11230 10334 11282 10386
rect 12238 10334 12290 10386
rect 13582 10334 13634 10386
rect 13694 10334 13746 10386
rect 16270 10334 16322 10386
rect 16942 10334 16994 10386
rect 17166 10334 17218 10386
rect 17278 10334 17330 10386
rect 26574 10334 26626 10386
rect 4466 10166 4518 10218
rect 4570 10166 4622 10218
rect 4674 10166 4726 10218
rect 24466 10166 24518 10218
rect 24570 10166 24622 10218
rect 24674 10166 24726 10218
rect 6526 9998 6578 10050
rect 7422 9998 7474 10050
rect 12686 9998 12738 10050
rect 13918 9998 13970 10050
rect 15262 9998 15314 10050
rect 16046 9998 16098 10050
rect 18958 9998 19010 10050
rect 27470 9998 27522 10050
rect 2270 9886 2322 9938
rect 5294 9886 5346 9938
rect 7086 9886 7138 9938
rect 9102 9886 9154 9938
rect 10110 9886 10162 9938
rect 13134 9886 13186 9938
rect 15150 9886 15202 9938
rect 17166 9886 17218 9938
rect 19406 9886 19458 9938
rect 26910 9886 26962 9938
rect 3838 9774 3890 9826
rect 4958 9774 5010 9826
rect 7310 9774 7362 9826
rect 7534 9774 7586 9826
rect 7870 9774 7922 9826
rect 9550 9774 9602 9826
rect 9998 9774 10050 9826
rect 10782 9774 10834 9826
rect 11342 9774 11394 9826
rect 12238 9774 12290 9826
rect 13246 9774 13298 9826
rect 13470 9774 13522 9826
rect 13806 9774 13858 9826
rect 14926 9774 14978 9826
rect 15710 9774 15762 9826
rect 16158 9774 16210 9826
rect 16606 9774 16658 9826
rect 17054 9774 17106 9826
rect 17278 9774 17330 9826
rect 18398 9774 18450 9826
rect 18846 9774 18898 9826
rect 20078 9774 20130 9826
rect 21086 9774 21138 9826
rect 25678 9774 25730 9826
rect 26574 9774 26626 9826
rect 1262 9662 1314 9714
rect 2830 9662 2882 9714
rect 17950 9662 18002 9714
rect 25118 9662 25170 9714
rect 26014 9662 26066 9714
rect 14030 9550 14082 9602
rect 14254 9550 14306 9602
rect 15486 9550 15538 9602
rect 3806 9382 3858 9434
rect 3910 9382 3962 9434
rect 4014 9382 4066 9434
rect 23806 9382 23858 9434
rect 23910 9382 23962 9434
rect 24014 9382 24066 9434
rect 1262 9214 1314 9266
rect 9662 9214 9714 9266
rect 13806 9214 13858 9266
rect 16494 9214 16546 9266
rect 17054 9214 17106 9266
rect 26462 9214 26514 9266
rect 3054 9102 3106 9154
rect 5518 9102 5570 9154
rect 6414 9102 6466 9154
rect 7422 9102 7474 9154
rect 18622 9102 18674 9154
rect 25342 9102 25394 9154
rect 2270 8990 2322 9042
rect 3838 8990 3890 9042
rect 5070 8990 5122 9042
rect 5854 8990 5906 9042
rect 6974 8990 7026 9042
rect 7310 8990 7362 9042
rect 7534 8990 7586 9042
rect 8094 8990 8146 9042
rect 10446 8990 10498 9042
rect 12798 8990 12850 9042
rect 14814 8990 14866 9042
rect 27246 8990 27298 9042
rect 10894 8878 10946 8930
rect 12126 8878 12178 8930
rect 18174 8878 18226 8930
rect 8542 8766 8594 8818
rect 15374 8766 15426 8818
rect 25902 8766 25954 8818
rect 4466 8598 4518 8650
rect 4570 8598 4622 8650
rect 4674 8598 4726 8650
rect 24466 8598 24518 8650
rect 24570 8598 24622 8650
rect 24674 8598 24726 8650
rect 12238 8430 12290 8482
rect 3054 8318 3106 8370
rect 6190 8318 6242 8370
rect 7198 8318 7250 8370
rect 8094 8318 8146 8370
rect 8206 8318 8258 8370
rect 11118 8318 11170 8370
rect 13246 8318 13298 8370
rect 14926 8318 14978 8370
rect 15598 8318 15650 8370
rect 15710 8318 15762 8370
rect 17614 8318 17666 8370
rect 19518 8318 19570 8370
rect 20526 8318 20578 8370
rect 2270 8206 2322 8258
rect 3614 8206 3666 8258
rect 6638 8206 6690 8258
rect 10558 8206 10610 8258
rect 15374 8206 15426 8258
rect 16942 8206 16994 8258
rect 17278 8206 17330 8258
rect 17390 8206 17442 8258
rect 19966 8206 20018 8258
rect 20302 8206 20354 8258
rect 20974 8206 21026 8258
rect 21646 8206 21698 8258
rect 22542 8206 22594 8258
rect 27358 8206 27410 8258
rect 7758 8094 7810 8146
rect 12910 8094 12962 8146
rect 17502 8094 17554 8146
rect 26462 8094 26514 8146
rect 1262 7982 1314 8034
rect 5070 7982 5122 8034
rect 8206 7982 8258 8034
rect 14478 7982 14530 8034
rect 15038 7982 15090 8034
rect 16158 7982 16210 8034
rect 16718 7982 16770 8034
rect 3806 7814 3858 7866
rect 3910 7814 3962 7866
rect 4014 7814 4066 7866
rect 23806 7814 23858 7866
rect 23910 7814 23962 7866
rect 24014 7814 24066 7866
rect 10894 7646 10946 7698
rect 12238 7646 12290 7698
rect 16606 7646 16658 7698
rect 16718 7646 16770 7698
rect 1486 7534 1538 7586
rect 2942 7534 2994 7586
rect 5518 7534 5570 7586
rect 7310 7534 7362 7586
rect 9326 7534 9378 7586
rect 17054 7534 17106 7586
rect 26014 7534 26066 7586
rect 27022 7534 27074 7586
rect 2270 7422 2322 7474
rect 3838 7422 3890 7474
rect 5070 7422 5122 7474
rect 6862 7422 6914 7474
rect 12126 7422 12178 7474
rect 12910 7422 12962 7474
rect 14590 7422 14642 7474
rect 15934 7422 15986 7474
rect 16158 7422 16210 7474
rect 16382 7422 16434 7474
rect 17390 7422 17442 7474
rect 9774 7310 9826 7362
rect 13358 7310 13410 7362
rect 15598 7310 15650 7362
rect 27470 7310 27522 7362
rect 15710 7198 15762 7250
rect 26574 7198 26626 7250
rect 4466 7030 4518 7082
rect 4570 7030 4622 7082
rect 4674 7030 4726 7082
rect 24466 7030 24518 7082
rect 24570 7030 24622 7082
rect 24674 7030 24726 7082
rect 13918 6862 13970 6914
rect 27470 6862 27522 6914
rect 12686 6750 12738 6802
rect 26014 6750 26066 6802
rect 26910 6750 26962 6802
rect 2046 6638 2098 6690
rect 3838 6638 3890 6690
rect 9662 6638 9714 6690
rect 10110 6638 10162 6690
rect 11006 6638 11058 6690
rect 11566 6638 11618 6690
rect 12350 6638 12402 6690
rect 26574 6638 26626 6690
rect 1374 6526 1426 6578
rect 2830 6414 2882 6466
rect 3806 6246 3858 6298
rect 3910 6246 3962 6298
rect 4014 6246 4066 6298
rect 23806 6246 23858 6298
rect 23910 6246 23962 6298
rect 24014 6246 24066 6298
rect 7758 6078 7810 6130
rect 26462 6078 26514 6130
rect 1598 5966 1650 6018
rect 9326 5966 9378 6018
rect 12014 5966 12066 6018
rect 13806 5966 13858 6018
rect 25342 5966 25394 6018
rect 2158 5854 2210 5906
rect 2606 5854 2658 5906
rect 14254 5854 14306 5906
rect 14702 5854 14754 5906
rect 16046 5854 16098 5906
rect 16942 5854 16994 5906
rect 27358 5854 27410 5906
rect 3166 5742 3218 5794
rect 15262 5742 15314 5794
rect 8878 5630 8930 5682
rect 11566 5630 11618 5682
rect 14814 5630 14866 5682
rect 25902 5630 25954 5682
rect 4466 5462 4518 5514
rect 4570 5462 4622 5514
rect 4674 5462 4726 5514
rect 24466 5462 24518 5514
rect 24570 5462 24622 5514
rect 24674 5462 24726 5514
rect 2606 5294 2658 5346
rect 7758 5294 7810 5346
rect 13806 5294 13858 5346
rect 14926 5294 14978 5346
rect 15374 5294 15426 5346
rect 1486 5182 1538 5234
rect 3166 5182 3218 5234
rect 3502 5182 3554 5234
rect 8318 5182 8370 5234
rect 12798 5182 12850 5234
rect 15934 5182 15986 5234
rect 26686 5182 26738 5234
rect 2046 5070 2098 5122
rect 4062 5070 4114 5122
rect 12350 5070 12402 5122
rect 13358 5070 13410 5122
rect 27470 5070 27522 5122
rect 3806 4678 3858 4730
rect 3910 4678 3962 4730
rect 4014 4678 4066 4730
rect 23806 4678 23858 4730
rect 23910 4678 23962 4730
rect 24014 4678 24066 4730
rect 27470 4286 27522 4338
rect 1486 4174 1538 4226
rect 2270 4174 2322 4226
rect 26910 4174 26962 4226
rect 4466 3894 4518 3946
rect 4570 3894 4622 3946
rect 4674 3894 4726 3946
rect 24466 3894 24518 3946
rect 24570 3894 24622 3946
rect 24674 3894 24726 3946
rect 27470 3726 27522 3778
rect 26910 3614 26962 3666
rect 2270 3502 2322 3554
rect 26574 3502 26626 3554
rect 26126 3390 26178 3442
rect 1262 3278 1314 3330
rect 3806 3110 3858 3162
rect 3910 3110 3962 3162
rect 4014 3110 4066 3162
rect 23806 3110 23858 3162
rect 23910 3110 23962 3162
rect 24014 3110 24066 3162
rect 1486 2830 1538 2882
rect 25230 2830 25282 2882
rect 26126 2830 26178 2882
rect 27022 2830 27074 2882
rect 1038 2718 1090 2770
rect 27470 2718 27522 2770
rect 25678 2494 25730 2546
rect 26574 2494 26626 2546
rect 4466 2326 4518 2378
rect 4570 2326 4622 2378
rect 4674 2326 4726 2378
rect 24466 2326 24518 2378
rect 24570 2326 24622 2378
rect 24674 2326 24726 2378
rect 1038 2158 1090 2210
rect 1598 2046 1650 2098
rect 11454 2046 11506 2098
rect 13246 2046 13298 2098
rect 27470 2046 27522 2098
rect 12014 1934 12066 1986
rect 13806 1934 13858 1986
rect 25566 1934 25618 1986
rect 26014 1934 26066 1986
rect 26910 1934 26962 1986
rect 25230 1822 25282 1874
rect 26462 1822 26514 1874
rect 3806 1542 3858 1594
rect 3910 1542 3962 1594
rect 4014 1542 4066 1594
rect 23806 1542 23858 1594
rect 23910 1542 23962 1594
rect 24014 1542 24066 1594
rect 7982 1262 8034 1314
rect 24894 1262 24946 1314
rect 25678 1262 25730 1314
rect 26574 1262 26626 1314
rect 27134 1150 27186 1202
rect 7534 926 7586 978
rect 25342 926 25394 978
rect 26238 926 26290 978
rect 4466 758 4518 810
rect 4570 758 4622 810
rect 4674 758 4726 810
rect 24466 758 24518 810
rect 24570 758 24622 810
rect 24674 758 24726 810
<< metal2 >>
rect 672 57344 784 57456
rect 2016 57344 2128 57456
rect 3360 57344 3472 57456
rect 4704 57344 4816 57456
rect 6048 57344 6160 57456
rect 7392 57344 7504 57456
rect 8736 57344 8848 57456
rect 10080 57344 10192 57456
rect 11424 57344 11536 57456
rect 12768 57344 12880 57456
rect 14112 57344 14224 57456
rect 15456 57344 15568 57456
rect 16800 57344 16912 57456
rect 18144 57344 18256 57456
rect 19488 57344 19600 57456
rect 19852 57372 20356 57428
rect 700 55972 756 57344
rect 1036 55972 1092 55982
rect 700 55970 1092 55972
rect 700 55918 1038 55970
rect 1090 55918 1092 55970
rect 700 55916 1092 55918
rect 1036 55906 1092 55916
rect 1372 55858 1428 55870
rect 1372 55806 1374 55858
rect 1426 55806 1428 55858
rect 1036 55298 1092 55310
rect 1036 55246 1038 55298
rect 1090 55246 1092 55298
rect 1036 55188 1092 55246
rect 1372 55300 1428 55806
rect 2044 55468 2100 57344
rect 3388 56308 3444 57344
rect 4732 56644 4788 57344
rect 4732 56588 5236 56644
rect 3804 56476 4068 56486
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 3804 56410 4068 56420
rect 3612 56308 3668 56318
rect 3388 56306 3668 56308
rect 3388 56254 3614 56306
rect 3666 56254 3668 56306
rect 3388 56252 3668 56254
rect 3612 56242 3668 56252
rect 5180 56306 5236 56588
rect 5180 56254 5182 56306
rect 5234 56254 5236 56306
rect 5180 56242 5236 56254
rect 3052 55972 3108 55982
rect 3052 55878 3108 55916
rect 4464 55692 4728 55702
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4464 55626 4728 55636
rect 2044 55412 2548 55468
rect 1372 55234 1428 55244
rect 1036 55122 1092 55132
rect 1484 55186 1540 55198
rect 1484 55134 1486 55186
rect 1538 55134 1540 55186
rect 1484 54852 1540 55134
rect 2492 55186 2548 55412
rect 2492 55134 2494 55186
rect 2546 55134 2548 55186
rect 2492 55122 2548 55134
rect 3500 55298 3556 55310
rect 3500 55246 3502 55298
rect 3554 55246 3556 55298
rect 364 54796 1540 54852
rect 364 50428 420 54796
rect 1484 54628 1540 54638
rect 1148 54626 1540 54628
rect 1148 54574 1486 54626
rect 1538 54574 1540 54626
rect 1148 54572 1540 54574
rect 1036 54292 1092 54302
rect 1036 54198 1092 54236
rect 1036 53730 1092 53742
rect 1036 53678 1038 53730
rect 1090 53678 1092 53730
rect 1036 53396 1092 53678
rect 1036 53330 1092 53340
rect 1036 52722 1092 52734
rect 1036 52670 1038 52722
rect 1090 52670 1092 52722
rect 1036 52500 1092 52670
rect 1036 52434 1092 52444
rect 1036 52162 1092 52174
rect 1036 52110 1038 52162
rect 1090 52110 1092 52162
rect 1036 51604 1092 52110
rect 1036 51538 1092 51548
rect 1036 51156 1092 51166
rect 924 51154 1092 51156
rect 924 51102 1038 51154
rect 1090 51102 1092 51154
rect 924 51100 1092 51102
rect 924 50708 980 51100
rect 1036 51090 1092 51100
rect 924 50642 980 50652
rect 28 50372 420 50428
rect 1036 50594 1092 50606
rect 1036 50542 1038 50594
rect 1090 50542 1092 50594
rect 28 38668 84 50372
rect 1036 49812 1092 50542
rect 1036 49746 1092 49756
rect 1036 49026 1092 49038
rect 1036 48974 1038 49026
rect 1090 48974 1092 49026
rect 1036 48916 1092 48974
rect 1036 48850 1092 48860
rect 1148 48468 1204 54572
rect 1484 54562 1540 54572
rect 1596 53618 1652 53630
rect 1596 53566 1598 53618
rect 1650 53566 1652 53618
rect 1596 53060 1652 53566
rect 1596 53004 1764 53060
rect 1596 52836 1652 52846
rect 1148 48402 1204 48412
rect 1260 52834 1652 52836
rect 1260 52782 1598 52834
rect 1650 52782 1652 52834
rect 1260 52780 1652 52782
rect 812 48132 868 48142
rect 812 43652 868 48076
rect 1036 48020 1092 48030
rect 1036 47926 1092 47964
rect 1036 47458 1092 47470
rect 1036 47406 1038 47458
rect 1090 47406 1092 47458
rect 1036 47124 1092 47406
rect 1036 47058 1092 47068
rect 1036 46452 1092 46462
rect 924 46450 1092 46452
rect 924 46398 1038 46450
rect 1090 46398 1092 46450
rect 924 46396 1092 46398
rect 924 45332 980 46396
rect 1036 46386 1092 46396
rect 924 45266 980 45276
rect 1148 45890 1204 45902
rect 1148 45838 1150 45890
rect 1202 45838 1204 45890
rect 1036 44884 1092 44894
rect 812 43586 868 43596
rect 924 44882 1092 44884
rect 924 44830 1038 44882
rect 1090 44830 1092 44882
rect 924 44828 1092 44830
rect 924 43540 980 44828
rect 1036 44818 1092 44828
rect 1148 44436 1204 45838
rect 1148 44370 1204 44380
rect 1036 44322 1092 44334
rect 1036 44270 1038 44322
rect 1090 44270 1092 44322
rect 1036 43540 1092 44270
rect 1036 43484 1204 43540
rect 924 43474 980 43484
rect 1036 43316 1092 43326
rect 364 43314 1092 43316
rect 364 43262 1038 43314
rect 1090 43262 1092 43314
rect 364 43260 1092 43262
rect 252 41076 308 41086
rect 28 38612 196 38668
rect 140 30772 196 38612
rect 252 35028 308 41020
rect 364 39060 420 43260
rect 1036 43250 1092 43260
rect 1036 42756 1092 42766
rect 364 38994 420 39004
rect 476 42754 1092 42756
rect 476 42702 1038 42754
rect 1090 42702 1092 42754
rect 476 42700 1092 42702
rect 476 37268 532 42700
rect 1036 42690 1092 42700
rect 1148 42644 1204 43484
rect 1148 42578 1204 42588
rect 1036 41748 1092 41758
rect 476 37202 532 37212
rect 588 41746 1092 41748
rect 588 41694 1038 41746
rect 1090 41694 1092 41746
rect 588 41692 1092 41694
rect 364 36820 420 36830
rect 364 35476 420 36764
rect 588 36372 644 41692
rect 1036 41682 1092 41692
rect 1036 41188 1092 41198
rect 812 41186 1092 41188
rect 812 41134 1038 41186
rect 1090 41134 1092 41186
rect 812 41132 1092 41134
rect 588 36306 644 36316
rect 700 40292 756 40302
rect 364 35410 420 35420
rect 588 35812 644 35822
rect 252 34972 532 35028
rect 140 30706 196 30716
rect 364 30772 420 30782
rect 140 27412 196 27422
rect 140 27076 196 27356
rect 140 27010 196 27020
rect 364 22148 420 30716
rect 476 26404 532 34972
rect 588 33348 644 35756
rect 588 33282 644 33292
rect 476 26338 532 26348
rect 588 33124 644 33134
rect 364 22082 420 22092
rect 364 20692 420 20702
rect 364 2884 420 20636
rect 588 13188 644 33068
rect 700 26908 756 40236
rect 812 36820 868 41132
rect 1036 41122 1092 41132
rect 1148 40402 1204 40414
rect 1148 40350 1150 40402
rect 1202 40350 1204 40402
rect 812 36754 868 36764
rect 1036 38610 1092 38622
rect 1036 38558 1038 38610
rect 1090 38558 1092 38610
rect 1036 36148 1092 38558
rect 812 36092 1092 36148
rect 812 33684 868 36092
rect 1148 35700 1204 40350
rect 1036 35644 1204 35700
rect 1260 35700 1316 52780
rect 1596 52770 1652 52780
rect 1708 52612 1764 53004
rect 1484 52556 1764 52612
rect 1484 46340 1540 52556
rect 1596 52164 1652 52174
rect 1596 52070 1652 52108
rect 1596 51268 1652 51278
rect 1596 51174 1652 51212
rect 1596 50484 1652 50494
rect 1596 50390 1652 50428
rect 2380 50484 2436 50494
rect 1596 48916 1652 48926
rect 1596 48914 1764 48916
rect 1596 48862 1598 48914
rect 1650 48862 1764 48914
rect 1596 48860 1764 48862
rect 1596 48850 1652 48860
rect 1596 48132 1652 48142
rect 1596 48038 1652 48076
rect 1596 46564 1652 46574
rect 1596 46470 1652 46508
rect 1484 46274 1540 46284
rect 1596 45780 1652 45790
rect 1596 45686 1652 45724
rect 1596 44994 1652 45006
rect 1596 44942 1598 44994
rect 1650 44942 1652 44994
rect 1596 44436 1652 44942
rect 1596 44370 1652 44380
rect 1596 44210 1652 44222
rect 1596 44158 1598 44210
rect 1650 44158 1652 44210
rect 1596 43764 1652 44158
rect 1596 43698 1652 43708
rect 1596 43428 1652 43438
rect 1596 43334 1652 43372
rect 1708 42868 1764 48860
rect 2044 47234 2100 47246
rect 2044 47182 2046 47234
rect 2098 47182 2100 47234
rect 1932 46450 1988 46462
rect 1932 46398 1934 46450
rect 1986 46398 1988 46450
rect 1932 46228 1988 46398
rect 1932 46162 1988 46172
rect 1708 42802 1764 42812
rect 1932 42756 1988 42766
rect 1820 42754 1988 42756
rect 1820 42702 1934 42754
rect 1986 42702 1988 42754
rect 1820 42700 1988 42702
rect 1596 42642 1652 42654
rect 1596 42590 1598 42642
rect 1650 42590 1652 42642
rect 1596 42196 1652 42590
rect 1596 42130 1652 42140
rect 1708 42644 1764 42654
rect 1372 42084 1428 42094
rect 1372 40628 1428 42028
rect 1596 41860 1652 41870
rect 1596 41766 1652 41804
rect 1596 41076 1652 41086
rect 1596 40982 1652 41020
rect 1708 40628 1764 42588
rect 1820 40852 1876 42700
rect 1932 42690 1988 42700
rect 2044 42196 2100 47182
rect 2380 42980 2436 50428
rect 2492 46564 2548 46574
rect 2492 46562 2996 46564
rect 2492 46510 2494 46562
rect 2546 46510 2996 46562
rect 2492 46508 2996 46510
rect 2492 46498 2548 46508
rect 2380 42914 2436 42924
rect 2604 43428 2660 43438
rect 2380 42644 2436 42654
rect 2380 42550 2436 42588
rect 2044 42130 2100 42140
rect 2492 41860 2548 41870
rect 2044 41858 2548 41860
rect 2044 41806 2494 41858
rect 2546 41806 2548 41858
rect 2044 41804 2548 41806
rect 1932 41748 1988 41758
rect 1932 41654 1988 41692
rect 2044 41412 2100 41804
rect 2492 41794 2548 41804
rect 1820 40786 1876 40796
rect 1932 41356 2100 41412
rect 2268 41636 2324 41646
rect 1708 40572 1876 40628
rect 1372 40562 1428 40572
rect 1596 40292 1652 40302
rect 1596 40198 1652 40236
rect 1708 39618 1764 39630
rect 1708 39566 1710 39618
rect 1762 39566 1764 39618
rect 1596 38948 1652 38958
rect 1596 38854 1652 38892
rect 1708 38612 1764 39566
rect 1708 38546 1764 38556
rect 1820 38162 1876 40572
rect 1820 38110 1822 38162
rect 1874 38110 1876 38162
rect 1820 38052 1876 38110
rect 1820 37986 1876 37996
rect 1932 40402 1988 41356
rect 1932 40350 1934 40402
rect 1986 40350 1988 40402
rect 1372 37938 1428 37950
rect 1372 37886 1374 37938
rect 1426 37886 1428 37938
rect 1372 35812 1428 37886
rect 1932 37940 1988 40350
rect 2044 41186 2100 41198
rect 2044 41134 2046 41186
rect 2098 41134 2100 41186
rect 2044 39956 2100 41134
rect 2044 39890 2100 39900
rect 2156 40292 2212 40302
rect 2156 39730 2212 40236
rect 2156 39678 2158 39730
rect 2210 39678 2212 39730
rect 2156 39666 2212 39678
rect 2268 39844 2324 41580
rect 2604 41300 2660 43372
rect 2156 38834 2212 38846
rect 2156 38782 2158 38834
rect 2210 38782 2212 38834
rect 2156 38612 2212 38782
rect 2156 38546 2212 38556
rect 1932 37874 1988 37884
rect 2268 37492 2324 39788
rect 1932 37436 2324 37492
rect 2380 41244 2660 41300
rect 1708 37378 1764 37390
rect 1708 37326 1710 37378
rect 1762 37326 1764 37378
rect 1708 37156 1764 37326
rect 1708 37090 1764 37100
rect 1372 35746 1428 35756
rect 1708 36932 1764 36942
rect 1036 35140 1092 35644
rect 1260 35634 1316 35644
rect 1148 35474 1204 35486
rect 1148 35422 1150 35474
rect 1202 35422 1204 35474
rect 1148 35364 1204 35422
rect 1148 35308 1428 35364
rect 1372 35140 1428 35308
rect 1036 35084 1204 35140
rect 1036 34916 1092 34926
rect 812 33618 868 33628
rect 924 34914 1092 34916
rect 924 34862 1038 34914
rect 1090 34862 1092 34914
rect 924 34860 1092 34862
rect 924 31892 980 34860
rect 1036 34850 1092 34860
rect 1148 34580 1204 35084
rect 1372 35074 1428 35084
rect 1148 34514 1204 34524
rect 1260 35028 1316 35038
rect 1148 34018 1204 34030
rect 1148 33966 1150 34018
rect 1202 33966 1204 34018
rect 1148 33572 1204 33966
rect 1260 33684 1316 34972
rect 1596 34804 1652 34814
rect 1596 34710 1652 34748
rect 1596 34468 1652 34478
rect 1484 34132 1540 34142
rect 1484 34038 1540 34076
rect 1260 33618 1316 33628
rect 1484 33684 1540 33694
rect 1148 33506 1204 33516
rect 924 31826 980 31836
rect 1036 33346 1092 33358
rect 1036 33294 1038 33346
rect 1090 33294 1092 33346
rect 1036 30996 1092 33294
rect 1148 33348 1204 33358
rect 1148 32562 1204 33292
rect 1148 32510 1150 32562
rect 1202 32510 1204 32562
rect 1148 32340 1204 32510
rect 1148 31780 1204 32284
rect 1148 31714 1204 31724
rect 1260 32452 1316 32462
rect 1036 30930 1092 30940
rect 1036 30770 1092 30782
rect 1036 30718 1038 30770
rect 1090 30718 1092 30770
rect 1036 30100 1092 30718
rect 1260 30324 1316 32396
rect 1484 30660 1540 33628
rect 1596 33460 1652 34412
rect 1708 33684 1764 36876
rect 1932 35252 1988 37436
rect 1932 35186 1988 35196
rect 2044 37266 2100 37278
rect 2044 37214 2046 37266
rect 2098 37214 2100 37266
rect 1932 34916 1988 34926
rect 1708 33618 1764 33628
rect 1820 34914 1988 34916
rect 1820 34862 1934 34914
rect 1986 34862 1988 34914
rect 1820 34860 1988 34862
rect 1596 33404 1764 33460
rect 1596 33236 1652 33246
rect 1596 33142 1652 33180
rect 1708 33012 1764 33404
rect 1596 32956 1764 33012
rect 1596 31106 1652 32956
rect 1820 32788 1876 34860
rect 1932 34850 1988 34860
rect 1932 34130 1988 34142
rect 1932 34078 1934 34130
rect 1986 34078 1988 34130
rect 1932 33908 1988 34078
rect 2044 34020 2100 37214
rect 2268 36708 2324 36718
rect 2156 36372 2212 36382
rect 2156 36278 2212 36316
rect 2268 35588 2324 36652
rect 2268 35494 2324 35532
rect 2156 35476 2212 35486
rect 2156 34244 2212 35420
rect 2268 35252 2324 35262
rect 2268 34468 2324 35196
rect 2268 34402 2324 34412
rect 2156 34188 2324 34244
rect 2156 34020 2212 34030
rect 2044 34018 2212 34020
rect 2044 33966 2158 34018
rect 2210 33966 2212 34018
rect 2044 33964 2212 33966
rect 2156 33954 2212 33964
rect 1932 33842 1988 33852
rect 2268 33796 2324 34188
rect 2156 33740 2324 33796
rect 1820 32722 1876 32732
rect 2044 33684 2100 33694
rect 1708 32452 1764 32462
rect 1708 32358 1764 32396
rect 2044 31892 2100 33628
rect 2044 31798 2100 31836
rect 1708 31780 1764 31790
rect 1708 31686 1764 31724
rect 1596 31054 1598 31106
rect 1650 31054 1652 31106
rect 1596 31042 1652 31054
rect 1484 30604 1652 30660
rect 1260 30258 1316 30268
rect 1036 30034 1092 30044
rect 1484 30098 1540 30110
rect 1484 30046 1486 30098
rect 1538 30046 1540 30098
rect 1036 29204 1092 29214
rect 1036 29110 1092 29148
rect 1036 28980 1092 28990
rect 1036 27970 1092 28924
rect 1484 28532 1540 30046
rect 1596 29538 1652 30604
rect 1596 29486 1598 29538
rect 1650 29486 1652 29538
rect 1596 29474 1652 29486
rect 1932 30100 1988 30110
rect 1540 28476 1652 28532
rect 1484 28466 1540 28476
rect 1036 27918 1038 27970
rect 1090 27918 1092 27970
rect 1036 27906 1092 27918
rect 1484 27860 1540 27870
rect 1148 27858 1540 27860
rect 1148 27806 1486 27858
rect 1538 27806 1540 27858
rect 1148 27804 1540 27806
rect 1148 27300 1204 27804
rect 1484 27794 1540 27804
rect 924 27244 1204 27300
rect 700 26852 868 26908
rect 588 13122 644 13132
rect 700 23940 756 23950
rect 700 5572 756 23884
rect 812 18676 868 26852
rect 812 18610 868 18620
rect 812 18452 868 18462
rect 812 9268 868 18396
rect 812 9202 868 9212
rect 700 5506 756 5516
rect 364 2818 420 2828
rect 924 1652 980 27244
rect 1036 27076 1092 27086
rect 1036 24162 1092 27020
rect 1260 27076 1316 27086
rect 1260 26982 1316 27020
rect 1596 26908 1652 28476
rect 1484 26852 1652 26908
rect 1708 27300 1764 27310
rect 1260 26516 1316 26526
rect 1260 25394 1316 26460
rect 1260 25342 1262 25394
rect 1314 25342 1316 25394
rect 1260 25330 1316 25342
rect 1036 24110 1038 24162
rect 1090 24110 1092 24162
rect 1036 24098 1092 24110
rect 1372 24948 1428 24958
rect 1036 23828 1092 23838
rect 1036 20188 1092 23772
rect 1148 23042 1204 23054
rect 1148 22990 1150 23042
rect 1202 22990 1204 23042
rect 1148 22372 1204 22990
rect 1148 22306 1204 22316
rect 1260 22260 1316 22270
rect 1260 22166 1316 22204
rect 1372 20690 1428 24892
rect 1484 23268 1540 26852
rect 1596 24164 1652 24174
rect 1596 24050 1652 24108
rect 1596 23998 1598 24050
rect 1650 23998 1652 24050
rect 1596 23986 1652 23998
rect 1484 22260 1540 23212
rect 1596 23604 1652 23614
rect 1596 23154 1652 23548
rect 1596 23102 1598 23154
rect 1650 23102 1652 23154
rect 1596 23090 1652 23102
rect 1708 23044 1764 27244
rect 1820 27076 1876 27086
rect 1820 25508 1876 27020
rect 1820 24722 1876 25452
rect 1820 24670 1822 24722
rect 1874 24670 1876 24722
rect 1820 24658 1876 24670
rect 1932 26292 1988 30044
rect 2044 28532 2100 28542
rect 2044 28438 2100 28476
rect 2156 28084 2212 33740
rect 2268 33572 2324 33582
rect 2268 33458 2324 33516
rect 2268 33406 2270 33458
rect 2322 33406 2324 33458
rect 2268 33394 2324 33406
rect 2268 30212 2324 30222
rect 2268 30118 2324 30156
rect 2380 28756 2436 41244
rect 2492 41076 2548 41086
rect 2492 41074 2660 41076
rect 2492 41022 2494 41074
rect 2546 41022 2660 41074
rect 2492 41020 2660 41022
rect 2492 41010 2548 41020
rect 2492 40516 2548 40526
rect 2492 40422 2548 40460
rect 2492 39844 2548 39854
rect 2492 39750 2548 39788
rect 2492 38052 2548 38062
rect 2492 35140 2548 37996
rect 2604 36708 2660 41020
rect 2828 40178 2884 40190
rect 2828 40126 2830 40178
rect 2882 40126 2884 40178
rect 2716 38610 2772 38622
rect 2716 38558 2718 38610
rect 2770 38558 2772 38610
rect 2716 38500 2772 38558
rect 2716 38434 2772 38444
rect 2828 38164 2884 40126
rect 2940 38668 2996 46508
rect 3052 41972 3108 41982
rect 3052 39730 3108 41916
rect 3052 39678 3054 39730
rect 3106 39678 3108 39730
rect 3052 39666 3108 39678
rect 3276 40514 3332 40526
rect 3276 40462 3278 40514
rect 3330 40462 3332 40514
rect 2940 38612 3108 38668
rect 2828 38098 2884 38108
rect 2828 37940 2884 37950
rect 2716 37380 2772 37390
rect 2716 37286 2772 37324
rect 2604 36642 2660 36652
rect 2604 36482 2660 36494
rect 2604 36430 2606 36482
rect 2658 36430 2660 36482
rect 2604 35364 2660 36430
rect 2716 35812 2772 35822
rect 2716 35718 2772 35756
rect 2604 35298 2660 35308
rect 2828 35252 2884 37884
rect 2828 35186 2884 35196
rect 2940 37826 2996 37838
rect 2940 37774 2942 37826
rect 2994 37774 2996 37826
rect 2492 35084 2660 35140
rect 2492 34802 2548 34814
rect 2492 34750 2494 34802
rect 2546 34750 2548 34802
rect 2492 34244 2548 34750
rect 2492 34178 2548 34188
rect 2492 34020 2548 34030
rect 2492 32564 2548 33964
rect 2604 33460 2660 35084
rect 2828 34804 2884 34814
rect 2716 34802 2884 34804
rect 2716 34750 2830 34802
rect 2882 34750 2884 34802
rect 2716 34748 2884 34750
rect 2716 33572 2772 34748
rect 2828 34738 2884 34748
rect 2828 34132 2884 34142
rect 2940 34132 2996 37774
rect 3052 36596 3108 38612
rect 3052 36530 3108 36540
rect 3164 37042 3220 37054
rect 3164 36990 3166 37042
rect 3218 36990 3220 37042
rect 3164 36484 3220 36990
rect 3052 36258 3108 36270
rect 3052 36206 3054 36258
rect 3106 36206 3108 36258
rect 3052 34916 3108 36206
rect 3164 35700 3220 36428
rect 3164 35634 3220 35644
rect 3164 34916 3220 34926
rect 3052 34914 3220 34916
rect 3052 34862 3166 34914
rect 3218 34862 3220 34914
rect 3052 34860 3220 34862
rect 3164 34850 3220 34860
rect 2828 34130 2996 34132
rect 2828 34078 2830 34130
rect 2882 34078 2996 34130
rect 2828 34076 2996 34078
rect 2828 34066 2884 34076
rect 2716 33506 2772 33516
rect 2940 33684 2996 33694
rect 3276 33684 3332 40462
rect 3500 39732 3556 55246
rect 6076 55188 6132 57344
rect 7420 56194 7476 57344
rect 8764 56644 8820 57344
rect 10108 56756 10164 57344
rect 10108 56700 10612 56756
rect 8764 56588 9044 56644
rect 8988 56306 9044 56588
rect 8988 56254 8990 56306
rect 9042 56254 9044 56306
rect 8988 56242 9044 56254
rect 10556 56306 10612 56700
rect 10556 56254 10558 56306
rect 10610 56254 10612 56306
rect 10556 56242 10612 56254
rect 7420 56142 7422 56194
rect 7474 56142 7476 56194
rect 7420 56130 7476 56142
rect 6188 55970 6244 55982
rect 6188 55918 6190 55970
rect 6242 55918 6244 55970
rect 6188 55860 6244 55918
rect 6188 55794 6244 55804
rect 8092 55970 8148 55982
rect 8092 55918 8094 55970
rect 8146 55918 8148 55970
rect 6076 55122 6132 55132
rect 6300 55298 6356 55310
rect 6300 55246 6302 55298
rect 6354 55246 6356 55298
rect 3804 54908 4068 54918
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 3804 54842 4068 54852
rect 4464 54124 4728 54134
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4464 54058 4728 54068
rect 3804 53340 4068 53350
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 3804 53274 4068 53284
rect 4464 52556 4728 52566
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4464 52490 4728 52500
rect 3804 51772 4068 51782
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 3804 51706 4068 51716
rect 5852 51268 5908 51278
rect 4464 50988 4728 50998
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4464 50922 4728 50932
rect 3804 50204 4068 50214
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 3804 50138 4068 50148
rect 4464 49420 4728 49430
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4464 49354 4728 49364
rect 3804 48636 4068 48646
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 3804 48570 4068 48580
rect 5628 48468 5684 48478
rect 4464 47852 4728 47862
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4464 47786 4728 47796
rect 3804 47068 4068 47078
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 3804 47002 4068 47012
rect 4464 46284 4728 46294
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4464 46218 4728 46228
rect 3804 45500 4068 45510
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 3804 45434 4068 45444
rect 4464 44716 4728 44726
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4464 44650 4728 44660
rect 3804 43932 4068 43942
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 3804 43866 4068 43876
rect 5628 43708 5684 48412
rect 5628 43652 5796 43708
rect 4464 43148 4728 43158
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4464 43082 4728 43092
rect 3804 42364 4068 42374
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 3804 42298 4068 42308
rect 5516 42084 5572 42094
rect 4464 41580 4728 41590
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4464 41514 4728 41524
rect 3804 40796 4068 40806
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 3804 40730 4068 40740
rect 4464 40012 4728 40022
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4464 39946 4728 39956
rect 3500 39666 3556 39676
rect 3948 39620 4004 39630
rect 3948 39526 4004 39564
rect 3500 39506 3556 39518
rect 3500 39454 3502 39506
rect 3554 39454 3556 39506
rect 3500 39396 3556 39454
rect 3500 39330 3556 39340
rect 5180 39396 5236 39406
rect 3804 39228 4068 39238
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 3804 39162 4068 39172
rect 3836 38610 3892 38622
rect 3836 38558 3838 38610
rect 3890 38558 3892 38610
rect 3836 37828 3892 38558
rect 3500 37772 3892 37828
rect 4172 38500 4228 38510
rect 3388 34132 3444 34142
rect 3388 34038 3444 34076
rect 2604 33394 2660 33404
rect 2716 33346 2772 33358
rect 2716 33294 2718 33346
rect 2770 33294 2772 33346
rect 2716 32788 2772 33294
rect 2828 32788 2884 32798
rect 2716 32786 2884 32788
rect 2716 32734 2830 32786
rect 2882 32734 2884 32786
rect 2716 32732 2884 32734
rect 2828 32722 2884 32732
rect 2492 32508 2884 32564
rect 2380 28662 2436 28700
rect 2492 31892 2548 31902
rect 2156 28028 2436 28084
rect 2268 27858 2324 27870
rect 2268 27806 2270 27858
rect 2322 27806 2324 27858
rect 2268 27076 2324 27806
rect 1708 22978 1764 22988
rect 1932 23828 1988 26236
rect 1596 22484 1652 22494
rect 1596 22390 1652 22428
rect 1484 22194 1540 22204
rect 1708 22260 1764 22270
rect 1596 22148 1652 22158
rect 1372 20638 1374 20690
rect 1426 20638 1428 20690
rect 1372 20626 1428 20638
rect 1484 22036 1540 22046
rect 1036 20132 1316 20188
rect 1148 19348 1204 19358
rect 1036 17556 1092 17566
rect 1036 8036 1092 17500
rect 1148 16660 1204 19292
rect 1260 19122 1316 20132
rect 1260 19070 1262 19122
rect 1314 19070 1316 19122
rect 1260 19058 1316 19070
rect 1260 17108 1316 17118
rect 1260 16994 1316 17052
rect 1260 16942 1262 16994
rect 1314 16942 1316 16994
rect 1260 16930 1316 16942
rect 1148 16604 1316 16660
rect 1148 12180 1204 12190
rect 1148 8260 1204 12124
rect 1260 9714 1316 16604
rect 1372 16324 1428 16334
rect 1372 16098 1428 16268
rect 1372 16046 1374 16098
rect 1426 16046 1428 16098
rect 1372 15316 1428 16046
rect 1372 15250 1428 15260
rect 1260 9662 1262 9714
rect 1314 9662 1316 9714
rect 1260 9650 1316 9662
rect 1372 13972 1428 13982
rect 1260 9268 1316 9278
rect 1260 9174 1316 9212
rect 1372 8428 1428 13916
rect 1484 13074 1540 21980
rect 1596 19012 1652 22092
rect 1596 18946 1652 18956
rect 1708 20018 1764 22204
rect 1820 20916 1876 20926
rect 1820 20822 1876 20860
rect 1708 19966 1710 20018
rect 1762 19966 1764 20018
rect 1596 18788 1652 18798
rect 1596 18450 1652 18732
rect 1596 18398 1598 18450
rect 1650 18398 1652 18450
rect 1596 18386 1652 18398
rect 1708 17108 1764 19966
rect 1820 17671 1876 17683
rect 1820 17619 1822 17671
rect 1874 17619 1876 17671
rect 1820 17444 1876 17619
rect 1820 17378 1876 17388
rect 1708 17042 1764 17052
rect 1820 16884 1876 16894
rect 1596 16772 1652 16782
rect 1596 15204 1652 16716
rect 1820 16436 1876 16828
rect 1708 16380 1876 16436
rect 1708 15314 1764 16380
rect 1820 16212 1876 16222
rect 1820 16118 1876 16156
rect 1708 15262 1710 15314
rect 1762 15262 1764 15314
rect 1708 15250 1764 15262
rect 1820 15316 1876 15326
rect 1596 15138 1652 15148
rect 1708 14532 1764 14542
rect 1820 14532 1876 15260
rect 1708 14530 1876 14532
rect 1708 14478 1710 14530
rect 1762 14478 1876 14530
rect 1708 14476 1876 14478
rect 1708 14466 1764 14476
rect 1932 14308 1988 23772
rect 2044 27020 2324 27076
rect 2044 26402 2100 27020
rect 2380 26964 2436 28028
rect 2268 26908 2436 26964
rect 2044 26350 2046 26402
rect 2098 26350 2100 26402
rect 2044 23044 2100 26350
rect 2156 26852 2324 26908
rect 2156 25506 2212 26852
rect 2492 26178 2548 31836
rect 2716 31892 2772 31902
rect 2716 31106 2772 31836
rect 2716 31054 2718 31106
rect 2770 31054 2772 31106
rect 2716 31042 2772 31054
rect 2716 30324 2772 30334
rect 2604 30212 2660 30222
rect 2604 29428 2660 30156
rect 2604 28980 2660 29372
rect 2604 28914 2660 28924
rect 2492 26126 2494 26178
rect 2546 26126 2548 26178
rect 2156 25454 2158 25506
rect 2210 25454 2212 25506
rect 2156 25442 2212 25454
rect 2268 25844 2324 25854
rect 2268 23604 2324 25788
rect 2380 24612 2436 24650
rect 2380 24546 2436 24556
rect 2380 24388 2436 24398
rect 2380 23940 2436 24332
rect 2380 23846 2436 23884
rect 2268 23548 2436 23604
rect 2268 23268 2324 23306
rect 2268 23202 2324 23212
rect 2268 23044 2324 23054
rect 2044 22988 2212 23044
rect 2044 22820 2100 22830
rect 2044 16772 2100 22764
rect 2156 21700 2212 22988
rect 2156 21634 2212 21644
rect 2156 20692 2212 20702
rect 2156 20598 2212 20636
rect 2156 19794 2212 19806
rect 2156 19742 2158 19794
rect 2210 19742 2212 19794
rect 2156 19124 2212 19742
rect 2268 19572 2324 22988
rect 2268 19506 2324 19516
rect 2268 19348 2324 19358
rect 2380 19348 2436 23548
rect 2268 19346 2436 19348
rect 2268 19294 2270 19346
rect 2322 19294 2436 19346
rect 2268 19292 2436 19294
rect 2268 19282 2324 19292
rect 2492 19124 2548 26126
rect 2716 27746 2772 30268
rect 2716 27694 2718 27746
rect 2770 27694 2772 27746
rect 2604 25394 2660 25406
rect 2604 25342 2606 25394
rect 2658 25342 2660 25394
rect 2604 24836 2660 25342
rect 2604 24770 2660 24780
rect 2716 24612 2772 27694
rect 2828 27188 2884 32508
rect 2940 30100 2996 33628
rect 3164 33628 3332 33684
rect 3052 33346 3108 33358
rect 3052 33294 3054 33346
rect 3106 33294 3108 33346
rect 3052 30548 3108 33294
rect 3164 30996 3220 33628
rect 3276 33460 3332 33470
rect 3276 33458 3444 33460
rect 3276 33406 3278 33458
rect 3330 33406 3444 33458
rect 3276 33404 3444 33406
rect 3276 33394 3332 33404
rect 3388 32562 3444 33404
rect 3388 32510 3390 32562
rect 3442 32510 3444 32562
rect 3388 32498 3444 32510
rect 3500 32340 3556 37772
rect 3804 37660 4068 37670
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 3804 37594 4068 37604
rect 4172 37156 4228 38444
rect 4464 38444 4728 38454
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4464 38378 4728 38388
rect 4732 38162 4788 38174
rect 4732 38110 4734 38162
rect 4786 38110 4788 38162
rect 4396 37938 4452 37950
rect 4396 37886 4398 37938
rect 4450 37886 4452 37938
rect 4396 37828 4452 37886
rect 4732 37940 4788 38110
rect 4732 37874 4788 37884
rect 4396 37762 4452 37772
rect 5068 37828 5124 37838
rect 4172 36706 4228 37100
rect 4844 37380 4900 37390
rect 4172 36654 4174 36706
rect 4226 36654 4228 36706
rect 3804 36092 4068 36102
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 3804 36026 4068 36036
rect 3948 35700 4004 35710
rect 4172 35700 4228 36654
rect 3948 35698 4228 35700
rect 3948 35646 3950 35698
rect 4002 35646 4228 35698
rect 3948 35644 4228 35646
rect 4284 37042 4340 37054
rect 4284 36990 4286 37042
rect 4338 36990 4340 37042
rect 3724 35364 3780 35374
rect 3612 35140 3668 35150
rect 3724 35140 3780 35308
rect 3836 35140 3892 35150
rect 3724 35138 3892 35140
rect 3724 35086 3838 35138
rect 3890 35086 3892 35138
rect 3724 35084 3892 35086
rect 3612 34914 3668 35084
rect 3836 35074 3892 35084
rect 3948 35028 4004 35644
rect 3948 34962 4004 34972
rect 4284 35026 4340 36990
rect 4464 36876 4728 36886
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4464 36810 4728 36820
rect 4732 36484 4788 36494
rect 4844 36484 4900 37324
rect 4732 36482 5012 36484
rect 4732 36430 4734 36482
rect 4786 36430 5012 36482
rect 4732 36428 5012 36430
rect 4732 36418 4788 36428
rect 4396 35700 4452 35710
rect 4396 35606 4452 35644
rect 4844 35588 4900 35598
rect 4464 35308 4728 35318
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4464 35242 4728 35252
rect 4844 35140 4900 35532
rect 4284 34974 4286 35026
rect 4338 34974 4340 35026
rect 4284 34962 4340 34974
rect 4508 35084 4900 35140
rect 3612 34862 3614 34914
rect 3666 34862 3668 34914
rect 3612 33908 3668 34862
rect 3804 34524 4068 34534
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 3804 34458 4068 34468
rect 4284 34468 4340 34478
rect 3612 33842 3668 33852
rect 4172 34356 4228 34366
rect 3724 33348 3780 33358
rect 3388 32284 3556 32340
rect 3612 33346 3780 33348
rect 3612 33294 3726 33346
rect 3778 33294 3780 33346
rect 3612 33292 3780 33294
rect 3276 31780 3332 31790
rect 3276 31686 3332 31724
rect 3164 30940 3332 30996
rect 3164 30772 3220 30782
rect 3164 30678 3220 30716
rect 3052 30492 3220 30548
rect 3052 30100 3108 30110
rect 2940 30098 3108 30100
rect 2940 30046 3054 30098
rect 3106 30046 3108 30098
rect 2940 30044 3108 30046
rect 3052 30034 3108 30044
rect 3164 30100 3220 30492
rect 3164 30034 3220 30044
rect 2828 27122 2884 27132
rect 3052 29876 3108 29886
rect 3052 26908 3108 29820
rect 3164 29316 3220 29326
rect 3276 29316 3332 30940
rect 3388 29988 3444 32284
rect 3612 31780 3668 33292
rect 3724 33282 3780 33292
rect 3804 32956 4068 32966
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 3804 32890 4068 32900
rect 3836 32676 3892 32686
rect 4172 32676 4228 34300
rect 4284 34130 4340 34412
rect 4284 34078 4286 34130
rect 4338 34078 4340 34130
rect 4284 34066 4340 34078
rect 4508 33908 4564 35084
rect 3836 32674 4228 32676
rect 3836 32622 3838 32674
rect 3890 32622 4228 32674
rect 3836 32620 4228 32622
rect 4284 33852 4564 33908
rect 4844 34914 4900 34926
rect 4844 34862 4846 34914
rect 4898 34862 4900 34914
rect 4844 34132 4900 34862
rect 3836 32610 3892 32620
rect 3612 31714 3668 31724
rect 4284 31444 4340 33852
rect 4464 33740 4728 33750
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4464 33674 4728 33684
rect 4508 33346 4564 33358
rect 4508 33294 4510 33346
rect 4562 33294 4564 33346
rect 4508 32900 4564 33294
rect 4844 32900 4900 34076
rect 4508 32844 4900 32900
rect 4464 32172 4728 32182
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4464 32106 4728 32116
rect 3804 31388 4068 31398
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 3804 31322 4068 31332
rect 4172 31388 4340 31444
rect 4172 30324 4228 31388
rect 4284 31220 4340 31230
rect 4284 31126 4340 31164
rect 4464 30604 4728 30614
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4464 30538 4728 30548
rect 3836 30212 3892 30222
rect 3612 30210 3892 30212
rect 3612 30158 3838 30210
rect 3890 30158 3892 30210
rect 3612 30156 3892 30158
rect 3388 29922 3444 29932
rect 3500 30098 3556 30110
rect 3500 30046 3502 30098
rect 3554 30046 3556 30098
rect 3164 29314 3332 29316
rect 3164 29262 3166 29314
rect 3218 29262 3332 29314
rect 3164 29260 3332 29262
rect 3164 27300 3220 29260
rect 3500 28868 3556 30046
rect 3500 28802 3556 28812
rect 3612 28866 3668 30156
rect 3836 30146 3892 30156
rect 3804 29820 4068 29830
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 3804 29754 4068 29764
rect 4172 29652 4228 30268
rect 4396 30436 4452 30446
rect 4284 30210 4340 30222
rect 4284 30158 4286 30210
rect 4338 30158 4340 30210
rect 4284 30100 4340 30158
rect 4284 30034 4340 30044
rect 3612 28814 3614 28866
rect 3666 28814 3668 28866
rect 3612 28802 3668 28814
rect 3724 29596 4228 29652
rect 4284 29652 4340 29662
rect 3724 28644 3780 29596
rect 4284 29558 4340 29596
rect 3164 27234 3220 27244
rect 3500 28588 3780 28644
rect 4172 29428 4228 29438
rect 4396 29428 4452 30380
rect 4508 30322 4564 30334
rect 4508 30270 4510 30322
rect 4562 30270 4564 30322
rect 4508 30212 4564 30270
rect 4508 30146 4564 30156
rect 4172 28642 4228 29372
rect 4172 28590 4174 28642
rect 4226 28590 4228 28642
rect 3276 27188 3332 27198
rect 3332 27132 3444 27188
rect 3276 27122 3332 27132
rect 3276 26964 3332 27002
rect 2828 26850 2884 26862
rect 3052 26852 3220 26908
rect 3276 26898 3332 26908
rect 2828 26798 2830 26850
rect 2882 26798 2884 26850
rect 2828 25508 2884 26798
rect 3052 26516 3108 26526
rect 3052 25844 3108 26460
rect 3052 25778 3108 25788
rect 2940 25508 2996 25518
rect 2828 25506 2996 25508
rect 2828 25454 2942 25506
rect 2994 25454 2996 25506
rect 2828 25452 2996 25454
rect 2940 25442 2996 25452
rect 2604 24556 2772 24612
rect 2604 22820 2660 24556
rect 3164 24164 3220 26852
rect 3388 26740 3444 27132
rect 3052 24108 3220 24164
rect 3276 26684 3444 26740
rect 2828 23938 2884 23950
rect 2828 23886 2830 23938
rect 2882 23886 2884 23938
rect 2716 23156 2772 23166
rect 2716 23042 2772 23100
rect 2716 22990 2718 23042
rect 2770 22990 2772 23042
rect 2716 22978 2772 22990
rect 2604 22754 2660 22764
rect 2828 22594 2884 23886
rect 2828 22542 2830 22594
rect 2882 22542 2884 22594
rect 2828 22530 2884 22542
rect 2940 23044 2996 23054
rect 2716 21700 2772 21710
rect 2156 19068 2548 19124
rect 2380 18900 2436 18910
rect 2156 18676 2212 18686
rect 2156 18450 2212 18620
rect 2156 18398 2158 18450
rect 2210 18398 2212 18450
rect 2156 18386 2212 18398
rect 2268 18564 2324 18574
rect 2044 16706 2100 16716
rect 2156 15428 2212 15438
rect 2268 15428 2324 18508
rect 2380 16212 2436 18844
rect 2380 16146 2436 16156
rect 2156 15426 2324 15428
rect 2156 15374 2158 15426
rect 2210 15374 2324 15426
rect 2156 15372 2324 15374
rect 2156 15362 2212 15372
rect 2268 15204 2324 15214
rect 2156 15092 2212 15102
rect 2156 14754 2212 15036
rect 2156 14702 2158 14754
rect 2210 14702 2212 14754
rect 2156 14690 2212 14702
rect 1932 14252 2212 14308
rect 1484 13022 1486 13074
rect 1538 13022 1540 13074
rect 1484 13010 1540 13022
rect 1708 13748 1764 13758
rect 1708 12516 1764 13692
rect 1820 13746 1876 13758
rect 1820 13694 1822 13746
rect 1874 13694 1876 13746
rect 1820 13300 1876 13694
rect 1820 13234 1876 13244
rect 2044 12962 2100 12974
rect 2044 12910 2046 12962
rect 2098 12910 2100 12962
rect 2044 12516 2100 12910
rect 1596 12460 1764 12516
rect 1932 12460 2100 12516
rect 1596 12180 1652 12460
rect 1596 12124 1876 12180
rect 1596 11620 1652 11630
rect 1596 11526 1652 11564
rect 1820 8428 1876 12124
rect 1932 11620 1988 12460
rect 2044 12180 2100 12190
rect 2044 12086 2100 12124
rect 1932 11554 1988 11564
rect 1932 10724 1988 10734
rect 1932 9380 1988 10668
rect 2044 10610 2100 10622
rect 2044 10558 2046 10610
rect 2098 10558 2100 10610
rect 2044 10500 2100 10558
rect 2044 10434 2100 10444
rect 1932 9324 2100 9380
rect 1372 8372 1540 8428
rect 1820 8372 1988 8428
rect 1148 8204 1428 8260
rect 1260 8036 1316 8046
rect 1036 8034 1316 8036
rect 1036 7982 1262 8034
rect 1314 7982 1316 8034
rect 1036 7980 1316 7982
rect 1260 7970 1316 7980
rect 1372 6578 1428 8204
rect 1484 7586 1540 8372
rect 1484 7534 1486 7586
rect 1538 7534 1540 7586
rect 1484 7522 1540 7534
rect 1596 8260 1652 8270
rect 1372 6526 1374 6578
rect 1426 6526 1428 6578
rect 1372 6514 1428 6526
rect 1484 6804 1540 6814
rect 1484 5234 1540 6748
rect 1596 6018 1652 8204
rect 1596 5966 1598 6018
rect 1650 5966 1652 6018
rect 1596 5954 1652 5966
rect 1484 5182 1486 5234
rect 1538 5182 1540 5234
rect 1484 5170 1540 5182
rect 1596 5572 1652 5582
rect 1036 5012 1092 5022
rect 1036 2770 1092 4956
rect 1484 4226 1540 4238
rect 1484 4174 1486 4226
rect 1538 4174 1540 4226
rect 1484 4116 1540 4174
rect 1484 4050 1540 4060
rect 1260 3330 1316 3342
rect 1260 3278 1262 3330
rect 1314 3278 1316 3330
rect 1260 3220 1316 3278
rect 1260 3154 1316 3164
rect 1484 2884 1540 2894
rect 1484 2790 1540 2828
rect 1036 2718 1038 2770
rect 1090 2718 1092 2770
rect 1036 2706 1092 2718
rect 1036 2324 1092 2334
rect 1036 2210 1092 2268
rect 1036 2158 1038 2210
rect 1090 2158 1092 2210
rect 1036 2146 1092 2158
rect 1596 2098 1652 5516
rect 1932 5124 1988 8372
rect 2044 6690 2100 9324
rect 2156 8708 2212 14252
rect 2268 13524 2324 15148
rect 2268 13430 2324 13468
rect 2268 13300 2324 13310
rect 2268 12180 2324 13244
rect 2268 12114 2324 12124
rect 2380 12964 2436 12974
rect 2380 11956 2436 12908
rect 2492 12964 2548 19068
rect 2604 20802 2660 20814
rect 2604 20750 2606 20802
rect 2658 20750 2660 20802
rect 2604 18340 2660 20750
rect 2716 18562 2772 21644
rect 2940 21588 2996 22988
rect 2716 18510 2718 18562
rect 2770 18510 2772 18562
rect 2716 18498 2772 18510
rect 2828 21532 2996 21588
rect 3052 22484 3108 24108
rect 3164 23938 3220 23950
rect 3164 23886 3166 23938
rect 3218 23886 3220 23938
rect 3164 23828 3220 23886
rect 3164 23762 3220 23772
rect 3276 23156 3332 26684
rect 3388 25506 3444 25518
rect 3388 25454 3390 25506
rect 3442 25454 3444 25506
rect 3388 25396 3444 25454
rect 3388 25330 3444 25340
rect 3500 25172 3556 28588
rect 4172 28578 4228 28590
rect 4284 29372 4452 29428
rect 3804 28252 4068 28262
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 3804 28186 4068 28196
rect 4284 27860 4340 29372
rect 4464 29036 4728 29046
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4464 28970 4728 28980
rect 3836 27804 4340 27860
rect 3612 27074 3668 27086
rect 3612 27022 3614 27074
rect 3666 27022 3668 27074
rect 3612 26514 3668 27022
rect 3836 26908 3892 27804
rect 3948 27636 4004 27646
rect 3948 27634 4228 27636
rect 3948 27582 3950 27634
rect 4002 27582 4228 27634
rect 3948 27580 4228 27582
rect 3948 27570 4004 27580
rect 4060 27188 4116 27198
rect 4060 27074 4116 27132
rect 4060 27022 4062 27074
rect 4114 27022 4116 27074
rect 4060 27010 4116 27022
rect 4172 27076 4228 27580
rect 4464 27468 4728 27478
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4464 27402 4728 27412
rect 4284 27300 4340 27310
rect 4284 27206 4340 27244
rect 4732 27076 4788 27086
rect 4172 27074 4788 27076
rect 4172 27022 4734 27074
rect 4786 27022 4788 27074
rect 4172 27020 4788 27022
rect 4732 27010 4788 27020
rect 3836 26852 4340 26908
rect 3804 26684 4068 26694
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 3804 26618 4068 26628
rect 3612 26462 3614 26514
rect 3666 26462 3668 26514
rect 3612 26450 3668 26462
rect 3612 25732 3668 25742
rect 3612 25638 3668 25676
rect 4060 25506 4116 25518
rect 4060 25454 4062 25506
rect 4114 25454 4116 25506
rect 4060 25284 4116 25454
rect 3388 25116 3556 25172
rect 3612 25228 4116 25284
rect 3388 24276 3444 25116
rect 3500 24948 3556 24958
rect 3612 24948 3668 25228
rect 4172 25172 4228 25182
rect 3804 25116 4068 25126
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 3804 25050 4068 25060
rect 3500 24946 3668 24948
rect 3500 24894 3502 24946
rect 3554 24894 3668 24946
rect 3500 24892 3668 24894
rect 3500 24882 3556 24892
rect 3724 24724 3780 24734
rect 3388 24220 3668 24276
rect 3388 24050 3444 24062
rect 3388 23998 3390 24050
rect 3442 23998 3444 24050
rect 3388 23604 3444 23998
rect 3388 23538 3444 23548
rect 3500 24052 3556 24062
rect 3276 23090 3332 23100
rect 2828 18564 2884 21532
rect 3052 21476 3108 22428
rect 3500 22258 3556 23996
rect 3500 22206 3502 22258
rect 3554 22206 3556 22258
rect 3500 22194 3556 22206
rect 2828 18498 2884 18508
rect 2940 21474 3108 21476
rect 2940 21422 3054 21474
rect 3106 21422 3108 21474
rect 2940 21420 3108 21422
rect 2604 18284 2884 18340
rect 2716 17780 2772 17790
rect 2716 17666 2772 17724
rect 2716 17614 2718 17666
rect 2770 17614 2772 17666
rect 2716 17602 2772 17614
rect 2828 17106 2884 18284
rect 2940 17892 2996 21420
rect 3052 21410 3108 21420
rect 3052 21028 3108 21038
rect 3612 21028 3668 24220
rect 3724 24052 3780 24668
rect 4172 24388 4228 25116
rect 4172 24322 4228 24332
rect 3724 23986 3780 23996
rect 4060 23940 4116 23950
rect 4060 23938 4228 23940
rect 4060 23886 4062 23938
rect 4114 23886 4228 23938
rect 4060 23884 4228 23886
rect 4060 23874 4116 23884
rect 3804 23548 4068 23558
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 3804 23482 4068 23492
rect 3836 23380 3892 23390
rect 4172 23380 4228 23884
rect 3836 23378 4228 23380
rect 3836 23326 3838 23378
rect 3890 23326 4228 23378
rect 3836 23324 4228 23326
rect 3836 23314 3892 23324
rect 4284 22370 4340 26852
rect 4464 25900 4728 25910
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4464 25834 4728 25844
rect 4844 25732 4900 32844
rect 4956 32788 5012 36428
rect 4956 32722 5012 32732
rect 5068 33908 5124 37772
rect 5068 32562 5124 33852
rect 5068 32510 5070 32562
rect 5122 32510 5124 32562
rect 5068 32498 5124 32510
rect 5180 34130 5236 39340
rect 5404 39284 5460 39294
rect 5404 38946 5460 39228
rect 5404 38894 5406 38946
rect 5458 38894 5460 38946
rect 5404 37828 5460 38894
rect 5404 37762 5460 37772
rect 5292 36258 5348 36270
rect 5292 36206 5294 36258
rect 5346 36206 5348 36258
rect 5292 35476 5348 36206
rect 5292 35410 5348 35420
rect 5404 36148 5460 36158
rect 5180 34078 5182 34130
rect 5234 34078 5236 34130
rect 4956 32450 5012 32462
rect 4956 32398 4958 32450
rect 5010 32398 5012 32450
rect 4956 31892 5012 32398
rect 4956 30660 5012 31836
rect 5068 31668 5124 31678
rect 5068 31574 5124 31612
rect 4956 30594 5012 30604
rect 5068 30994 5124 31006
rect 5068 30942 5070 30994
rect 5122 30942 5124 30994
rect 4956 30210 5012 30222
rect 4956 30158 4958 30210
rect 5010 30158 5012 30210
rect 4956 29652 5012 30158
rect 5068 30212 5124 30942
rect 5068 30146 5124 30156
rect 4956 29586 5012 29596
rect 5068 29988 5124 29998
rect 4956 29428 5012 29438
rect 4956 28530 5012 29372
rect 4956 28478 4958 28530
rect 5010 28478 5012 28530
rect 4956 27860 5012 28478
rect 4956 27794 5012 27804
rect 4956 27634 5012 27646
rect 4956 27582 4958 27634
rect 5010 27582 5012 27634
rect 4956 27300 5012 27582
rect 4956 27234 5012 27244
rect 4732 25676 4900 25732
rect 4956 26066 5012 26078
rect 4956 26014 4958 26066
rect 5010 26014 5012 26066
rect 4956 25732 5012 26014
rect 4620 25506 4676 25518
rect 4620 25454 4622 25506
rect 4674 25454 4676 25506
rect 4620 24612 4676 25454
rect 4732 25508 4788 25676
rect 4956 25666 5012 25676
rect 4732 25452 5012 25508
rect 4620 24546 4676 24556
rect 4464 24332 4728 24342
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4464 24266 4728 24276
rect 4620 23938 4676 23950
rect 4620 23886 4622 23938
rect 4674 23886 4676 23938
rect 4620 23604 4676 23886
rect 4620 23538 4676 23548
rect 4464 22764 4728 22774
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4464 22698 4728 22708
rect 4284 22318 4286 22370
rect 4338 22318 4340 22370
rect 4284 22306 4340 22318
rect 3804 21980 4068 21990
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 3804 21914 4068 21924
rect 4956 21812 5012 25452
rect 5068 24722 5124 29932
rect 5180 28980 5236 34078
rect 5292 34916 5348 34926
rect 5292 34468 5348 34860
rect 5292 33346 5348 34412
rect 5292 33294 5294 33346
rect 5346 33294 5348 33346
rect 5292 30996 5348 33294
rect 5404 32116 5460 36092
rect 5516 35810 5572 42028
rect 5516 35758 5518 35810
rect 5570 35758 5572 35810
rect 5516 35746 5572 35758
rect 5628 34132 5684 34142
rect 5516 33908 5572 33918
rect 5516 33814 5572 33852
rect 5516 32340 5572 32350
rect 5516 32246 5572 32284
rect 5404 32060 5572 32116
rect 5404 31778 5460 31790
rect 5404 31726 5406 31778
rect 5458 31726 5460 31778
rect 5404 31220 5460 31726
rect 5404 31154 5460 31164
rect 5516 31106 5572 32060
rect 5516 31054 5518 31106
rect 5570 31054 5572 31106
rect 5516 31042 5572 31054
rect 5628 31668 5684 34076
rect 5292 30940 5460 30996
rect 5292 30660 5348 30670
rect 5292 29428 5348 30604
rect 5292 29362 5348 29372
rect 5180 28914 5236 28924
rect 5068 24670 5070 24722
rect 5122 24670 5124 24722
rect 5068 24658 5124 24670
rect 5180 28756 5236 28766
rect 5180 23156 5236 28700
rect 5292 27076 5348 27086
rect 5292 26982 5348 27020
rect 5404 26908 5460 30940
rect 5516 30884 5572 30894
rect 5516 30210 5572 30828
rect 5628 30660 5684 31612
rect 5740 30884 5796 43652
rect 5852 41412 5908 51212
rect 6300 43708 6356 55246
rect 6860 55188 6916 55198
rect 6860 55094 6916 55132
rect 7756 51268 7812 51278
rect 5852 41346 5908 41356
rect 5964 43652 6356 43708
rect 7644 45780 7700 45790
rect 5964 40292 6020 43652
rect 6748 42980 6804 42990
rect 5964 40226 6020 40236
rect 6076 40402 6132 40414
rect 6412 40404 6468 40414
rect 6076 40350 6078 40402
rect 6130 40350 6132 40402
rect 6076 40180 6132 40350
rect 6076 40114 6132 40124
rect 6188 40402 6468 40404
rect 6188 40350 6414 40402
rect 6466 40350 6468 40402
rect 6188 40348 6468 40350
rect 5852 39844 5908 39854
rect 5852 38722 5908 39788
rect 6188 39060 6244 40348
rect 6412 40338 6468 40348
rect 5852 38670 5854 38722
rect 5906 38670 5908 38722
rect 5852 38658 5908 38670
rect 5964 39004 6244 39060
rect 6300 40180 6356 40190
rect 5964 38274 6020 39004
rect 5964 38222 5966 38274
rect 6018 38222 6020 38274
rect 5964 38210 6020 38222
rect 6300 38724 6356 40124
rect 5964 35474 6020 35486
rect 5964 35422 5966 35474
rect 6018 35422 6020 35474
rect 5852 34916 5908 34926
rect 5852 34822 5908 34860
rect 5964 33908 6020 35422
rect 6300 34132 6356 38668
rect 6412 39508 6468 39518
rect 6412 36594 6468 39452
rect 6524 39506 6580 39518
rect 6524 39454 6526 39506
rect 6578 39454 6580 39506
rect 6524 37940 6580 39454
rect 6636 39396 6692 39406
rect 6636 38050 6692 39340
rect 6636 37998 6638 38050
rect 6690 37998 6692 38050
rect 6636 37986 6692 37998
rect 6524 37874 6580 37884
rect 6524 37380 6580 37390
rect 6524 37286 6580 37324
rect 6412 36542 6414 36594
rect 6466 36542 6468 36594
rect 6412 36484 6468 36542
rect 6412 36418 6468 36428
rect 6524 35812 6580 35822
rect 6524 34914 6580 35756
rect 6524 34862 6526 34914
rect 6578 34862 6580 34914
rect 6524 34850 6580 34862
rect 6300 34066 6356 34076
rect 6188 33908 6244 33918
rect 6636 33908 6692 33918
rect 5964 33852 6188 33908
rect 5964 31892 6020 31902
rect 5964 31778 6020 31836
rect 5964 31726 5966 31778
rect 6018 31726 6020 31778
rect 5964 31714 6020 31726
rect 6076 31890 6132 31902
rect 6076 31838 6078 31890
rect 6130 31838 6132 31890
rect 5964 30996 6020 31006
rect 6076 30996 6132 31838
rect 5964 30994 6132 30996
rect 5964 30942 5966 30994
rect 6018 30942 6132 30994
rect 5964 30940 6132 30942
rect 5964 30930 6020 30940
rect 5796 30828 5908 30884
rect 5740 30818 5796 30828
rect 5628 30604 5796 30660
rect 5516 30158 5518 30210
rect 5570 30158 5572 30210
rect 5516 27972 5572 30158
rect 5628 29428 5684 29438
rect 5628 29334 5684 29372
rect 5628 28642 5684 28654
rect 5628 28590 5630 28642
rect 5682 28590 5684 28642
rect 5628 28420 5684 28590
rect 5628 28354 5684 28364
rect 5740 28196 5796 30604
rect 5852 29316 5908 30828
rect 5964 29316 6020 29326
rect 5852 29314 6020 29316
rect 5852 29262 5966 29314
rect 6018 29262 6020 29314
rect 5852 29260 6020 29262
rect 5852 28756 5908 29260
rect 5964 29250 6020 29260
rect 5852 28690 5908 28700
rect 6076 28980 6132 28990
rect 5740 28130 5796 28140
rect 5964 28308 6020 28318
rect 5516 27916 5908 27972
rect 5516 27746 5572 27758
rect 5516 27694 5518 27746
rect 5570 27694 5572 27746
rect 5516 27412 5572 27694
rect 5516 27346 5572 27356
rect 5740 27748 5796 27758
rect 5404 26852 5684 26908
rect 5516 26740 5572 26750
rect 5516 26402 5572 26684
rect 5516 26350 5518 26402
rect 5570 26350 5572 26402
rect 5516 26338 5572 26350
rect 5516 25620 5572 25630
rect 5404 25060 5460 25070
rect 5292 24724 5348 24734
rect 5292 23266 5348 24668
rect 5404 23940 5460 25004
rect 5516 24946 5572 25564
rect 5516 24894 5518 24946
rect 5570 24894 5572 24946
rect 5516 24882 5572 24894
rect 5628 24164 5684 26852
rect 5740 25732 5796 27692
rect 5740 25666 5796 25676
rect 5740 25508 5796 25518
rect 5740 25414 5796 25452
rect 5852 25172 5908 27916
rect 5852 25106 5908 25116
rect 5964 27188 6020 28252
rect 5628 24108 5796 24164
rect 5516 23940 5572 23950
rect 5404 23884 5516 23940
rect 5516 23846 5572 23884
rect 5740 23604 5796 24108
rect 5292 23214 5294 23266
rect 5346 23214 5348 23266
rect 5292 23202 5348 23214
rect 5404 23548 5796 23604
rect 5852 24052 5908 24062
rect 4956 21746 5012 21756
rect 5068 23100 5236 23156
rect 4956 21588 5012 21598
rect 4284 21362 4340 21374
rect 4284 21310 4286 21362
rect 4338 21310 4340 21362
rect 3612 20972 4228 21028
rect 3052 20802 3108 20972
rect 3164 20916 3220 20926
rect 3164 20822 3220 20860
rect 3052 20750 3054 20802
rect 3106 20750 3108 20802
rect 3052 20738 3108 20750
rect 3612 20802 3668 20814
rect 3612 20750 3614 20802
rect 3666 20750 3668 20802
rect 3612 20188 3668 20750
rect 3804 20412 4068 20422
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 3804 20346 4068 20356
rect 3276 20132 3668 20188
rect 3276 20130 3332 20132
rect 3276 20078 3278 20130
rect 3330 20078 3332 20130
rect 3276 20066 3332 20078
rect 3388 19572 3444 19582
rect 3388 19346 3444 19516
rect 3388 19294 3390 19346
rect 3442 19294 3444 19346
rect 3052 19122 3108 19134
rect 3052 19070 3054 19122
rect 3106 19070 3108 19122
rect 3052 18564 3108 19070
rect 3388 18788 3444 19294
rect 3804 18844 4068 18854
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 3804 18778 4068 18788
rect 3388 18722 3444 18732
rect 3052 18498 3108 18508
rect 3836 18564 3892 18574
rect 3164 18226 3220 18238
rect 3164 18174 3166 18226
rect 3218 18174 3220 18226
rect 2940 17836 3108 17892
rect 2828 17054 2830 17106
rect 2882 17054 2884 17106
rect 2828 17042 2884 17054
rect 2940 17668 2996 17678
rect 2940 16322 2996 17612
rect 2940 16270 2942 16322
rect 2994 16270 2996 16322
rect 2940 16258 2996 16270
rect 2828 16212 2884 16222
rect 2828 15988 2884 16156
rect 2828 15932 2996 15988
rect 2828 15764 2884 15774
rect 2604 15316 2660 15326
rect 2604 15222 2660 15260
rect 2716 15092 2772 15102
rect 2604 12964 2660 12974
rect 2492 12962 2660 12964
rect 2492 12910 2606 12962
rect 2658 12910 2660 12962
rect 2492 12908 2660 12910
rect 2492 12292 2548 12908
rect 2604 12898 2660 12908
rect 2492 12066 2548 12236
rect 2492 12014 2494 12066
rect 2546 12014 2548 12066
rect 2492 12002 2548 12014
rect 2604 12740 2660 12750
rect 2268 11900 2436 11956
rect 2268 9938 2324 11900
rect 2268 9886 2270 9938
rect 2322 9886 2324 9938
rect 2268 9874 2324 9886
rect 2380 11620 2436 11630
rect 2268 9044 2324 9054
rect 2380 9044 2436 11564
rect 2492 10386 2548 10398
rect 2492 10334 2494 10386
rect 2546 10334 2548 10386
rect 2492 10052 2548 10334
rect 2492 9986 2548 9996
rect 2268 9042 2436 9044
rect 2268 8990 2270 9042
rect 2322 8990 2436 9042
rect 2268 8988 2436 8990
rect 2268 8978 2324 8988
rect 2156 8642 2212 8652
rect 2604 8596 2660 12684
rect 2716 11618 2772 15036
rect 2716 11566 2718 11618
rect 2770 11566 2772 11618
rect 2716 11508 2772 11566
rect 2716 11442 2772 11452
rect 2492 8540 2660 8596
rect 2716 10052 2772 10062
rect 2492 8428 2548 8540
rect 2716 8428 2772 9996
rect 2828 9714 2884 15708
rect 2940 10052 2996 15932
rect 3052 15204 3108 17836
rect 3164 16884 3220 18174
rect 3724 17780 3780 17790
rect 3388 17778 3780 17780
rect 3388 17726 3726 17778
rect 3778 17726 3780 17778
rect 3388 17724 3780 17726
rect 3164 16818 3220 16828
rect 3276 17666 3332 17678
rect 3276 17614 3278 17666
rect 3330 17614 3332 17666
rect 3052 15138 3108 15148
rect 3276 14754 3332 17614
rect 3388 16882 3444 17724
rect 3724 17714 3780 17724
rect 3836 17556 3892 18508
rect 3388 16830 3390 16882
rect 3442 16830 3444 16882
rect 3388 16818 3444 16830
rect 3612 17500 3892 17556
rect 3948 17666 4004 17678
rect 3948 17614 3950 17666
rect 4002 17614 4004 17666
rect 3948 17556 4004 17614
rect 3612 16100 3668 17500
rect 3948 17490 4004 17500
rect 3804 17276 4068 17286
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 3804 17210 4068 17220
rect 3836 16996 3892 17006
rect 3836 16902 3892 16940
rect 4060 16324 4116 16334
rect 4172 16324 4228 20972
rect 4284 20020 4340 21310
rect 4464 21196 4728 21206
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4464 21130 4728 21140
rect 4956 20916 5012 21532
rect 4396 20802 4452 20814
rect 4396 20750 4398 20802
rect 4450 20750 4452 20802
rect 4396 20692 4452 20750
rect 4396 20626 4452 20636
rect 4284 19954 4340 19964
rect 4844 20244 4900 20254
rect 4464 19628 4728 19638
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4464 19562 4728 19572
rect 4620 19236 4676 19246
rect 4620 19142 4676 19180
rect 4284 18226 4340 18238
rect 4284 18174 4286 18226
rect 4338 18174 4340 18226
rect 4284 17892 4340 18174
rect 4464 18060 4728 18070
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4464 17994 4728 18004
rect 4284 17826 4340 17836
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 4732 17554 4788 17566
rect 4732 17502 4734 17554
rect 4786 17502 4788 17554
rect 4732 17220 4788 17502
rect 4732 17154 4788 17164
rect 4464 16492 4728 16502
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4464 16426 4728 16436
rect 4060 16322 4172 16324
rect 4060 16270 4062 16322
rect 4114 16270 4172 16322
rect 4060 16268 4172 16270
rect 4060 16258 4116 16268
rect 4172 16230 4228 16268
rect 3612 16006 3668 16044
rect 3804 15708 4068 15718
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 3804 15642 4068 15652
rect 4060 15540 4116 15550
rect 3276 14702 3278 14754
rect 3330 14702 3332 14754
rect 3276 14690 3332 14702
rect 3500 15428 3556 15438
rect 3388 13636 3444 13646
rect 3388 13542 3444 13580
rect 3164 13188 3220 13198
rect 2940 9986 2996 9996
rect 3052 13076 3108 13086
rect 2828 9662 2830 9714
rect 2882 9662 2884 9714
rect 2828 9650 2884 9662
rect 2044 6638 2046 6690
rect 2098 6638 2100 6690
rect 2044 6626 2100 6638
rect 2156 8372 2548 8428
rect 2604 8372 2772 8428
rect 2940 9492 2996 9502
rect 2156 5906 2212 8372
rect 2268 8260 2324 8270
rect 2268 8258 2436 8260
rect 2268 8206 2270 8258
rect 2322 8206 2436 8258
rect 2268 8204 2436 8206
rect 2268 8194 2324 8204
rect 2268 8036 2324 8046
rect 2268 7474 2324 7980
rect 2380 7700 2436 8204
rect 2380 7634 2436 7644
rect 2268 7422 2270 7474
rect 2322 7422 2324 7474
rect 2268 7410 2324 7422
rect 2492 7588 2548 7598
rect 2156 5854 2158 5906
rect 2210 5854 2212 5906
rect 2156 5842 2212 5854
rect 2492 5348 2548 7532
rect 2604 5906 2660 8372
rect 2940 7586 2996 9436
rect 3052 9154 3108 13020
rect 3164 13074 3220 13132
rect 3164 13022 3166 13074
rect 3218 13022 3220 13074
rect 3164 13010 3220 13022
rect 3500 13074 3556 15372
rect 4060 15428 4116 15484
rect 4172 15428 4228 15438
rect 4060 15426 4228 15428
rect 4060 15374 4174 15426
rect 4226 15374 4228 15426
rect 4060 15372 4228 15374
rect 3724 15204 3780 15242
rect 3724 15138 3780 15148
rect 3948 14532 4004 14542
rect 3612 14530 4004 14532
rect 3612 14478 3950 14530
rect 4002 14478 4004 14530
rect 3612 14476 4004 14478
rect 3612 13186 3668 14476
rect 3948 14466 4004 14476
rect 4060 14308 4116 15372
rect 4172 15362 4228 15372
rect 4464 14924 4728 14934
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4464 14858 4728 14868
rect 4172 14756 4228 14766
rect 4172 14642 4228 14700
rect 4172 14590 4174 14642
rect 4226 14590 4228 14642
rect 4172 14578 4228 14590
rect 4284 14532 4340 14542
rect 4284 14438 4340 14476
rect 4732 14308 4788 14318
rect 4060 14252 4228 14308
rect 3804 14140 4068 14150
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 3804 14074 4068 14084
rect 3612 13134 3614 13186
rect 3666 13134 3668 13186
rect 3612 13122 3668 13134
rect 3724 13972 3780 13982
rect 3500 13022 3502 13074
rect 3554 13022 3556 13074
rect 3500 13010 3556 13022
rect 3724 12852 3780 13916
rect 3948 13860 4004 13870
rect 3948 13746 4004 13804
rect 3948 13694 3950 13746
rect 4002 13694 4004 13746
rect 3948 13682 4004 13694
rect 4172 12962 4228 14252
rect 4732 14214 4788 14252
rect 4396 14196 4452 14206
rect 4396 13858 4452 14140
rect 4844 13972 4900 20188
rect 4956 16548 5012 20860
rect 5068 19348 5124 23100
rect 5404 23044 5460 23548
rect 5180 22988 5460 23044
rect 5628 23380 5684 23390
rect 5180 20580 5236 22988
rect 5516 22932 5572 22942
rect 5404 21586 5460 21598
rect 5404 21534 5406 21586
rect 5458 21534 5460 21586
rect 5292 21476 5348 21486
rect 5292 20802 5348 21420
rect 5404 21140 5460 21534
rect 5404 21074 5460 21084
rect 5292 20750 5294 20802
rect 5346 20750 5348 20802
rect 5292 20738 5348 20750
rect 5180 20524 5460 20580
rect 5180 20020 5236 20030
rect 5404 20020 5460 20524
rect 5516 20242 5572 22876
rect 5628 22708 5684 23324
rect 5740 22932 5796 22942
rect 5740 22838 5796 22876
rect 5628 22652 5796 22708
rect 5628 22260 5684 22270
rect 5628 21700 5684 22204
rect 5628 21634 5684 21644
rect 5516 20190 5518 20242
rect 5570 20190 5572 20242
rect 5516 20178 5572 20190
rect 5180 20018 5348 20020
rect 5180 19966 5182 20018
rect 5234 19966 5348 20018
rect 5180 19964 5348 19966
rect 5404 19964 5572 20020
rect 5180 19954 5236 19964
rect 5068 19292 5236 19348
rect 5068 19122 5124 19134
rect 5068 19070 5070 19122
rect 5122 19070 5124 19122
rect 5068 18900 5124 19070
rect 5068 18834 5124 18844
rect 5068 18564 5124 18574
rect 5068 18470 5124 18508
rect 5068 18340 5124 18350
rect 5068 17780 5124 18284
rect 5068 17686 5124 17724
rect 5180 17332 5236 19292
rect 5292 17892 5348 19964
rect 5404 19236 5460 19246
rect 5404 19142 5460 19180
rect 5516 19012 5572 19964
rect 5404 18956 5572 19012
rect 5740 19012 5796 22652
rect 5852 21028 5908 23996
rect 5852 20962 5908 20972
rect 5852 20580 5908 20590
rect 5852 20486 5908 20524
rect 5964 20356 6020 27132
rect 6076 23938 6132 28924
rect 6188 28642 6244 33852
rect 6300 33906 6692 33908
rect 6300 33854 6638 33906
rect 6690 33854 6692 33906
rect 6300 33852 6692 33854
rect 6300 30436 6356 33852
rect 6636 33842 6692 33852
rect 6412 33684 6468 33694
rect 6412 31106 6468 33628
rect 6524 33124 6580 33134
rect 6524 33122 6692 33124
rect 6524 33070 6526 33122
rect 6578 33070 6692 33122
rect 6524 33068 6692 33070
rect 6524 33058 6580 33068
rect 6412 31054 6414 31106
rect 6466 31054 6468 31106
rect 6412 31042 6468 31054
rect 6524 31778 6580 31790
rect 6524 31726 6526 31778
rect 6578 31726 6580 31778
rect 6524 30436 6580 31726
rect 6300 30370 6356 30380
rect 6412 30380 6580 30436
rect 6412 29652 6468 30380
rect 6524 30212 6580 30222
rect 6524 30118 6580 30156
rect 6412 29586 6468 29596
rect 6636 29428 6692 33068
rect 6188 28590 6190 28642
rect 6242 28590 6244 28642
rect 6188 25284 6244 28590
rect 6412 29372 6692 29428
rect 6188 25218 6244 25228
rect 6300 27074 6356 27086
rect 6300 27022 6302 27074
rect 6354 27022 6356 27074
rect 6300 24052 6356 27022
rect 6412 26628 6468 29372
rect 6524 28420 6580 28430
rect 6524 27858 6580 28364
rect 6524 27806 6526 27858
rect 6578 27806 6580 27858
rect 6524 26908 6580 27806
rect 6524 26852 6692 26908
rect 6412 26562 6468 26572
rect 6412 26404 6468 26414
rect 6412 25508 6468 26348
rect 6524 25508 6580 25518
rect 6412 25506 6580 25508
rect 6412 25454 6526 25506
rect 6578 25454 6580 25506
rect 6412 25452 6580 25454
rect 6524 25442 6580 25452
rect 6636 24276 6692 26852
rect 6748 26516 6804 42924
rect 6860 40402 6916 40414
rect 6860 40350 6862 40402
rect 6914 40350 6916 40402
rect 6860 38836 6916 40350
rect 7532 40292 7588 40302
rect 7196 40290 7588 40292
rect 7196 40238 7534 40290
rect 7586 40238 7588 40290
rect 7196 40236 7588 40238
rect 7084 40180 7140 40190
rect 6972 40178 7140 40180
rect 6972 40126 7086 40178
rect 7138 40126 7140 40178
rect 6972 40124 7140 40126
rect 6972 39842 7028 40124
rect 7084 40114 7140 40124
rect 6972 39790 6974 39842
rect 7026 39790 7028 39842
rect 6972 39778 7028 39790
rect 7196 39396 7252 40236
rect 7532 40226 7588 40236
rect 7308 39732 7364 39742
rect 7308 39638 7364 39676
rect 6972 39340 7252 39396
rect 6972 39058 7028 39340
rect 7644 39060 7700 45724
rect 6972 39006 6974 39058
rect 7026 39006 7028 39058
rect 6972 38994 7028 39006
rect 7196 39004 7700 39060
rect 6860 38770 6916 38780
rect 7196 38668 7252 39004
rect 7756 38668 7812 51212
rect 8092 42868 8148 55918
rect 9996 55970 10052 55982
rect 9996 55918 9998 55970
rect 10050 55918 10052 55970
rect 9100 52164 9156 52174
rect 8876 46564 8932 46574
rect 8092 42802 8148 42812
rect 8540 44996 8596 45006
rect 8316 42196 8372 42206
rect 8316 41748 8372 42140
rect 8540 42084 8596 44940
rect 8540 42018 8596 42028
rect 8652 42532 8708 42542
rect 8316 41692 8484 41748
rect 7868 41076 7924 41086
rect 7868 39844 7924 41020
rect 8204 40402 8260 40414
rect 8204 40350 8206 40402
rect 8258 40350 8260 40402
rect 7868 39842 8036 39844
rect 7868 39790 7870 39842
rect 7922 39790 8036 39842
rect 7868 39788 8036 39790
rect 7868 39778 7924 39788
rect 6860 38612 6916 38622
rect 7196 38612 7588 38668
rect 6860 36484 6916 38556
rect 6972 38162 7028 38174
rect 6972 38110 6974 38162
rect 7026 38110 7028 38162
rect 6972 37042 7028 38110
rect 6972 36990 6974 37042
rect 7026 36990 7028 37042
rect 6972 36596 7028 36990
rect 6972 36540 7252 36596
rect 6860 36482 7140 36484
rect 6860 36430 6862 36482
rect 6914 36430 7140 36482
rect 6860 36428 7140 36430
rect 6860 36418 6916 36428
rect 6860 35586 6916 35598
rect 6860 35534 6862 35586
rect 6914 35534 6916 35586
rect 6860 33460 6916 35534
rect 6972 35026 7028 35038
rect 6972 34974 6974 35026
rect 7026 34974 7028 35026
rect 6972 33908 7028 34974
rect 7084 34468 7140 36428
rect 7084 34402 7140 34412
rect 6972 33842 7028 33852
rect 6860 33394 6916 33404
rect 7196 33348 7252 36540
rect 7196 33282 7252 33292
rect 7420 36370 7476 36382
rect 7420 36318 7422 36370
rect 7474 36318 7476 36370
rect 7196 32562 7252 32574
rect 7196 32510 7198 32562
rect 7250 32510 7252 32562
rect 6972 30996 7028 31006
rect 7196 30996 7252 32510
rect 7308 31778 7364 31790
rect 7308 31726 7310 31778
rect 7362 31726 7364 31778
rect 7308 31444 7364 31726
rect 7420 31668 7476 36318
rect 7532 34580 7588 38612
rect 7532 34514 7588 34524
rect 7644 38612 7812 38668
rect 7868 39060 7924 39070
rect 7644 33684 7700 38612
rect 7756 33908 7812 33918
rect 7756 33814 7812 33852
rect 7420 31602 7476 31612
rect 7532 33628 7700 33684
rect 7364 31388 7476 31444
rect 7308 31378 7364 31388
rect 6972 30994 7252 30996
rect 6972 30942 6974 30994
rect 7026 30942 7252 30994
rect 6972 30940 7252 30942
rect 6972 29764 7028 30940
rect 7308 30884 7364 30894
rect 7308 30790 7364 30828
rect 6972 29698 7028 29708
rect 7308 30210 7364 30222
rect 7308 30158 7310 30210
rect 7362 30158 7364 30210
rect 7196 29652 7252 29662
rect 7196 29558 7252 29596
rect 7308 29540 7364 30158
rect 7308 29474 7364 29484
rect 7308 28642 7364 28654
rect 7308 28590 7310 28642
rect 7362 28590 7364 28642
rect 7308 28420 7364 28590
rect 7308 28354 7364 28364
rect 7420 28308 7476 31388
rect 7420 28242 7476 28252
rect 7420 28084 7476 28094
rect 7420 27990 7476 28028
rect 6748 26460 7028 26516
rect 6300 23986 6356 23996
rect 6412 24220 6692 24276
rect 6748 26178 6804 26190
rect 6748 26126 6750 26178
rect 6802 26126 6804 26178
rect 6748 26068 6804 26126
rect 6076 23886 6078 23938
rect 6130 23886 6132 23938
rect 6076 23874 6132 23886
rect 6188 23828 6244 23838
rect 6188 23826 6356 23828
rect 6188 23774 6190 23826
rect 6242 23774 6356 23826
rect 6188 23772 6356 23774
rect 6188 23762 6244 23772
rect 6076 23156 6132 23166
rect 6076 22482 6132 23100
rect 6300 23156 6356 23772
rect 6300 23062 6356 23100
rect 6076 22430 6078 22482
rect 6130 22430 6132 22482
rect 6076 21028 6132 22430
rect 6076 20972 6356 21028
rect 5852 20300 6020 20356
rect 6188 20804 6244 20814
rect 5852 19234 5908 20300
rect 6076 19348 6132 19358
rect 5852 19182 5854 19234
rect 5906 19182 5908 19234
rect 5852 19170 5908 19182
rect 5964 19346 6132 19348
rect 5964 19294 6078 19346
rect 6130 19294 6132 19346
rect 5964 19292 6132 19294
rect 5404 18340 5460 18956
rect 5740 18946 5796 18956
rect 5964 18788 6020 19292
rect 6076 19282 6132 19292
rect 5516 18732 6020 18788
rect 6076 18788 6132 18798
rect 5516 18450 5572 18732
rect 6076 18564 6132 18732
rect 5516 18398 5518 18450
rect 5570 18398 5572 18450
rect 5516 18386 5572 18398
rect 5852 18562 6132 18564
rect 5852 18510 6078 18562
rect 6130 18510 6132 18562
rect 5852 18508 6132 18510
rect 5404 18274 5460 18284
rect 5292 17836 5684 17892
rect 5180 17266 5236 17276
rect 5404 17666 5460 17678
rect 5404 17614 5406 17666
rect 5458 17614 5460 17666
rect 5404 16996 5460 17614
rect 5180 16940 5460 16996
rect 5516 17332 5572 17342
rect 4956 16482 5012 16492
rect 5068 16882 5124 16894
rect 5068 16830 5070 16882
rect 5122 16830 5124 16882
rect 4844 13906 4900 13916
rect 4956 16324 5012 16334
rect 4396 13806 4398 13858
rect 4450 13806 4452 13858
rect 4396 13794 4452 13806
rect 4956 13860 5012 16268
rect 4956 13794 5012 13804
rect 4956 13636 5012 13646
rect 4956 13542 5012 13580
rect 4844 13524 4900 13534
rect 4464 13356 4728 13366
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4464 13290 4728 13300
rect 4620 13076 4676 13086
rect 4844 13076 4900 13468
rect 4620 13074 4900 13076
rect 4620 13022 4622 13074
rect 4674 13022 4900 13074
rect 4620 13020 4900 13022
rect 4620 13010 4676 13020
rect 4172 12910 4174 12962
rect 4226 12910 4228 12962
rect 4172 12898 4228 12910
rect 3500 12796 3780 12852
rect 3164 12180 3220 12190
rect 3164 11394 3220 12124
rect 3164 11342 3166 11394
rect 3218 11342 3220 11394
rect 3164 11330 3220 11342
rect 3052 9102 3054 9154
rect 3106 9102 3108 9154
rect 3052 9090 3108 9102
rect 3276 11284 3332 11294
rect 3276 8932 3332 11228
rect 3052 8876 3332 8932
rect 3052 8370 3108 8876
rect 3052 8318 3054 8370
rect 3106 8318 3108 8370
rect 3052 8306 3108 8318
rect 3164 8708 3220 8718
rect 2940 7534 2942 7586
rect 2994 7534 2996 7586
rect 2940 7522 2996 7534
rect 3164 7028 3220 8652
rect 3500 8260 3556 12796
rect 3804 12572 4068 12582
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 3804 12506 4068 12516
rect 4172 12516 4228 12526
rect 3612 12404 3668 12414
rect 4172 12404 4228 12460
rect 3612 12310 3668 12348
rect 3836 12348 4228 12404
rect 3612 11956 3668 11966
rect 3612 10834 3668 11900
rect 3836 11394 3892 12348
rect 3836 11342 3838 11394
rect 3890 11342 3892 11394
rect 3836 11330 3892 11342
rect 4172 12068 4228 12078
rect 3804 11004 4068 11014
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 3804 10938 4068 10948
rect 3612 10782 3614 10834
rect 3666 10782 3668 10834
rect 3612 10770 3668 10782
rect 3836 9828 3892 9838
rect 3836 9734 3892 9772
rect 3804 9436 4068 9446
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 3804 9370 4068 9380
rect 3836 9044 3892 9054
rect 4172 9044 4228 12012
rect 4464 11788 4728 11798
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4464 11722 4728 11732
rect 4284 11282 4340 11294
rect 4284 11230 4286 11282
rect 4338 11230 4340 11282
rect 4284 11172 4340 11230
rect 4284 11106 4340 11116
rect 4844 11060 4900 13020
rect 5068 12404 5124 16830
rect 5180 16322 5236 16940
rect 5180 16270 5182 16322
rect 5234 16270 5236 16322
rect 5180 16258 5236 16270
rect 5292 16660 5348 16670
rect 5180 15540 5236 15550
rect 5180 15426 5236 15484
rect 5180 15374 5182 15426
rect 5234 15374 5236 15426
rect 5180 14530 5236 15374
rect 5180 14478 5182 14530
rect 5234 14478 5236 14530
rect 5180 14466 5236 14478
rect 5068 12338 5124 12348
rect 5292 12290 5348 16604
rect 5516 16548 5572 17276
rect 5404 16492 5572 16548
rect 5404 15316 5460 16492
rect 5628 16436 5684 17836
rect 5404 15250 5460 15260
rect 5516 16380 5684 16436
rect 5740 16884 5796 16894
rect 5516 15148 5572 16380
rect 5292 12238 5294 12290
rect 5346 12238 5348 12290
rect 5292 12226 5348 12238
rect 5404 15092 5572 15148
rect 5628 15988 5684 15998
rect 5628 15202 5684 15932
rect 5628 15150 5630 15202
rect 5682 15150 5684 15202
rect 5628 15138 5684 15150
rect 5404 11956 5460 15092
rect 5740 14754 5796 16828
rect 5852 16324 5908 18508
rect 6076 18498 6132 18508
rect 5964 18340 6020 18350
rect 5964 17666 6020 18284
rect 6076 17780 6132 17790
rect 6076 17686 6132 17724
rect 5964 17614 5966 17666
rect 6018 17614 6020 17666
rect 5964 17556 6020 17614
rect 5964 17490 6020 17500
rect 5964 17108 6020 17118
rect 6188 17108 6244 20748
rect 5964 17106 6244 17108
rect 5964 17054 5966 17106
rect 6018 17054 6244 17106
rect 5964 17052 6244 17054
rect 5964 17042 6020 17052
rect 5852 16258 5908 16268
rect 5964 16212 6020 16222
rect 5964 16210 6132 16212
rect 5964 16158 5966 16210
rect 6018 16158 6132 16210
rect 5964 16156 6132 16158
rect 5964 16146 6020 16156
rect 5852 16098 5908 16110
rect 5852 16046 5854 16098
rect 5906 16046 5908 16098
rect 5852 15316 5908 16046
rect 5852 15250 5908 15260
rect 5740 14702 5742 14754
rect 5794 14702 5796 14754
rect 5740 14690 5796 14702
rect 5516 13972 5572 13982
rect 5516 13878 5572 13916
rect 5740 13300 5796 13310
rect 5740 13186 5796 13244
rect 5740 13134 5742 13186
rect 5794 13134 5796 13186
rect 5740 13122 5796 13134
rect 6076 12404 6132 16156
rect 6188 16098 6244 16110
rect 6188 16046 6190 16098
rect 6242 16046 6244 16098
rect 6188 14868 6244 16046
rect 6300 15988 6356 20972
rect 6300 15922 6356 15932
rect 6412 15148 6468 24220
rect 6748 24164 6804 26012
rect 6748 24098 6804 24108
rect 6860 25732 6916 25742
rect 6524 24052 6580 24062
rect 6524 23958 6580 23996
rect 6860 23940 6916 25676
rect 6972 25060 7028 26460
rect 7420 26068 7476 26078
rect 7084 25618 7140 25630
rect 7084 25566 7086 25618
rect 7138 25566 7140 25618
rect 7084 25284 7140 25566
rect 7084 25218 7140 25228
rect 6972 25004 7140 25060
rect 6972 24836 7028 24846
rect 6972 24610 7028 24780
rect 6972 24558 6974 24610
rect 7026 24558 7028 24610
rect 6972 24388 7028 24558
rect 6972 24322 7028 24332
rect 6636 23884 6916 23940
rect 6524 21588 6580 21598
rect 6524 21494 6580 21532
rect 6524 20580 6580 20590
rect 6524 19346 6580 20524
rect 6524 19294 6526 19346
rect 6578 19294 6580 19346
rect 6524 19282 6580 19294
rect 6636 19012 6692 23884
rect 7084 23828 7140 25004
rect 7420 24722 7476 26012
rect 7420 24670 7422 24722
rect 7474 24670 7476 24722
rect 7420 24658 7476 24670
rect 6748 23772 7140 23828
rect 7196 23940 7252 23950
rect 6748 19124 6804 23772
rect 7196 23716 7252 23884
rect 6972 23660 7252 23716
rect 6860 23042 6916 23054
rect 6860 22990 6862 23042
rect 6914 22990 6916 23042
rect 6860 22820 6916 22990
rect 6860 22754 6916 22764
rect 6860 21588 6916 21598
rect 6860 20692 6916 21532
rect 6972 21364 7028 23660
rect 7532 23548 7588 33628
rect 7644 33460 7700 33470
rect 7644 33366 7700 33404
rect 7644 32452 7700 32462
rect 7644 32358 7700 32396
rect 7868 31892 7924 39004
rect 7980 38948 8036 39788
rect 8204 39060 8260 40350
rect 8204 38994 8260 39004
rect 7980 38892 8148 38948
rect 7980 38724 8036 38734
rect 7980 38630 8036 38668
rect 8092 38164 8148 38892
rect 8316 38834 8372 38846
rect 8316 38782 8318 38834
rect 8370 38782 8372 38834
rect 8204 38276 8260 38286
rect 8204 38182 8260 38220
rect 7980 38108 8148 38164
rect 7980 36706 8036 38108
rect 8316 38052 8372 38782
rect 8092 37996 8372 38052
rect 8092 37490 8148 37996
rect 8092 37438 8094 37490
rect 8146 37438 8148 37490
rect 8092 37426 8148 37438
rect 7980 36654 7982 36706
rect 8034 36654 8036 36706
rect 7980 35812 8036 36654
rect 7980 35746 8036 35756
rect 8316 35924 8372 35934
rect 8092 35474 8148 35486
rect 8092 35422 8094 35474
rect 8146 35422 8148 35474
rect 8092 34132 8148 35422
rect 8204 34692 8260 34730
rect 8204 34626 8260 34636
rect 8092 34066 8148 34076
rect 8204 34468 8260 34478
rect 8204 34130 8260 34412
rect 8204 34078 8206 34130
rect 8258 34078 8260 34130
rect 8204 33346 8260 34078
rect 8204 33294 8206 33346
rect 8258 33294 8260 33346
rect 7868 31836 8148 31892
rect 8092 31778 8148 31836
rect 8092 31726 8094 31778
rect 8146 31726 8148 31778
rect 7980 31668 8036 31678
rect 7756 29764 7812 29774
rect 7308 23492 7588 23548
rect 7644 28196 7700 28206
rect 7084 23268 7140 23278
rect 7084 21586 7140 23212
rect 7084 21534 7086 21586
rect 7138 21534 7140 21586
rect 7084 21522 7140 21534
rect 7196 22146 7252 22158
rect 7196 22094 7198 22146
rect 7250 22094 7252 22146
rect 6972 21308 7140 21364
rect 6972 20916 7028 20926
rect 6972 20822 7028 20860
rect 6860 20244 6916 20636
rect 6972 20244 7028 20254
rect 6860 20188 6972 20244
rect 6972 20130 7028 20188
rect 6972 20078 6974 20130
rect 7026 20078 7028 20130
rect 6972 20066 7028 20078
rect 7084 19234 7140 21308
rect 7196 20916 7252 22094
rect 7196 20850 7252 20860
rect 7308 20692 7364 23492
rect 7532 22932 7588 22942
rect 7532 21474 7588 22876
rect 7532 21422 7534 21474
rect 7586 21422 7588 21474
rect 7532 21410 7588 21422
rect 7644 21586 7700 28140
rect 7756 26404 7812 29708
rect 7980 28530 8036 31612
rect 8092 30324 8148 31726
rect 8204 31668 8260 33294
rect 8204 31602 8260 31612
rect 8092 30258 8148 30268
rect 8092 29986 8148 29998
rect 8092 29934 8094 29986
rect 8146 29934 8148 29986
rect 8092 29764 8148 29934
rect 8092 29698 8148 29708
rect 7980 28478 7982 28530
rect 8034 28478 8036 28530
rect 7980 28308 8036 28478
rect 7980 28242 8036 28252
rect 8092 28532 8148 28542
rect 8092 27858 8148 28476
rect 8092 27806 8094 27858
rect 8146 27806 8148 27858
rect 8092 27794 8148 27806
rect 8316 27186 8372 35868
rect 8316 27134 8318 27186
rect 8370 27134 8372 27186
rect 8316 27122 8372 27134
rect 7868 27074 7924 27086
rect 7868 27022 7870 27074
rect 7922 27022 7924 27074
rect 7868 26908 7924 27022
rect 8428 26908 8484 41692
rect 8652 38668 8708 42476
rect 8764 39172 8820 39182
rect 8764 38836 8820 39116
rect 8764 38742 8820 38780
rect 8540 38612 8708 38668
rect 8540 32788 8596 38612
rect 8652 37268 8708 37278
rect 8652 35698 8708 37212
rect 8652 35646 8654 35698
rect 8706 35646 8708 35698
rect 8652 35634 8708 35646
rect 8764 36596 8820 36606
rect 8652 35476 8708 35486
rect 8652 34020 8708 35420
rect 8764 34244 8820 36540
rect 8876 34468 8932 46508
rect 9100 45332 9156 52108
rect 9100 45266 9156 45276
rect 9772 42756 9828 42766
rect 8988 40964 9044 40974
rect 8988 40962 9492 40964
rect 8988 40910 8990 40962
rect 9042 40910 9492 40962
rect 8988 40908 9492 40910
rect 8988 40898 9044 40908
rect 9212 40402 9268 40414
rect 9212 40350 9214 40402
rect 9266 40350 9268 40402
rect 8988 39618 9044 39630
rect 8988 39566 8990 39618
rect 9042 39566 9044 39618
rect 8988 38722 9044 39566
rect 8988 38670 8990 38722
rect 9042 38670 9044 38722
rect 8988 38658 9044 38670
rect 9212 38724 9268 40350
rect 9436 38834 9492 40908
rect 9548 39956 9604 39966
rect 9548 39730 9604 39900
rect 9548 39678 9550 39730
rect 9602 39678 9604 39730
rect 9548 39666 9604 39678
rect 9436 38782 9438 38834
rect 9490 38782 9492 38834
rect 9436 38770 9492 38782
rect 9772 38668 9828 42700
rect 9884 42644 9940 42654
rect 9884 39508 9940 42588
rect 9996 39732 10052 55918
rect 10220 55300 10276 55310
rect 10108 41300 10164 41310
rect 10108 41206 10164 41244
rect 9996 39666 10052 39676
rect 9884 39452 10052 39508
rect 9212 38658 9268 38668
rect 9436 38612 9828 38668
rect 9884 38724 9940 38734
rect 9324 37156 9380 37166
rect 9212 37154 9380 37156
rect 9212 37102 9326 37154
rect 9378 37102 9380 37154
rect 9212 37100 9380 37102
rect 9212 35140 9268 37100
rect 9324 37090 9380 37100
rect 9324 35586 9380 35598
rect 9324 35534 9326 35586
rect 9378 35534 9380 35586
rect 9324 35476 9380 35534
rect 9324 35410 9380 35420
rect 9212 35074 9268 35084
rect 9324 35028 9380 35038
rect 8876 34402 8932 34412
rect 9100 34692 9156 34702
rect 8764 34188 8932 34244
rect 8652 33954 8708 33964
rect 8764 34018 8820 34030
rect 8764 33966 8766 34018
rect 8818 33966 8820 34018
rect 8540 32722 8596 32732
rect 8652 33684 8708 33694
rect 8540 30770 8596 30782
rect 8540 30718 8542 30770
rect 8594 30718 8596 30770
rect 8540 30100 8596 30718
rect 8540 30034 8596 30044
rect 8540 29540 8596 29550
rect 8540 29446 8596 29484
rect 8652 27748 8708 33628
rect 8764 32900 8820 33966
rect 8876 33684 8932 34188
rect 9100 34130 9156 34636
rect 9100 34078 9102 34130
rect 9154 34078 9156 34130
rect 9100 34066 9156 34078
rect 8876 33618 8932 33628
rect 9324 33684 9380 34972
rect 9324 33618 9380 33628
rect 8876 33460 8932 33470
rect 9436 33460 9492 38612
rect 8876 33366 8932 33404
rect 9324 33404 9492 33460
rect 9548 38164 9604 38174
rect 8764 32834 8820 32844
rect 8652 27654 8708 27692
rect 8764 32676 8820 32686
rect 7868 26852 8148 26908
rect 8428 26852 8596 26908
rect 7756 26338 7812 26348
rect 7980 26068 8036 26078
rect 7980 25974 8036 26012
rect 7756 25172 7812 25182
rect 7756 24722 7812 25116
rect 7756 24670 7758 24722
rect 7810 24670 7812 24722
rect 7756 24658 7812 24670
rect 7980 24612 8036 24622
rect 8092 24612 8148 26852
rect 8204 25282 8260 25294
rect 8204 25230 8206 25282
rect 8258 25230 8260 25282
rect 8204 24724 8260 25230
rect 8204 24658 8260 24668
rect 8428 24724 8484 24734
rect 8428 24630 8484 24668
rect 7980 24610 8148 24612
rect 7980 24558 7982 24610
rect 8034 24558 8148 24610
rect 7980 24556 8148 24558
rect 7980 24546 8036 24556
rect 8316 24500 8372 24510
rect 7756 23714 7812 23726
rect 7756 23662 7758 23714
rect 7810 23662 7812 23714
rect 7756 23268 7812 23662
rect 7756 23202 7812 23212
rect 7756 22932 7812 22942
rect 7756 22930 8148 22932
rect 7756 22878 7758 22930
rect 7810 22878 8148 22930
rect 7756 22876 8148 22878
rect 7756 22866 7812 22876
rect 7644 21534 7646 21586
rect 7698 21534 7700 21586
rect 7644 21252 7700 21534
rect 7532 21196 7700 21252
rect 7756 21924 7812 21934
rect 7084 19182 7086 19234
rect 7138 19182 7140 19234
rect 7084 19170 7140 19182
rect 7196 20636 7364 20692
rect 7420 20690 7476 20702
rect 7420 20638 7422 20690
rect 7474 20638 7476 20690
rect 6748 19068 6916 19124
rect 6636 18956 6804 19012
rect 6524 18228 6580 18238
rect 6524 18134 6580 18172
rect 6524 17892 6580 17902
rect 6524 17778 6580 17836
rect 6524 17726 6526 17778
rect 6578 17726 6580 17778
rect 6524 17714 6580 17726
rect 6636 15988 6692 15998
rect 6748 15988 6804 18956
rect 6860 18004 6916 19068
rect 6860 17948 7028 18004
rect 6692 15932 6804 15988
rect 6860 16658 6916 16670
rect 6860 16606 6862 16658
rect 6914 16606 6916 16658
rect 6636 15894 6692 15932
rect 6748 15764 6804 15774
rect 6748 15538 6804 15708
rect 6748 15486 6750 15538
rect 6802 15486 6804 15538
rect 6748 15474 6804 15486
rect 6860 15148 6916 16606
rect 6972 16212 7028 17948
rect 6972 16118 7028 16156
rect 7084 15764 7140 15774
rect 7084 15314 7140 15708
rect 7084 15262 7086 15314
rect 7138 15262 7140 15314
rect 7084 15250 7140 15262
rect 6188 14802 6244 14812
rect 6300 15092 6468 15148
rect 6748 15092 6916 15148
rect 6972 15204 7028 15214
rect 6076 12348 6244 12404
rect 5404 11890 5460 11900
rect 5628 12292 5684 12302
rect 5404 11508 5460 11518
rect 5404 11414 5460 11452
rect 5068 11284 5124 11294
rect 5068 11282 5236 11284
rect 5068 11230 5070 11282
rect 5122 11230 5236 11282
rect 5068 11228 5236 11230
rect 5068 11218 5124 11228
rect 4844 11004 5124 11060
rect 4956 10836 5012 10846
rect 4464 10220 4728 10230
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4464 10154 4728 10164
rect 4956 9826 5012 10780
rect 4956 9774 4958 9826
rect 5010 9774 5012 9826
rect 4956 9762 5012 9774
rect 3836 9042 4228 9044
rect 3836 8990 3838 9042
rect 3890 8990 4228 9042
rect 3836 8988 4228 8990
rect 5068 9042 5124 11004
rect 5180 10836 5236 11228
rect 5180 10722 5236 10780
rect 5180 10670 5182 10722
rect 5234 10670 5236 10722
rect 5180 10658 5236 10670
rect 5628 10498 5684 12236
rect 6076 12178 6132 12190
rect 6076 12126 6078 12178
rect 6130 12126 6132 12178
rect 5628 10446 5630 10498
rect 5682 10446 5684 10498
rect 5628 10434 5684 10446
rect 5852 11508 5908 11518
rect 5068 8990 5070 9042
rect 5122 8990 5124 9042
rect 3836 8978 3892 8988
rect 5068 8978 5124 8990
rect 5180 10388 5236 10398
rect 4464 8652 4728 8662
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4464 8586 4728 8596
rect 3612 8260 3668 8270
rect 3500 8258 3668 8260
rect 3500 8206 3614 8258
rect 3666 8206 3668 8258
rect 3500 8204 3668 8206
rect 3612 8194 3668 8204
rect 5068 8036 5124 8046
rect 5068 7942 5124 7980
rect 3804 7868 4068 7878
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 3804 7802 4068 7812
rect 3836 7476 3892 7486
rect 3836 7382 3892 7420
rect 5068 7476 5124 7486
rect 5180 7476 5236 10332
rect 5292 9940 5348 9950
rect 5292 9846 5348 9884
rect 5516 9156 5572 9166
rect 5516 9062 5572 9100
rect 5852 9042 5908 11452
rect 5852 8990 5854 9042
rect 5906 8990 5908 9042
rect 5852 8978 5908 8990
rect 5516 8484 5572 8494
rect 5516 7586 5572 8428
rect 5516 7534 5518 7586
rect 5570 7534 5572 7586
rect 5516 7522 5572 7534
rect 5068 7474 5236 7476
rect 5068 7422 5070 7474
rect 5122 7422 5236 7474
rect 5068 7420 5236 7422
rect 5068 7410 5124 7420
rect 3052 6972 3220 7028
rect 4464 7084 4728 7094
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4464 7018 4728 7028
rect 2604 5854 2606 5906
rect 2658 5854 2660 5906
rect 2604 5842 2660 5854
rect 2828 6466 2884 6478
rect 2828 6414 2830 6466
rect 2882 6414 2884 6466
rect 2828 5908 2884 6414
rect 2828 5842 2884 5852
rect 2604 5348 2660 5358
rect 2492 5346 2660 5348
rect 2492 5294 2606 5346
rect 2658 5294 2660 5346
rect 2492 5292 2660 5294
rect 2604 5282 2660 5292
rect 3052 5236 3108 6972
rect 3836 6690 3892 6702
rect 3836 6638 3838 6690
rect 3890 6638 3892 6690
rect 3836 6580 3892 6638
rect 3836 6514 3892 6524
rect 3500 6468 3556 6478
rect 3164 5796 3220 5806
rect 3164 5702 3220 5740
rect 3164 5236 3220 5246
rect 3052 5234 3220 5236
rect 3052 5182 3166 5234
rect 3218 5182 3220 5234
rect 3052 5180 3220 5182
rect 3164 5170 3220 5180
rect 3500 5234 3556 6412
rect 3804 6300 4068 6310
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 3804 6234 4068 6244
rect 6076 6132 6132 12126
rect 6188 10276 6244 12348
rect 6188 10210 6244 10220
rect 6188 8372 6244 8382
rect 6188 8278 6244 8316
rect 6076 6066 6132 6076
rect 4464 5516 4728 5526
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4464 5450 4728 5460
rect 3500 5182 3502 5234
rect 3554 5182 3556 5234
rect 3500 5170 3556 5182
rect 2044 5124 2100 5134
rect 1932 5122 2100 5124
rect 1932 5070 2046 5122
rect 2098 5070 2100 5122
rect 1932 5068 2100 5070
rect 2044 5058 2100 5068
rect 4060 5124 4116 5134
rect 4060 5030 4116 5068
rect 3804 4732 4068 4742
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 3804 4666 4068 4676
rect 1596 2046 1598 2098
rect 1650 2046 1652 2098
rect 1596 2034 1652 2046
rect 2044 4340 2100 4350
rect 924 1586 980 1596
rect 700 644 756 654
rect 700 112 756 588
rect 2044 112 2100 4284
rect 2268 4228 2324 4238
rect 2268 4134 2324 4172
rect 4464 3948 4728 3958
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4464 3882 4728 3892
rect 2268 3556 2324 3566
rect 2268 3462 2324 3500
rect 6300 3388 6356 15092
rect 6412 14644 6468 14654
rect 6412 12850 6468 14588
rect 6412 12798 6414 12850
rect 6466 12798 6468 12850
rect 6412 12786 6468 12798
rect 6412 12180 6468 12190
rect 6412 12068 6468 12124
rect 6524 12068 6580 12078
rect 6412 12066 6580 12068
rect 6412 12014 6526 12066
rect 6578 12014 6580 12066
rect 6412 12012 6580 12014
rect 6412 9828 6468 12012
rect 6524 12002 6580 12012
rect 6748 12068 6804 15092
rect 6860 14644 6916 14654
rect 6860 14550 6916 14588
rect 6972 13858 7028 15148
rect 6972 13806 6974 13858
rect 7026 13806 7028 13858
rect 6972 12404 7028 13806
rect 6972 12338 7028 12348
rect 7084 15092 7140 15102
rect 7084 12180 7140 15036
rect 7196 13524 7252 20636
rect 7308 20020 7364 20030
rect 7308 19926 7364 19964
rect 7420 19684 7476 20638
rect 7532 20132 7588 21196
rect 7756 21028 7812 21868
rect 8092 21586 8148 22876
rect 8092 21534 8094 21586
rect 8146 21534 8148 21586
rect 8092 21522 8148 21534
rect 7532 20066 7588 20076
rect 7644 20972 7812 21028
rect 7476 19628 7588 19684
rect 7420 19618 7476 19628
rect 7308 19236 7364 19246
rect 7308 19234 7476 19236
rect 7308 19182 7310 19234
rect 7362 19182 7476 19234
rect 7308 19180 7476 19182
rect 7308 19170 7364 19180
rect 7308 17666 7364 17678
rect 7308 17614 7310 17666
rect 7362 17614 7364 17666
rect 7308 17220 7364 17614
rect 7308 17154 7364 17164
rect 7420 16324 7476 19180
rect 7420 16258 7476 16268
rect 7532 16100 7588 19628
rect 7644 18450 7700 20972
rect 7980 20804 8036 20814
rect 7756 20244 7812 20254
rect 7756 19796 7812 20188
rect 7868 20132 7924 20142
rect 7868 20018 7924 20076
rect 7868 19966 7870 20018
rect 7922 19966 7924 20018
rect 7868 19954 7924 19966
rect 7980 19906 8036 20748
rect 7980 19854 7982 19906
rect 8034 19854 8036 19906
rect 7980 19842 8036 19854
rect 7756 19740 7924 19796
rect 7644 18398 7646 18450
rect 7698 18398 7700 18450
rect 7644 18386 7700 18398
rect 7532 15540 7588 16044
rect 7420 15484 7588 15540
rect 7756 17444 7812 17454
rect 7756 16996 7812 17388
rect 7308 15202 7364 15214
rect 7308 15150 7310 15202
rect 7362 15150 7364 15202
rect 7308 14532 7364 15150
rect 7420 15204 7476 15484
rect 7420 15138 7476 15148
rect 7532 15316 7588 15326
rect 7308 14466 7364 14476
rect 7420 14980 7476 14990
rect 7308 14308 7364 14318
rect 7308 14214 7364 14252
rect 7420 13636 7476 14924
rect 7532 14532 7588 15260
rect 7756 15314 7812 16940
rect 7868 15428 7924 19740
rect 8204 19234 8260 19246
rect 8204 19182 8206 19234
rect 8258 19182 8260 19234
rect 8204 19012 8260 19182
rect 8204 18946 8260 18956
rect 8316 18788 8372 24444
rect 8540 22484 8596 26852
rect 8540 22418 8596 22428
rect 8652 25508 8708 25518
rect 8540 21476 8596 21486
rect 8540 21382 8596 21420
rect 8428 20916 8484 20926
rect 8428 20018 8484 20860
rect 8428 19966 8430 20018
rect 8482 19966 8484 20018
rect 8428 19954 8484 19966
rect 8652 19236 8708 25452
rect 8316 18722 8372 18732
rect 8540 19180 8708 19236
rect 8316 18562 8372 18574
rect 8316 18510 8318 18562
rect 8370 18510 8372 18562
rect 8092 18340 8148 18350
rect 8092 16770 8148 18284
rect 8204 17668 8260 17678
rect 8204 17574 8260 17612
rect 8092 16718 8094 16770
rect 8146 16718 8148 16770
rect 8092 16706 8148 16718
rect 8204 16884 8260 16894
rect 8204 16322 8260 16828
rect 8204 16270 8206 16322
rect 8258 16270 8260 16322
rect 8204 16258 8260 16270
rect 8092 15988 8148 15998
rect 7868 15362 7924 15372
rect 7980 15876 8036 15886
rect 7756 15262 7758 15314
rect 7810 15262 7812 15314
rect 7644 15204 7700 15242
rect 7644 15138 7700 15148
rect 7756 15092 7812 15262
rect 7980 15148 8036 15820
rect 8092 15316 8148 15932
rect 8316 15540 8372 18510
rect 8316 15474 8372 15484
rect 8428 16882 8484 16894
rect 8428 16830 8430 16882
rect 8482 16830 8484 16882
rect 8316 15316 8372 15326
rect 8092 15314 8372 15316
rect 8092 15262 8318 15314
rect 8370 15262 8372 15314
rect 8092 15260 8372 15262
rect 8316 15250 8372 15260
rect 7756 15026 7812 15036
rect 7868 15092 8036 15148
rect 7756 14644 7812 14654
rect 7532 14476 7700 14532
rect 7420 13542 7476 13580
rect 7532 14306 7588 14318
rect 7532 14254 7534 14306
rect 7586 14254 7588 14306
rect 7196 13458 7252 13468
rect 6972 12124 7140 12180
rect 7196 13188 7252 13198
rect 6972 12068 7028 12124
rect 6748 12002 6804 12012
rect 6860 12012 7028 12068
rect 6524 11732 6580 11742
rect 6524 10724 6580 11676
rect 6636 11508 6692 11518
rect 6636 11414 6692 11452
rect 6524 10668 6692 10724
rect 6524 10500 6580 10668
rect 6524 10434 6580 10444
rect 6524 10052 6580 10062
rect 6524 9958 6580 9996
rect 6412 9772 6580 9828
rect 6412 9156 6468 9166
rect 6412 9062 6468 9100
rect 6524 5012 6580 9772
rect 6636 8258 6692 10668
rect 6748 10500 6804 10510
rect 6748 10406 6804 10444
rect 6860 9380 6916 12012
rect 6972 11508 7028 11518
rect 6972 10500 7028 11452
rect 7084 11508 7140 11518
rect 7196 11508 7252 13132
rect 7420 12962 7476 12974
rect 7420 12910 7422 12962
rect 7474 12910 7476 12962
rect 7420 12628 7476 12910
rect 7420 12562 7476 12572
rect 7308 12066 7364 12078
rect 7308 12014 7310 12066
rect 7362 12014 7364 12066
rect 7308 11956 7364 12014
rect 7308 11890 7364 11900
rect 7532 11618 7588 14254
rect 7644 13188 7700 14476
rect 7756 14530 7812 14588
rect 7756 14478 7758 14530
rect 7810 14478 7812 14530
rect 7756 14466 7812 14478
rect 7868 13412 7924 15092
rect 7644 13122 7700 13132
rect 7756 13356 7924 13412
rect 7980 14530 8036 14542
rect 7980 14478 7982 14530
rect 8034 14478 8036 14530
rect 7532 11566 7534 11618
rect 7586 11566 7588 11618
rect 7532 11554 7588 11566
rect 7084 11506 7252 11508
rect 7084 11454 7086 11506
rect 7138 11454 7252 11506
rect 7084 11452 7252 11454
rect 7084 11442 7140 11452
rect 7308 11394 7364 11406
rect 7308 11342 7310 11394
rect 7362 11342 7364 11394
rect 7196 10948 7252 10958
rect 7196 10834 7252 10892
rect 7196 10782 7198 10834
rect 7250 10782 7252 10834
rect 7196 10770 7252 10782
rect 6972 10444 7140 10500
rect 7084 10164 7140 10444
rect 6860 9314 6916 9324
rect 6972 10052 7028 10062
rect 6972 9042 7028 9996
rect 7084 9938 7140 10108
rect 7084 9886 7086 9938
rect 7138 9886 7140 9938
rect 7084 9874 7140 9886
rect 7308 9826 7364 11342
rect 7756 11394 7812 13356
rect 7868 13188 7924 13198
rect 7980 13188 8036 14478
rect 8204 14532 8260 14542
rect 8204 14438 8260 14476
rect 8092 14418 8148 14430
rect 8092 14366 8094 14418
rect 8146 14366 8148 14418
rect 8092 13748 8148 14366
rect 8428 14420 8484 16830
rect 8540 16436 8596 19180
rect 8764 19124 8820 32620
rect 8876 32340 8932 32350
rect 8876 32246 8932 32284
rect 9100 31780 9156 31790
rect 9100 30994 9156 31724
rect 9100 30942 9102 30994
rect 9154 30942 9156 30994
rect 8876 30210 8932 30222
rect 8876 30158 8878 30210
rect 8930 30158 8932 30210
rect 8876 28420 8932 30158
rect 9100 30212 9156 30942
rect 9100 30146 9156 30156
rect 8988 29204 9044 29214
rect 8988 29202 9156 29204
rect 8988 29150 8990 29202
rect 9042 29150 9156 29202
rect 8988 29148 9156 29150
rect 8988 29138 9044 29148
rect 9100 28756 9156 29148
rect 9100 28690 9156 28700
rect 8876 28354 8932 28364
rect 9324 26908 9380 33404
rect 9436 33236 9492 33246
rect 9548 33236 9604 38108
rect 9660 37938 9716 37950
rect 9660 37886 9662 37938
rect 9714 37886 9716 37938
rect 9660 37268 9716 37886
rect 9660 37202 9716 37212
rect 9660 34916 9716 34926
rect 9660 34914 9828 34916
rect 9660 34862 9662 34914
rect 9714 34862 9828 34914
rect 9660 34860 9828 34862
rect 9660 34850 9716 34860
rect 9660 34130 9716 34142
rect 9660 34078 9662 34130
rect 9714 34078 9716 34130
rect 9660 34020 9716 34078
rect 9660 33954 9716 33964
rect 9772 34018 9828 34860
rect 9772 33966 9774 34018
rect 9826 33966 9828 34018
rect 9772 33954 9828 33966
rect 9436 33234 9604 33236
rect 9436 33182 9438 33234
rect 9490 33182 9604 33234
rect 9436 33180 9604 33182
rect 9660 33684 9716 33694
rect 9436 33170 9492 33180
rect 9660 31890 9716 33628
rect 9884 32788 9940 38668
rect 9996 34802 10052 39452
rect 10108 39060 10164 39070
rect 10108 38836 10164 39004
rect 10108 38742 10164 38780
rect 10220 36706 10276 55244
rect 11452 55188 11508 57344
rect 12796 56644 12852 57344
rect 14140 56756 14196 57344
rect 14140 56700 14644 56756
rect 12796 56588 13076 56644
rect 13020 56306 13076 56588
rect 13020 56254 13022 56306
rect 13074 56254 13076 56306
rect 13020 56242 13076 56254
rect 14588 56306 14644 56700
rect 14588 56254 14590 56306
rect 14642 56254 14644 56306
rect 14588 56242 14644 56254
rect 15484 56308 15540 57344
rect 16828 57204 16884 57344
rect 16828 57148 16996 57204
rect 15484 56242 15540 56252
rect 16492 56308 16548 56318
rect 16492 56214 16548 56252
rect 11452 55122 11508 55132
rect 11564 55970 11620 55982
rect 11564 55918 11566 55970
rect 11618 55918 11620 55970
rect 11564 54516 11620 55918
rect 14028 55972 14084 55982
rect 14028 55878 14084 55916
rect 15596 55970 15652 55982
rect 15596 55918 15598 55970
rect 15650 55918 15652 55970
rect 14700 55860 14756 55870
rect 12796 55298 12852 55310
rect 12796 55246 12798 55298
rect 12850 55246 12852 55298
rect 11900 55188 11956 55198
rect 11900 55094 11956 55132
rect 11564 54450 11620 54460
rect 11900 54292 11956 54302
rect 11116 53172 11172 53182
rect 10892 52388 10948 52398
rect 10780 43652 10836 43662
rect 10668 41186 10724 41198
rect 10668 41134 10670 41186
rect 10722 41134 10724 41186
rect 10444 40402 10500 40414
rect 10444 40350 10446 40402
rect 10498 40350 10500 40402
rect 10444 39396 10500 40350
rect 10444 39330 10500 39340
rect 10556 39506 10612 39518
rect 10556 39454 10558 39506
rect 10610 39454 10612 39506
rect 10220 36654 10222 36706
rect 10274 36654 10276 36706
rect 10220 36642 10276 36654
rect 10444 38612 10500 38622
rect 9996 34750 9998 34802
rect 10050 34750 10052 34802
rect 9996 34738 10052 34750
rect 10444 34804 10500 38556
rect 10556 36706 10612 39454
rect 10668 37380 10724 41134
rect 10668 37314 10724 37324
rect 10556 36654 10558 36706
rect 10610 36654 10612 36706
rect 10556 36642 10612 36654
rect 10220 34132 10276 34142
rect 10220 34038 10276 34076
rect 10332 33348 10388 33358
rect 9660 31838 9662 31890
rect 9714 31838 9716 31890
rect 9660 31826 9716 31838
rect 9772 32732 9940 32788
rect 10108 33346 10388 33348
rect 10108 33294 10334 33346
rect 10386 33294 10388 33346
rect 10108 33292 10388 33294
rect 9660 30212 9716 30222
rect 9436 30098 9492 30110
rect 9436 30046 9438 30098
rect 9490 30046 9492 30098
rect 9436 29988 9492 30046
rect 9436 29922 9492 29932
rect 9548 28530 9604 28542
rect 9548 28478 9550 28530
rect 9602 28478 9604 28530
rect 9548 28084 9604 28478
rect 9548 28018 9604 28028
rect 9548 27748 9604 27758
rect 8988 26852 9044 26862
rect 9324 26852 9492 26908
rect 8988 26850 9156 26852
rect 8988 26798 8990 26850
rect 9042 26798 9156 26850
rect 8988 26796 9156 26798
rect 8988 26786 9044 26796
rect 9100 26292 9156 26796
rect 9324 26292 9380 26302
rect 9100 26290 9380 26292
rect 9100 26238 9326 26290
rect 9378 26238 9380 26290
rect 9100 26236 9380 26238
rect 9324 26226 9380 26236
rect 8988 26180 9044 26190
rect 8988 26178 9156 26180
rect 8988 26126 8990 26178
rect 9042 26126 9156 26178
rect 8988 26124 9156 26126
rect 8988 26114 9044 26124
rect 8988 25506 9044 25518
rect 8988 25454 8990 25506
rect 9042 25454 9044 25506
rect 8988 25396 9044 25454
rect 8988 25330 9044 25340
rect 8876 25284 8932 25294
rect 8876 23042 8932 25228
rect 8876 22990 8878 23042
rect 8930 22990 8932 23042
rect 8876 22978 8932 22990
rect 8988 25060 9044 25070
rect 8988 21812 9044 25004
rect 8876 21756 9044 21812
rect 8876 21252 8932 21756
rect 9100 21700 9156 26124
rect 9436 25956 9492 26852
rect 9324 25900 9492 25956
rect 9324 24948 9380 25900
rect 9324 24882 9380 24892
rect 9548 25730 9604 27692
rect 9660 27636 9716 30156
rect 9772 27860 9828 32732
rect 9884 32562 9940 32574
rect 9884 32510 9886 32562
rect 9938 32510 9940 32562
rect 9884 31668 9940 32510
rect 9884 31602 9940 31612
rect 10108 31220 10164 33292
rect 10332 33282 10388 33292
rect 10332 32340 10388 32350
rect 10444 32340 10500 34748
rect 10668 35140 10724 35150
rect 10668 34132 10724 35084
rect 10780 34356 10836 43596
rect 10892 41972 10948 52332
rect 10892 41906 10948 41916
rect 10892 41300 10948 41310
rect 10892 40290 10948 41244
rect 10892 40238 10894 40290
rect 10946 40238 10948 40290
rect 10892 38612 10948 40238
rect 11004 38834 11060 38846
rect 11004 38782 11006 38834
rect 11058 38782 11060 38834
rect 11004 38724 11060 38782
rect 11004 38658 11060 38668
rect 10892 38546 10948 38556
rect 10892 36482 10948 36494
rect 10892 36430 10894 36482
rect 10946 36430 10948 36482
rect 10892 34916 10948 36430
rect 11116 35364 11172 53116
rect 11788 41188 11844 41198
rect 11788 41094 11844 41132
rect 11788 39508 11844 39518
rect 11788 38834 11844 39452
rect 11788 38782 11790 38834
rect 11842 38782 11844 38834
rect 11788 38770 11844 38782
rect 11788 37268 11844 37278
rect 11788 35810 11844 37212
rect 11788 35758 11790 35810
rect 11842 35758 11844 35810
rect 11788 35746 11844 35758
rect 11116 35298 11172 35308
rect 10892 34822 10948 34860
rect 10780 34300 11396 34356
rect 10780 34132 10836 34142
rect 10668 34130 10836 34132
rect 10668 34078 10782 34130
rect 10834 34078 10836 34130
rect 10668 34076 10836 34078
rect 10780 34066 10836 34076
rect 11004 34130 11060 34142
rect 11004 34078 11006 34130
rect 11058 34078 11060 34130
rect 10332 32338 10500 32340
rect 10332 32286 10334 32338
rect 10386 32286 10500 32338
rect 10332 32284 10500 32286
rect 10892 33458 10948 33470
rect 10892 33406 10894 33458
rect 10946 33406 10948 33458
rect 10892 33348 10948 33406
rect 9884 31164 10164 31220
rect 10220 31778 10276 31790
rect 10220 31726 10222 31778
rect 10274 31726 10276 31778
rect 10220 31220 10276 31726
rect 10332 31444 10388 32284
rect 10892 32228 10948 33292
rect 10892 32162 10948 32172
rect 10668 31668 10724 31678
rect 10668 31574 10724 31612
rect 10332 31388 10836 31444
rect 9884 29988 9940 31164
rect 10220 31154 10276 31164
rect 9996 30996 10052 31006
rect 9996 30902 10052 30940
rect 10556 30996 10612 31006
rect 10556 30902 10612 30940
rect 9884 29922 9940 29932
rect 10108 30884 10164 30894
rect 10108 29650 10164 30828
rect 10108 29598 10110 29650
rect 10162 29598 10164 29650
rect 10108 29586 10164 29598
rect 10332 30660 10388 30670
rect 9884 28756 9940 28766
rect 9940 28700 10164 28756
rect 9884 28662 9940 28700
rect 9772 27804 9940 27860
rect 9772 27636 9828 27646
rect 9660 27634 9828 27636
rect 9660 27582 9774 27634
rect 9826 27582 9828 27634
rect 9660 27580 9828 27582
rect 9772 27570 9828 27580
rect 9884 26908 9940 27804
rect 10108 27300 10164 28700
rect 10108 27206 10164 27244
rect 9548 25678 9550 25730
rect 9602 25678 9604 25730
rect 9212 24722 9268 24734
rect 9212 24670 9214 24722
rect 9266 24670 9268 24722
rect 9212 24612 9268 24670
rect 9212 24276 9268 24556
rect 9212 24210 9268 24220
rect 9548 23548 9604 25678
rect 9436 23492 9604 23548
rect 9772 26852 9940 26908
rect 9436 23380 9492 23492
rect 9212 23324 9492 23380
rect 9212 22484 9268 23324
rect 9660 23268 9716 23278
rect 9324 23154 9380 23166
rect 9324 23102 9326 23154
rect 9378 23102 9380 23154
rect 9324 22820 9380 23102
rect 9324 22754 9380 22764
rect 9436 22932 9492 22942
rect 9212 22428 9380 22484
rect 8876 21186 8932 21196
rect 8988 21644 9156 21700
rect 8876 20804 8932 20814
rect 8876 20710 8932 20748
rect 8652 19068 8820 19124
rect 8652 18004 8708 19068
rect 8764 18340 8820 18350
rect 8764 18246 8820 18284
rect 8652 17948 8820 18004
rect 8540 16370 8596 16380
rect 8652 17668 8708 17678
rect 8428 14354 8484 14364
rect 8092 13682 8148 13692
rect 8204 14308 8260 14318
rect 7868 13186 8036 13188
rect 7868 13134 7870 13186
rect 7922 13134 8036 13186
rect 7868 13132 8036 13134
rect 8092 13188 8148 13198
rect 7868 13122 7924 13132
rect 8092 13076 8148 13132
rect 7980 13020 8148 13076
rect 7980 12962 8036 13020
rect 8204 12964 8260 14252
rect 8652 14084 8708 17612
rect 8764 15202 8820 17948
rect 8876 17780 8932 17790
rect 8876 17686 8932 17724
rect 8988 16996 9044 21644
rect 8988 16930 9044 16940
rect 9100 21476 9156 21486
rect 9100 20018 9156 21420
rect 9100 19966 9102 20018
rect 9154 19966 9156 20018
rect 8988 16770 9044 16782
rect 8988 16718 8990 16770
rect 9042 16718 9044 16770
rect 8876 15874 8932 15886
rect 8876 15822 8878 15874
rect 8930 15822 8932 15874
rect 8876 15316 8932 15822
rect 8876 15250 8932 15260
rect 8764 15150 8766 15202
rect 8818 15150 8820 15202
rect 8764 14980 8820 15150
rect 8764 14914 8820 14924
rect 8876 14644 8932 14654
rect 8876 14550 8932 14588
rect 8764 14532 8820 14542
rect 8764 14438 8820 14476
rect 8428 14028 8708 14084
rect 8428 13636 8484 14028
rect 8540 13860 8596 13870
rect 8540 13766 8596 13804
rect 8988 13636 9044 16718
rect 9100 15652 9156 19966
rect 9212 17668 9268 17678
rect 9212 16996 9268 17612
rect 9324 17556 9380 22428
rect 9436 20914 9492 22876
rect 9548 22820 9604 22830
rect 9548 22370 9604 22764
rect 9548 22318 9550 22370
rect 9602 22318 9604 22370
rect 9548 21364 9604 22318
rect 9548 21298 9604 21308
rect 9436 20862 9438 20914
rect 9490 20862 9492 20914
rect 9436 20850 9492 20862
rect 9436 19572 9492 19582
rect 9436 19234 9492 19516
rect 9436 19182 9438 19234
rect 9490 19182 9492 19234
rect 9436 18340 9492 19182
rect 9436 18274 9492 18284
rect 9660 18116 9716 23212
rect 9436 18060 9716 18116
rect 9436 17778 9492 18060
rect 9436 17726 9438 17778
rect 9490 17726 9492 17778
rect 9436 17714 9492 17726
rect 9324 17500 9604 17556
rect 9212 16098 9268 16940
rect 9324 16884 9380 16894
rect 9324 16790 9380 16828
rect 9212 16046 9214 16098
rect 9266 16046 9268 16098
rect 9212 16034 9268 16046
rect 9324 16212 9380 16222
rect 9212 15876 9268 15886
rect 9212 15782 9268 15820
rect 9100 15596 9268 15652
rect 9100 15204 9156 15214
rect 9100 14754 9156 15148
rect 9100 14702 9102 14754
rect 9154 14702 9156 14754
rect 9100 14690 9156 14702
rect 9212 14756 9268 15596
rect 9324 15148 9380 16156
rect 9548 15204 9604 17500
rect 9324 15092 9492 15148
rect 9212 14690 9268 14700
rect 9324 14868 9380 14878
rect 9324 14642 9380 14812
rect 9324 14590 9326 14642
rect 9378 14590 9380 14642
rect 9324 14578 9380 14590
rect 9324 13860 9380 13870
rect 9324 13746 9380 13804
rect 9324 13694 9326 13746
rect 9378 13694 9380 13746
rect 9324 13682 9380 13694
rect 8428 13580 8932 13636
rect 8764 13412 8820 13422
rect 7980 12910 7982 12962
rect 8034 12910 8036 12962
rect 7980 12898 8036 12910
rect 8092 12908 8260 12964
rect 8316 13188 8372 13198
rect 7868 12740 7924 12750
rect 8092 12740 8148 12908
rect 7868 12738 8148 12740
rect 7868 12686 7870 12738
rect 7922 12686 8148 12738
rect 7868 12684 8148 12686
rect 8204 12740 8260 12750
rect 7868 12674 7924 12684
rect 7756 11342 7758 11394
rect 7810 11342 7812 11394
rect 7756 11330 7812 11342
rect 7644 11172 7700 11182
rect 7980 11172 8036 12684
rect 8204 12646 8260 12684
rect 8316 12068 8372 13132
rect 8316 12002 8372 12012
rect 8428 13076 8484 13086
rect 7644 11170 8036 11172
rect 7644 11118 7646 11170
rect 7698 11118 8036 11170
rect 7644 11116 8036 11118
rect 8092 11954 8148 11966
rect 8092 11902 8094 11954
rect 8146 11902 8148 11954
rect 7644 11106 7700 11116
rect 8092 10948 8148 11902
rect 8316 11844 8372 11854
rect 8316 11618 8372 11788
rect 8316 11566 8318 11618
rect 8370 11566 8372 11618
rect 8316 11554 8372 11566
rect 8204 11508 8260 11518
rect 8204 11414 8260 11452
rect 8316 11284 8372 11294
rect 8316 11172 8372 11228
rect 8092 10882 8148 10892
rect 8204 11116 8372 11172
rect 7980 10724 8036 10734
rect 7980 10630 8036 10668
rect 7420 10610 7476 10622
rect 7420 10558 7422 10610
rect 7474 10558 7476 10610
rect 7420 10050 7476 10558
rect 7756 10610 7812 10622
rect 7756 10558 7758 10610
rect 7810 10558 7812 10610
rect 7756 10500 7812 10558
rect 7868 10612 7924 10622
rect 7868 10518 7924 10556
rect 7756 10434 7812 10444
rect 8092 10388 8148 10398
rect 8092 10294 8148 10332
rect 8204 10276 8260 11116
rect 7644 10164 7700 10174
rect 7420 9998 7422 10050
rect 7474 9998 7476 10050
rect 7420 9986 7476 9998
rect 7532 10052 7588 10062
rect 7308 9774 7310 9826
rect 7362 9774 7364 9826
rect 7308 9716 7364 9774
rect 7532 9826 7588 9996
rect 7532 9774 7534 9826
rect 7586 9774 7588 9826
rect 7532 9762 7588 9774
rect 6972 8990 6974 9042
rect 7026 8990 7028 9042
rect 6972 8978 7028 8990
rect 7084 9660 7364 9716
rect 6636 8206 6638 8258
rect 6690 8206 6692 8258
rect 6636 8194 6692 8206
rect 6860 8372 6916 8382
rect 6860 7474 6916 8316
rect 7084 8260 7140 9660
rect 7308 9380 7364 9390
rect 7308 9042 7364 9324
rect 7420 9156 7476 9166
rect 7420 9062 7476 9100
rect 7308 8990 7310 9042
rect 7362 8990 7364 9042
rect 7308 8978 7364 8990
rect 7532 9044 7588 9054
rect 7644 9044 7700 10108
rect 7868 9940 7924 9950
rect 7868 9826 7924 9884
rect 7868 9774 7870 9826
rect 7922 9774 7924 9826
rect 7868 9762 7924 9774
rect 7532 9042 8036 9044
rect 7532 8990 7534 9042
rect 7586 8990 8036 9042
rect 7532 8988 8036 8990
rect 7532 8978 7588 8988
rect 7196 8708 7252 8718
rect 7196 8370 7252 8652
rect 7196 8318 7198 8370
rect 7250 8318 7252 8370
rect 7196 8306 7252 8318
rect 7980 8372 8036 8988
rect 8092 9042 8148 9054
rect 8092 8990 8094 9042
rect 8146 8990 8148 9042
rect 8092 8596 8148 8990
rect 8092 8530 8148 8540
rect 8092 8372 8148 8382
rect 7980 8370 8148 8372
rect 7980 8318 8094 8370
rect 8146 8318 8148 8370
rect 7980 8316 8148 8318
rect 8092 8306 8148 8316
rect 8204 8370 8260 10220
rect 8204 8318 8206 8370
rect 8258 8318 8260 8370
rect 8204 8306 8260 8318
rect 8316 10164 8372 10174
rect 7084 8194 7140 8204
rect 7756 8148 7812 8158
rect 7756 8054 7812 8092
rect 8204 8036 8260 8046
rect 8316 8036 8372 10108
rect 8428 8484 8484 13020
rect 8764 12178 8820 13356
rect 8876 12962 8932 13580
rect 8988 13634 9156 13636
rect 8988 13582 8990 13634
rect 9042 13582 9156 13634
rect 8988 13580 9156 13582
rect 8988 13570 9044 13580
rect 8876 12910 8878 12962
rect 8930 12910 8932 12962
rect 8876 12898 8932 12910
rect 8764 12126 8766 12178
rect 8818 12126 8820 12178
rect 8764 12114 8820 12126
rect 8876 12738 8932 12750
rect 8876 12686 8878 12738
rect 8930 12686 8932 12738
rect 8540 12068 8596 12078
rect 8540 11974 8596 12012
rect 8652 12066 8708 12078
rect 8652 12014 8654 12066
rect 8706 12014 8708 12066
rect 8652 11844 8708 12014
rect 8652 11778 8708 11788
rect 8764 11956 8820 11966
rect 8764 10948 8820 11900
rect 8764 10882 8820 10892
rect 8764 10724 8820 10734
rect 8764 10610 8820 10668
rect 8764 10558 8766 10610
rect 8818 10558 8820 10610
rect 8764 10546 8820 10558
rect 8876 9940 8932 12686
rect 9100 12180 9156 13580
rect 9100 12114 9156 12124
rect 9212 12738 9268 12750
rect 9212 12686 9214 12738
rect 9266 12686 9268 12738
rect 8988 12068 9044 12078
rect 8988 11394 9044 12012
rect 9212 11508 9268 12686
rect 8988 11342 8990 11394
rect 9042 11342 9044 11394
rect 8988 10052 9044 11342
rect 9100 11396 9156 11406
rect 9212 11396 9268 11452
rect 9100 11394 9268 11396
rect 9100 11342 9102 11394
rect 9154 11342 9268 11394
rect 9100 11340 9268 11342
rect 9324 12740 9380 12750
rect 9324 11844 9380 12684
rect 9436 12516 9492 15092
rect 9436 12450 9492 12460
rect 9436 12292 9492 12302
rect 9436 12198 9492 12236
rect 9324 11394 9380 11788
rect 9324 11342 9326 11394
rect 9378 11342 9380 11394
rect 9100 11330 9156 11340
rect 9324 11330 9380 11342
rect 9436 11170 9492 11182
rect 9436 11118 9438 11170
rect 9490 11118 9492 11170
rect 8988 9986 9044 9996
rect 9100 11060 9156 11070
rect 8876 9874 8932 9884
rect 9100 9938 9156 11004
rect 9100 9886 9102 9938
rect 9154 9886 9156 9938
rect 9100 9874 9156 9886
rect 9212 10948 9268 10958
rect 8540 8818 8596 8830
rect 8540 8766 8542 8818
rect 8594 8766 8596 8818
rect 8540 8708 8596 8766
rect 8540 8642 8596 8652
rect 8428 8418 8484 8428
rect 8204 8034 8372 8036
rect 8204 7982 8206 8034
rect 8258 7982 8372 8034
rect 8204 7980 8372 7982
rect 8204 7970 8260 7980
rect 7308 7700 7364 7710
rect 7308 7586 7364 7644
rect 7308 7534 7310 7586
rect 7362 7534 7364 7586
rect 7308 7522 7364 7534
rect 6860 7422 6862 7474
rect 6914 7422 6916 7474
rect 6860 7410 6916 7422
rect 7756 6132 7812 6142
rect 7756 6038 7812 6076
rect 9212 6020 9268 10892
rect 9436 10612 9492 11118
rect 9548 10724 9604 15148
rect 9772 17332 9828 26852
rect 9884 26292 9940 26302
rect 9884 26198 9940 26236
rect 10220 26180 10276 26190
rect 9884 26068 9940 26078
rect 9884 19572 9940 26012
rect 9996 26068 10052 26078
rect 9996 26066 10164 26068
rect 9996 26014 9998 26066
rect 10050 26014 10164 26066
rect 9996 26012 10164 26014
rect 9996 26002 10052 26012
rect 9996 25508 10052 25518
rect 9996 24722 10052 25452
rect 9996 24670 9998 24722
rect 10050 24670 10052 24722
rect 9996 24658 10052 24670
rect 10108 24724 10164 26012
rect 10108 24658 10164 24668
rect 10220 24052 10276 26124
rect 10220 23986 10276 23996
rect 10332 24050 10388 30604
rect 10556 30098 10612 30110
rect 10556 30046 10558 30098
rect 10610 30046 10612 30098
rect 10556 29764 10612 30046
rect 10556 29698 10612 29708
rect 10556 28532 10612 28542
rect 10332 23998 10334 24050
rect 10386 23998 10388 24050
rect 10332 23986 10388 23998
rect 10444 28084 10500 28094
rect 10444 27858 10500 28028
rect 10444 27806 10446 27858
rect 10498 27806 10500 27858
rect 10220 23828 10276 23838
rect 10108 23492 10164 23502
rect 9996 22484 10052 22494
rect 10108 22484 10164 23436
rect 10052 22428 10164 22484
rect 9996 22390 10052 22428
rect 10108 20692 10164 22428
rect 10220 20916 10276 23772
rect 10332 23156 10388 23166
rect 10332 23062 10388 23100
rect 10444 22260 10500 27806
rect 10556 26962 10612 28476
rect 10556 26910 10558 26962
rect 10610 26910 10612 26962
rect 10556 25396 10612 26910
rect 10668 26290 10724 26302
rect 10668 26238 10670 26290
rect 10722 26238 10724 26290
rect 10668 25730 10724 26238
rect 10668 25678 10670 25730
rect 10722 25678 10724 25730
rect 10668 25666 10724 25678
rect 10556 25330 10612 25340
rect 10668 25508 10724 25518
rect 10556 24724 10612 24734
rect 10556 24630 10612 24668
rect 10500 22204 10612 22260
rect 10444 22194 10500 22204
rect 10444 21588 10500 21626
rect 10444 21522 10500 21532
rect 10444 21364 10500 21374
rect 10220 20850 10276 20860
rect 10332 21028 10388 21038
rect 10332 20914 10388 20972
rect 10332 20862 10334 20914
rect 10386 20862 10388 20914
rect 10332 20850 10388 20862
rect 10108 20636 10276 20692
rect 9996 20013 10052 20025
rect 10220 20020 10276 20636
rect 9996 19961 9998 20013
rect 10050 19961 10052 20013
rect 9996 19908 10052 19961
rect 9996 19842 10052 19852
rect 10108 19964 10276 20020
rect 9884 19506 9940 19516
rect 9884 19348 9940 19358
rect 9884 19254 9940 19292
rect 9884 18226 9940 18238
rect 9884 18174 9886 18226
rect 9938 18174 9940 18226
rect 9884 18004 9940 18174
rect 9884 17938 9940 17948
rect 9772 13746 9828 17276
rect 9996 17666 10052 17678
rect 9996 17614 9998 17666
rect 10050 17614 10052 17666
rect 9996 17444 10052 17614
rect 9996 17108 10052 17388
rect 9996 17042 10052 17052
rect 9884 16884 9940 16894
rect 9884 16790 9940 16828
rect 9996 16658 10052 16670
rect 9996 16606 9998 16658
rect 10050 16606 10052 16658
rect 9996 16098 10052 16606
rect 9996 16046 9998 16098
rect 10050 16046 10052 16098
rect 9996 16034 10052 16046
rect 9884 15988 9940 15998
rect 9884 15538 9940 15932
rect 9884 15486 9886 15538
rect 9938 15486 9940 15538
rect 9884 15474 9940 15486
rect 9772 13694 9774 13746
rect 9826 13694 9828 13746
rect 9772 12628 9828 13694
rect 9884 14530 9940 14542
rect 9884 14478 9886 14530
rect 9938 14478 9940 14530
rect 9884 13636 9940 14478
rect 10108 14084 10164 19964
rect 10220 19796 10276 19806
rect 10220 14418 10276 19740
rect 10332 19234 10388 19246
rect 10332 19182 10334 19234
rect 10386 19182 10388 19234
rect 10332 17444 10388 19182
rect 10444 18676 10500 21308
rect 10556 20018 10612 22204
rect 10556 19966 10558 20018
rect 10610 19966 10612 20018
rect 10556 19954 10612 19966
rect 10668 19236 10724 25452
rect 10780 22484 10836 31388
rect 10892 30772 10948 30782
rect 10892 30322 10948 30716
rect 10892 30270 10894 30322
rect 10946 30270 10948 30322
rect 10892 30258 10948 30270
rect 10892 29428 10948 29438
rect 10892 26292 10948 29372
rect 11004 29204 11060 34078
rect 11228 32788 11284 32798
rect 11116 31892 11172 31902
rect 11116 31798 11172 31836
rect 11228 31444 11284 32732
rect 11340 32116 11396 34300
rect 11788 34132 11844 34142
rect 11788 34038 11844 34076
rect 11452 32340 11508 32350
rect 11452 32338 11732 32340
rect 11452 32286 11454 32338
rect 11506 32286 11732 32338
rect 11452 32284 11732 32286
rect 11452 32274 11508 32284
rect 11340 32060 11620 32116
rect 11116 31388 11284 31444
rect 11340 31668 11396 31678
rect 11116 30100 11172 31388
rect 11228 31220 11284 31230
rect 11228 30882 11284 31164
rect 11228 30830 11230 30882
rect 11282 30830 11284 30882
rect 11228 30818 11284 30830
rect 11340 30994 11396 31612
rect 11340 30942 11342 30994
rect 11394 30942 11396 30994
rect 11340 30436 11396 30942
rect 11452 31666 11508 31678
rect 11452 31614 11454 31666
rect 11506 31614 11508 31666
rect 11452 30996 11508 31614
rect 11452 30930 11508 30940
rect 11564 30772 11620 32060
rect 11676 31780 11732 32284
rect 11788 31780 11844 31790
rect 11676 31778 11844 31780
rect 11676 31726 11790 31778
rect 11842 31726 11844 31778
rect 11676 31724 11844 31726
rect 11788 31714 11844 31724
rect 11788 30994 11844 31006
rect 11788 30942 11790 30994
rect 11842 30942 11844 30994
rect 11788 30884 11844 30942
rect 11340 30370 11396 30380
rect 11452 30716 11620 30772
rect 11676 30828 11844 30884
rect 11116 30044 11284 30100
rect 11004 29138 11060 29148
rect 11116 28644 11172 28654
rect 11116 28550 11172 28588
rect 11004 27748 11060 27758
rect 11004 27654 11060 27692
rect 10892 26226 10948 26236
rect 11116 26628 11172 26638
rect 11116 26290 11172 26572
rect 11116 26238 11118 26290
rect 11170 26238 11172 26290
rect 11116 26226 11172 26238
rect 11116 24836 11172 24846
rect 11228 24836 11284 30044
rect 11340 29988 11396 29998
rect 11340 28756 11396 29932
rect 11340 25506 11396 28700
rect 11340 25454 11342 25506
rect 11394 25454 11396 25506
rect 11340 25442 11396 25454
rect 11452 25620 11508 30716
rect 11676 30212 11732 30828
rect 11900 30772 11956 54236
rect 12572 52836 12628 52846
rect 12460 47012 12516 47022
rect 12460 43708 12516 46956
rect 12348 43652 12516 43708
rect 12124 41076 12180 41086
rect 12124 40982 12180 41020
rect 12236 40292 12292 40302
rect 12124 40180 12180 40190
rect 12124 40086 12180 40124
rect 12236 38946 12292 40236
rect 12236 38894 12238 38946
rect 12290 38894 12292 38946
rect 12236 38882 12292 38894
rect 12012 37380 12068 37390
rect 12012 37286 12068 37324
rect 12012 33124 12068 33134
rect 12012 33122 12180 33124
rect 12012 33070 12014 33122
rect 12066 33070 12180 33122
rect 12012 33068 12180 33070
rect 12012 33058 12068 33068
rect 11676 30146 11732 30156
rect 11788 30716 11956 30772
rect 12012 32900 12068 32910
rect 11564 29652 11620 29662
rect 11564 28868 11620 29596
rect 11564 28754 11620 28812
rect 11564 28702 11566 28754
rect 11618 28702 11620 28754
rect 11564 28690 11620 28702
rect 11676 29314 11732 29326
rect 11676 29262 11678 29314
rect 11730 29262 11732 29314
rect 11676 27972 11732 29262
rect 11676 27906 11732 27916
rect 11564 26964 11620 26974
rect 11564 26870 11620 26908
rect 11788 26908 11844 30716
rect 12012 30660 12068 32844
rect 12124 32116 12180 33068
rect 12124 32050 12180 32060
rect 12236 31778 12292 31790
rect 12236 31726 12238 31778
rect 12290 31726 12292 31778
rect 12236 31668 12292 31726
rect 12236 31602 12292 31612
rect 12348 31444 12404 43652
rect 12572 39844 12628 52780
rect 12796 43708 12852 55246
rect 14364 53844 14420 53854
rect 13692 45332 13748 45342
rect 12796 43652 12964 43708
rect 12796 40292 12852 40302
rect 12572 39778 12628 39788
rect 12684 40290 12852 40292
rect 12684 40238 12798 40290
rect 12850 40238 12852 40290
rect 12684 40236 12852 40238
rect 12572 38948 12628 38958
rect 12572 36596 12628 38892
rect 12572 36530 12628 36540
rect 12684 35140 12740 40236
rect 12796 40226 12852 40236
rect 12908 40068 12964 43652
rect 12908 40002 12964 40012
rect 13244 41412 13300 41422
rect 13132 38834 13188 38846
rect 13132 38782 13134 38834
rect 13186 38782 13188 38834
rect 12796 38724 12852 38734
rect 12796 38722 13076 38724
rect 12796 38670 12798 38722
rect 12850 38670 13076 38722
rect 12796 38668 13076 38670
rect 12796 38658 12852 38668
rect 12908 38612 13076 38668
rect 12684 35074 12740 35084
rect 12796 37268 12852 37278
rect 12684 34132 12740 34142
rect 12572 34130 12740 34132
rect 12572 34078 12686 34130
rect 12738 34078 12740 34130
rect 12572 34076 12740 34078
rect 12572 33346 12628 34076
rect 12684 34066 12740 34076
rect 12572 33294 12574 33346
rect 12626 33294 12628 33346
rect 12572 32676 12628 33294
rect 12684 33684 12740 33694
rect 12684 33012 12740 33628
rect 12684 32946 12740 32956
rect 12572 32610 12628 32620
rect 12796 32004 12852 37212
rect 12908 32900 12964 38612
rect 13132 38276 13188 38782
rect 13132 38210 13188 38220
rect 12908 32834 12964 32844
rect 13020 37380 13076 37390
rect 12796 31938 12852 31948
rect 12908 32116 12964 32126
rect 12460 31892 12516 31902
rect 12460 31798 12516 31836
rect 12908 31890 12964 32060
rect 12908 31838 12910 31890
rect 12962 31838 12964 31890
rect 12908 31826 12964 31838
rect 13020 31668 13076 37324
rect 13132 37266 13188 37278
rect 13132 37214 13134 37266
rect 13186 37214 13188 37266
rect 13132 33684 13188 37214
rect 13132 33618 13188 33628
rect 13244 33460 13300 41356
rect 13468 40628 13524 40638
rect 13356 40178 13412 40190
rect 13356 40126 13358 40178
rect 13410 40126 13412 40178
rect 13356 38724 13412 40126
rect 13356 38658 13412 38668
rect 11900 30604 12068 30660
rect 12124 31388 12404 31444
rect 12572 31612 13076 31668
rect 13132 33404 13300 33460
rect 13356 34132 13412 34142
rect 11900 29652 11956 30604
rect 12124 30436 12180 31388
rect 12236 31220 12292 31230
rect 12236 31106 12292 31164
rect 12236 31054 12238 31106
rect 12290 31054 12292 31106
rect 12236 31042 12292 31054
rect 11900 29586 11956 29596
rect 12012 30380 12180 30436
rect 11900 28644 11956 28654
rect 11900 28550 11956 28588
rect 12012 27860 12068 30380
rect 12236 30324 12292 30334
rect 12124 30212 12180 30222
rect 12124 30118 12180 30156
rect 12236 29428 12292 30268
rect 12572 30212 12628 31612
rect 12796 30436 12852 30446
rect 12572 30210 12740 30212
rect 12572 30158 12574 30210
rect 12626 30158 12740 30210
rect 12572 30156 12740 30158
rect 12572 30146 12628 30156
rect 12124 29372 12292 29428
rect 12124 28644 12180 29372
rect 12236 29204 12292 29214
rect 12236 29202 12628 29204
rect 12236 29150 12238 29202
rect 12290 29150 12628 29202
rect 12236 29148 12628 29150
rect 12236 29138 12292 29148
rect 12572 28866 12628 29148
rect 12572 28814 12574 28866
rect 12626 28814 12628 28866
rect 12572 28802 12628 28814
rect 12348 28644 12404 28654
rect 12124 28642 12404 28644
rect 12124 28590 12350 28642
rect 12402 28590 12404 28642
rect 12124 28588 12404 28590
rect 12124 28420 12180 28430
rect 12124 28082 12180 28364
rect 12124 28030 12126 28082
rect 12178 28030 12180 28082
rect 12124 28018 12180 28030
rect 12012 27804 12180 27860
rect 12012 27300 12068 27310
rect 12012 27206 12068 27244
rect 11788 26852 11956 26908
rect 11452 25508 11508 25564
rect 11676 26180 11732 26190
rect 11676 25618 11732 26124
rect 11676 25566 11678 25618
rect 11730 25566 11732 25618
rect 11676 25554 11732 25566
rect 11452 25452 11620 25508
rect 11564 25396 11620 25452
rect 11564 25340 11732 25396
rect 11116 24834 11284 24836
rect 11116 24782 11118 24834
rect 11170 24782 11284 24834
rect 11116 24780 11284 24782
rect 11452 25172 11508 25182
rect 11116 24770 11172 24780
rect 10892 23940 10948 23950
rect 10892 23938 11172 23940
rect 10892 23886 10894 23938
rect 10946 23886 11172 23938
rect 10892 23884 11172 23886
rect 10892 23874 10948 23884
rect 10892 22930 10948 22942
rect 10892 22878 10894 22930
rect 10946 22878 10948 22930
rect 10892 22596 10948 22878
rect 11116 22820 11172 23884
rect 11228 23828 11284 23838
rect 11228 23734 11284 23772
rect 11116 22764 11396 22820
rect 11228 22596 11284 22606
rect 10892 22540 11228 22596
rect 10780 22418 10836 22428
rect 11116 22148 11172 22158
rect 11004 22146 11172 22148
rect 11004 22094 11118 22146
rect 11170 22094 11172 22146
rect 11004 22092 11172 22094
rect 11004 21700 11060 22092
rect 11116 22082 11172 22092
rect 10780 21644 11060 21700
rect 10780 20802 10836 21644
rect 10780 20750 10782 20802
rect 10834 20750 10836 20802
rect 10780 20738 10836 20750
rect 10892 21476 10948 21486
rect 10892 20244 10948 21420
rect 11004 21364 11060 21374
rect 11004 21270 11060 21308
rect 11116 21252 11172 21262
rect 11116 20802 11172 21196
rect 11116 20750 11118 20802
rect 11170 20750 11172 20802
rect 11116 20738 11172 20750
rect 11228 20804 11284 22540
rect 11340 21026 11396 22764
rect 11452 21700 11508 25116
rect 11564 23938 11620 23950
rect 11564 23886 11566 23938
rect 11618 23886 11620 23938
rect 11564 21924 11620 23886
rect 11676 22708 11732 25340
rect 11676 22642 11732 22652
rect 11788 23604 11844 23614
rect 11788 22484 11844 23548
rect 11676 22428 11844 22484
rect 11676 22036 11732 22428
rect 11788 22260 11844 22270
rect 11788 22166 11844 22204
rect 11676 21980 11844 22036
rect 11564 21858 11620 21868
rect 11452 21644 11620 21700
rect 11340 20974 11342 21026
rect 11394 20974 11396 21026
rect 11340 20962 11396 20974
rect 11228 20748 11396 20804
rect 11228 20468 11284 20478
rect 11116 20244 11172 20254
rect 10892 20188 11116 20244
rect 10892 19908 10948 19918
rect 10892 19458 10948 19852
rect 11004 19684 11060 20188
rect 11116 20150 11172 20188
rect 11004 19618 11060 19628
rect 10892 19406 10894 19458
rect 10946 19406 10948 19458
rect 10892 19394 10948 19406
rect 10668 19180 10948 19236
rect 10444 18564 10500 18620
rect 10780 18676 10836 18686
rect 10556 18564 10612 18574
rect 10444 18562 10612 18564
rect 10444 18510 10558 18562
rect 10610 18510 10612 18562
rect 10444 18508 10612 18510
rect 10556 18498 10612 18508
rect 10332 17378 10388 17388
rect 10444 18340 10500 18350
rect 10444 17890 10500 18284
rect 10444 17838 10446 17890
rect 10498 17838 10500 17890
rect 10444 17108 10500 17838
rect 10332 17052 10500 17108
rect 10332 15148 10388 17052
rect 10556 16882 10612 16894
rect 10556 16830 10558 16882
rect 10610 16830 10612 16882
rect 10444 16212 10500 16222
rect 10444 16118 10500 16156
rect 10556 15988 10612 16830
rect 10556 15922 10612 15932
rect 10556 15540 10612 15550
rect 10556 15426 10612 15484
rect 10556 15374 10558 15426
rect 10610 15374 10612 15426
rect 10556 15362 10612 15374
rect 10332 15092 10612 15148
rect 10220 14366 10222 14418
rect 10274 14366 10276 14418
rect 10220 14354 10276 14366
rect 10108 14028 10388 14084
rect 9996 13636 10052 13646
rect 9884 13634 10052 13636
rect 9884 13582 9998 13634
rect 10050 13582 10052 13634
rect 9884 13580 10052 13582
rect 9996 13570 10052 13580
rect 10220 13636 10276 13646
rect 9996 12852 10052 12862
rect 9996 12758 10052 12796
rect 9772 12572 10052 12628
rect 9660 12516 9716 12526
rect 9660 12068 9716 12460
rect 9772 12068 9828 12078
rect 9660 12066 9828 12068
rect 9660 12014 9774 12066
rect 9826 12014 9828 12066
rect 9660 12012 9828 12014
rect 9772 12002 9828 12012
rect 9772 11844 9828 11854
rect 9772 11618 9828 11788
rect 9772 11566 9774 11618
rect 9826 11566 9828 11618
rect 9772 11554 9828 11566
rect 9884 11508 9940 11518
rect 9884 11414 9940 11452
rect 9548 10668 9828 10724
rect 9436 10546 9492 10556
rect 9324 10498 9380 10510
rect 9324 10446 9326 10498
rect 9378 10446 9380 10498
rect 9324 9044 9380 10446
rect 9660 10500 9716 10510
rect 9660 10406 9716 10444
rect 9548 10388 9604 10398
rect 9548 10294 9604 10332
rect 9548 9826 9604 9838
rect 9548 9774 9550 9826
rect 9602 9774 9604 9826
rect 9548 9268 9604 9774
rect 9660 9268 9716 9278
rect 9548 9266 9716 9268
rect 9548 9214 9662 9266
rect 9714 9214 9716 9266
rect 9548 9212 9716 9214
rect 9660 9202 9716 9212
rect 9324 8978 9380 8988
rect 9660 8596 9716 8606
rect 9324 8484 9380 8494
rect 9324 7586 9380 8428
rect 9324 7534 9326 7586
rect 9378 7534 9380 7586
rect 9324 7522 9380 7534
rect 9660 6690 9716 8540
rect 9772 8372 9828 10668
rect 9884 10386 9940 10398
rect 9884 10334 9886 10386
rect 9938 10334 9940 10386
rect 9884 9156 9940 10334
rect 9996 9826 10052 12572
rect 10108 10498 10164 10510
rect 10108 10446 10110 10498
rect 10162 10446 10164 10498
rect 10108 10164 10164 10446
rect 10108 10098 10164 10108
rect 9996 9774 9998 9826
rect 10050 9774 10052 9826
rect 9996 9762 10052 9774
rect 10108 9938 10164 9950
rect 10108 9886 10110 9938
rect 10162 9886 10164 9938
rect 9884 9090 9940 9100
rect 9996 9604 10052 9614
rect 9996 8484 10052 9548
rect 9996 8418 10052 8428
rect 9772 8306 9828 8316
rect 9772 7364 9828 7374
rect 9772 7270 9828 7308
rect 9660 6638 9662 6690
rect 9714 6638 9716 6690
rect 9660 6626 9716 6638
rect 10108 6690 10164 9886
rect 10220 8372 10276 13580
rect 10332 13074 10388 14028
rect 10332 13022 10334 13074
rect 10386 13022 10388 13074
rect 10332 13010 10388 13022
rect 10444 13524 10500 13534
rect 10332 12516 10388 12526
rect 10332 9604 10388 12460
rect 10332 9538 10388 9548
rect 10444 9268 10500 13468
rect 10220 8306 10276 8316
rect 10332 9212 10500 9268
rect 10108 6638 10110 6690
rect 10162 6638 10164 6690
rect 10108 6626 10164 6638
rect 9324 6020 9380 6030
rect 9212 6018 9380 6020
rect 9212 5966 9326 6018
rect 9378 5966 9380 6018
rect 9212 5964 9380 5966
rect 9324 5954 9380 5964
rect 8876 5682 8932 5694
rect 8876 5630 8878 5682
rect 8930 5630 8932 5682
rect 8316 5460 8372 5470
rect 7756 5348 7812 5358
rect 7756 5254 7812 5292
rect 8316 5234 8372 5404
rect 8876 5348 8932 5630
rect 8876 5282 8932 5292
rect 8316 5182 8318 5234
rect 8370 5182 8372 5234
rect 8316 5170 8372 5182
rect 6524 4946 6580 4956
rect 6636 5124 6692 5134
rect 6636 4452 6692 5068
rect 8764 5124 8820 5134
rect 6636 4386 6692 4396
rect 7980 5012 8036 5022
rect 6300 3332 6468 3388
rect 6412 3220 6468 3332
rect 3804 3164 4068 3174
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 3804 3098 4068 3108
rect 6076 3164 6468 3220
rect 4464 2380 4728 2390
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4464 2314 4728 2324
rect 3388 1652 3444 1662
rect 3388 112 3444 1596
rect 3804 1596 4068 1606
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 3804 1530 4068 1540
rect 4464 812 4728 822
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4464 746 4728 756
rect 4732 420 4788 430
rect 4732 112 4788 364
rect 6076 112 6132 3164
rect 7980 1314 8036 4956
rect 7980 1262 7982 1314
rect 8034 1262 8036 1314
rect 7980 1250 8036 1262
rect 7532 980 7588 990
rect 7420 978 7588 980
rect 7420 926 7534 978
rect 7586 926 7588 978
rect 7420 924 7588 926
rect 7420 112 7476 924
rect 7532 914 7588 924
rect 8764 112 8820 5068
rect 10332 2100 10388 9212
rect 10444 9044 10500 9054
rect 10444 8260 10500 8988
rect 10556 8484 10612 15092
rect 10780 14530 10836 18620
rect 10892 18004 10948 19180
rect 11004 18228 11060 18238
rect 11004 18226 11172 18228
rect 11004 18174 11006 18226
rect 11058 18174 11172 18226
rect 11004 18172 11172 18174
rect 11004 18162 11060 18172
rect 11116 18004 11172 18172
rect 10892 17948 11060 18004
rect 10892 15204 10948 15242
rect 10892 15138 10948 15148
rect 10780 14478 10782 14530
rect 10834 14478 10836 14530
rect 10668 13746 10724 13758
rect 10668 13694 10670 13746
rect 10722 13694 10724 13746
rect 10668 12292 10724 13694
rect 10780 12516 10836 14478
rect 11004 13746 11060 17948
rect 11116 17938 11172 17948
rect 11116 17444 11172 17454
rect 11116 17108 11172 17388
rect 11116 16098 11172 17052
rect 11228 16882 11284 20412
rect 11228 16830 11230 16882
rect 11282 16830 11284 16882
rect 11228 16818 11284 16830
rect 11340 16660 11396 20748
rect 11116 16046 11118 16098
rect 11170 16046 11172 16098
rect 11116 16034 11172 16046
rect 11228 16604 11396 16660
rect 11452 18004 11508 18014
rect 11564 18004 11620 21644
rect 11508 17948 11620 18004
rect 11676 18228 11732 18238
rect 11228 15148 11284 16604
rect 11004 13694 11006 13746
rect 11058 13694 11060 13746
rect 11004 13682 11060 13694
rect 11116 15092 11284 15148
rect 10780 12450 10836 12460
rect 11004 12292 11060 12302
rect 10668 12290 11060 12292
rect 10668 12238 11006 12290
rect 11058 12238 11060 12290
rect 10668 12236 11060 12238
rect 11004 12226 11060 12236
rect 11116 11956 11172 15092
rect 11340 14642 11396 14654
rect 11340 14590 11342 14642
rect 11394 14590 11396 14642
rect 10668 11900 11172 11956
rect 11228 13746 11284 13758
rect 11228 13694 11230 13746
rect 11282 13694 11284 13746
rect 10668 10724 10724 11900
rect 11116 11732 11172 11742
rect 11004 11506 11060 11518
rect 11004 11454 11006 11506
rect 11058 11454 11060 11506
rect 10668 10658 10724 10668
rect 10780 11394 10836 11406
rect 10780 11342 10782 11394
rect 10834 11342 10836 11394
rect 10668 10500 10724 10510
rect 10780 10500 10836 11342
rect 10892 10948 10948 10958
rect 10892 10610 10948 10892
rect 10892 10558 10894 10610
rect 10946 10558 10948 10610
rect 10892 10546 10948 10558
rect 10668 10498 10836 10500
rect 10668 10446 10670 10498
rect 10722 10446 10836 10498
rect 10668 10444 10836 10446
rect 10668 10434 10724 10444
rect 10892 10388 10948 10398
rect 10780 9826 10836 9838
rect 10780 9774 10782 9826
rect 10834 9774 10836 9826
rect 10556 8428 10724 8484
rect 10556 8260 10612 8270
rect 10444 8258 10612 8260
rect 10444 8206 10558 8258
rect 10610 8206 10612 8258
rect 10444 8204 10612 8206
rect 10556 8194 10612 8204
rect 10668 7364 10724 8428
rect 10780 7700 10836 9774
rect 10892 8930 10948 10332
rect 11004 9044 11060 11454
rect 11116 11506 11172 11676
rect 11116 11454 11118 11506
rect 11170 11454 11172 11506
rect 11116 11442 11172 11454
rect 11116 11060 11172 11070
rect 11116 10724 11172 11004
rect 11228 10724 11284 13694
rect 11340 13636 11396 14590
rect 11340 13570 11396 13580
rect 11452 13076 11508 17948
rect 11564 17444 11620 17454
rect 11564 17350 11620 17388
rect 11676 16322 11732 18172
rect 11676 16270 11678 16322
rect 11730 16270 11732 16322
rect 11676 13412 11732 16270
rect 11676 13346 11732 13356
rect 11676 13076 11732 13086
rect 11452 13020 11676 13076
rect 11564 12740 11620 12750
rect 11340 12738 11620 12740
rect 11340 12686 11566 12738
rect 11618 12686 11620 12738
rect 11340 12684 11620 12686
rect 11340 11060 11396 12684
rect 11564 12674 11620 12684
rect 11564 12180 11620 12190
rect 11676 12180 11732 13020
rect 11564 12178 11732 12180
rect 11564 12126 11566 12178
rect 11618 12126 11732 12178
rect 11564 12124 11732 12126
rect 11564 12114 11620 12124
rect 11340 10994 11396 11004
rect 11452 11732 11508 11742
rect 11452 11618 11508 11676
rect 11452 11566 11454 11618
rect 11506 11566 11508 11618
rect 11228 10668 11396 10724
rect 11116 10498 11172 10668
rect 11116 10446 11118 10498
rect 11170 10446 11172 10498
rect 11116 10434 11172 10446
rect 11228 10388 11284 10398
rect 11228 10294 11284 10332
rect 11340 9826 11396 10668
rect 11452 10610 11508 11566
rect 11676 11396 11732 11434
rect 11676 11330 11732 11340
rect 11564 11282 11620 11294
rect 11564 11230 11566 11282
rect 11618 11230 11620 11282
rect 11564 10948 11620 11230
rect 11564 10882 11620 10892
rect 11676 11172 11732 11182
rect 11676 10724 11732 11116
rect 11788 11060 11844 21980
rect 11788 10994 11844 11004
rect 11900 10836 11956 26852
rect 12012 26852 12068 26862
rect 12012 26290 12068 26796
rect 12012 26238 12014 26290
rect 12066 26238 12068 26290
rect 12012 26226 12068 26238
rect 12012 25060 12068 25070
rect 12012 23938 12068 25004
rect 12012 23886 12014 23938
rect 12066 23886 12068 23938
rect 12012 23874 12068 23886
rect 12012 22930 12068 22942
rect 12012 22878 12014 22930
rect 12066 22878 12068 22930
rect 12012 20802 12068 22878
rect 12124 21924 12180 27804
rect 12348 26908 12404 28588
rect 12684 28308 12740 30156
rect 12684 28242 12740 28252
rect 12796 26908 12852 30380
rect 12908 30210 12964 30222
rect 12908 30158 12910 30210
rect 12962 30158 12964 30210
rect 12908 30100 12964 30158
rect 12908 30034 12964 30044
rect 13020 28642 13076 28654
rect 13020 28590 13022 28642
rect 13074 28590 13076 28642
rect 13020 28420 13076 28590
rect 13020 28354 13076 28364
rect 13132 27524 13188 33404
rect 13244 33234 13300 33246
rect 13244 33182 13246 33234
rect 13298 33182 13300 33234
rect 13244 32564 13300 33182
rect 13244 32498 13300 32508
rect 13356 32340 13412 34076
rect 13244 32284 13412 32340
rect 13244 29988 13300 32284
rect 13468 32116 13524 40572
rect 13580 38836 13636 38846
rect 13580 38742 13636 38780
rect 13580 38500 13636 38510
rect 13580 37156 13636 38444
rect 13580 37062 13636 37100
rect 13580 36370 13636 36382
rect 13580 36318 13582 36370
rect 13634 36318 13636 36370
rect 13580 35698 13636 36318
rect 13580 35646 13582 35698
rect 13634 35646 13636 35698
rect 13580 35634 13636 35646
rect 13468 32050 13524 32060
rect 13580 34018 13636 34030
rect 13580 33966 13582 34018
rect 13634 33966 13636 34018
rect 13356 32004 13412 32014
rect 13356 30324 13412 31948
rect 13468 31778 13524 31790
rect 13468 31726 13470 31778
rect 13522 31726 13524 31778
rect 13468 31332 13524 31726
rect 13580 31668 13636 33966
rect 13580 31602 13636 31612
rect 13468 31266 13524 31276
rect 13468 30996 13524 31006
rect 13468 30994 13636 30996
rect 13468 30942 13470 30994
rect 13522 30942 13636 30994
rect 13468 30940 13636 30942
rect 13468 30930 13524 30940
rect 13580 30884 13636 30940
rect 13580 30818 13636 30828
rect 13356 30210 13412 30268
rect 13356 30158 13358 30210
rect 13410 30158 13412 30210
rect 13356 30146 13412 30158
rect 13580 30322 13636 30334
rect 13580 30270 13582 30322
rect 13634 30270 13636 30322
rect 13244 29932 13412 29988
rect 13132 27468 13300 27524
rect 12908 27300 12964 27310
rect 13132 27300 13188 27310
rect 12964 27244 13076 27300
rect 12908 27234 12964 27244
rect 12348 26852 12516 26908
rect 12796 26852 12964 26908
rect 12460 26404 12516 26852
rect 12460 26338 12516 26348
rect 12684 25732 12740 25742
rect 12236 24164 12292 24174
rect 12236 24070 12292 24108
rect 12572 23940 12628 23950
rect 12236 22596 12292 22606
rect 12236 22502 12292 22540
rect 12124 21858 12180 21868
rect 12124 21588 12180 21598
rect 12124 21494 12180 21532
rect 12012 20750 12014 20802
rect 12066 20750 12068 20802
rect 12012 20738 12068 20750
rect 12348 21140 12404 21150
rect 12348 20804 12404 21084
rect 12348 20802 12516 20804
rect 12348 20750 12350 20802
rect 12402 20750 12516 20802
rect 12348 20748 12516 20750
rect 12348 20738 12404 20748
rect 12460 20468 12516 20748
rect 12460 20402 12516 20412
rect 12572 19572 12628 23884
rect 12684 19684 12740 25676
rect 12908 25508 12964 26852
rect 12908 25442 12964 25452
rect 12908 25282 12964 25294
rect 12908 25230 12910 25282
rect 12962 25230 12964 25282
rect 12796 24498 12852 24510
rect 12796 24446 12798 24498
rect 12850 24446 12852 24498
rect 12796 24164 12852 24446
rect 12796 24098 12852 24108
rect 12908 23938 12964 25230
rect 12908 23886 12910 23938
rect 12962 23886 12964 23938
rect 12908 23874 12964 23886
rect 13020 23548 13076 27244
rect 13132 27206 13188 27244
rect 13244 26908 13300 27468
rect 13132 26852 13300 26908
rect 13132 25732 13188 26852
rect 13356 26740 13412 29932
rect 13580 29426 13636 30270
rect 13580 29374 13582 29426
rect 13634 29374 13636 29426
rect 13580 29362 13636 29374
rect 13580 28644 13636 28654
rect 13580 28550 13636 28588
rect 13580 28308 13636 28318
rect 13580 27970 13636 28252
rect 13580 27918 13582 27970
rect 13634 27918 13636 27970
rect 13580 27748 13636 27918
rect 13580 27682 13636 27692
rect 13356 26684 13524 26740
rect 13356 26516 13412 26526
rect 13132 25666 13188 25676
rect 13244 26290 13300 26302
rect 13244 26238 13246 26290
rect 13298 26238 13300 26290
rect 13244 25844 13300 26238
rect 12908 23492 13076 23548
rect 13132 25508 13188 25518
rect 12684 19618 12740 19628
rect 12796 20020 12852 20030
rect 12796 19906 12852 19964
rect 12796 19854 12798 19906
rect 12850 19854 12852 19906
rect 12572 19506 12628 19516
rect 12796 19460 12852 19854
rect 12796 19394 12852 19404
rect 12012 19348 12068 19358
rect 12012 19346 12628 19348
rect 12012 19294 12014 19346
rect 12066 19294 12628 19346
rect 12012 19292 12628 19294
rect 12012 19282 12068 19292
rect 12572 19236 12628 19292
rect 12796 19236 12852 19246
rect 12572 19234 12852 19236
rect 12572 19182 12798 19234
rect 12850 19182 12852 19234
rect 12572 19180 12852 19182
rect 12796 19170 12852 19180
rect 12012 19124 12068 19134
rect 12012 16882 12068 19068
rect 12460 19124 12516 19134
rect 12460 19030 12516 19068
rect 12908 18900 12964 23492
rect 13132 20356 13188 25452
rect 13244 25396 13300 25788
rect 13244 25330 13300 25340
rect 13356 24836 13412 26460
rect 13244 24780 13412 24836
rect 13244 23266 13300 24780
rect 13244 23214 13246 23266
rect 13298 23214 13300 23266
rect 13244 23202 13300 23214
rect 13356 24610 13412 24622
rect 13356 24558 13358 24610
rect 13410 24558 13412 24610
rect 13356 22820 13412 24558
rect 13468 23940 13524 26684
rect 13692 26178 13748 45276
rect 14140 41970 14196 41982
rect 14140 41918 14142 41970
rect 14194 41918 14196 41970
rect 13916 41076 13972 41086
rect 13916 40982 13972 41020
rect 14028 39618 14084 39630
rect 14028 39566 14030 39618
rect 14082 39566 14084 39618
rect 13916 38836 13972 38846
rect 13804 38724 13860 38734
rect 13804 38630 13860 38668
rect 13804 37044 13860 37054
rect 13804 32564 13860 36988
rect 13804 32498 13860 32508
rect 13916 31220 13972 38780
rect 14028 35026 14084 39566
rect 14140 39284 14196 41918
rect 14364 41524 14420 53788
rect 14700 41972 14756 55804
rect 14700 41906 14756 41916
rect 14364 41458 14420 41468
rect 14588 41858 14644 41870
rect 14588 41806 14590 41858
rect 14642 41806 14644 41858
rect 14364 41300 14420 41310
rect 14588 41300 14644 41806
rect 15596 41748 15652 55918
rect 16940 55468 16996 57148
rect 18172 56308 18228 57344
rect 19516 57316 19572 57344
rect 19516 57250 19572 57260
rect 19852 57316 19908 57372
rect 19852 57250 19908 57260
rect 18508 56308 18564 56318
rect 18172 56306 18564 56308
rect 18172 56254 18510 56306
rect 18562 56254 18564 56306
rect 18172 56252 18564 56254
rect 18508 56242 18564 56252
rect 20300 56306 20356 57372
rect 20832 57344 20944 57456
rect 22176 57344 22288 57456
rect 22540 57372 23044 57428
rect 20300 56254 20302 56306
rect 20354 56254 20356 56306
rect 20300 56242 20356 56254
rect 20860 56308 20916 57344
rect 22204 57204 22260 57344
rect 22540 57204 22596 57372
rect 22204 57148 22596 57204
rect 20860 56242 20916 56252
rect 22204 56308 22260 56318
rect 22204 56214 22260 56252
rect 22540 56196 22596 56206
rect 21756 56082 21812 56094
rect 21756 56030 21758 56082
rect 21810 56030 21812 56082
rect 17500 55970 17556 55982
rect 17500 55918 17502 55970
rect 17554 55918 17556 55970
rect 16940 55412 17332 55468
rect 17276 55186 17332 55412
rect 17276 55134 17278 55186
rect 17330 55134 17332 55186
rect 17276 55122 17332 55134
rect 16828 53732 16884 53742
rect 16044 50484 16100 50494
rect 15596 41682 15652 41692
rect 15708 45892 15764 45902
rect 14364 41298 14644 41300
rect 14364 41246 14366 41298
rect 14418 41246 14644 41298
rect 14364 41244 14644 41246
rect 15036 41412 15092 41422
rect 14364 41234 14420 41244
rect 14364 41076 14420 41086
rect 14364 40402 14420 41020
rect 14364 40350 14366 40402
rect 14418 40350 14420 40402
rect 14364 40338 14420 40350
rect 14140 39218 14196 39228
rect 14252 40180 14308 40190
rect 14252 38834 14308 40124
rect 14476 39508 14532 41244
rect 14476 39442 14532 39452
rect 14588 40404 14644 40414
rect 14252 38782 14254 38834
rect 14306 38782 14308 38834
rect 14252 38770 14308 38782
rect 14028 34974 14030 35026
rect 14082 34974 14084 35026
rect 14028 34962 14084 34974
rect 14140 32116 14196 32126
rect 13972 31164 14084 31220
rect 13916 31154 13972 31164
rect 13916 30770 13972 30782
rect 13916 30718 13918 30770
rect 13970 30718 13972 30770
rect 13916 30660 13972 30718
rect 13916 30594 13972 30604
rect 14028 30436 14084 31164
rect 13916 30380 14084 30436
rect 13916 28980 13972 30380
rect 14028 30212 14084 30222
rect 14028 30118 14084 30156
rect 14028 29540 14084 29550
rect 14140 29540 14196 32060
rect 14476 31780 14532 31790
rect 14476 31686 14532 31724
rect 14364 30884 14420 30894
rect 14028 29538 14196 29540
rect 14028 29486 14030 29538
rect 14082 29486 14196 29538
rect 14028 29484 14196 29486
rect 14252 30212 14308 30222
rect 14028 29474 14084 29484
rect 13804 28756 13860 28766
rect 13804 27074 13860 28700
rect 13916 28644 13972 28924
rect 13916 28578 13972 28588
rect 13916 27858 13972 27870
rect 13916 27806 13918 27858
rect 13970 27806 13972 27858
rect 13916 27300 13972 27806
rect 14252 27860 14308 30156
rect 14364 29876 14420 30828
rect 14588 30772 14644 40348
rect 14924 40178 14980 40190
rect 14924 40126 14926 40178
rect 14978 40126 14980 40178
rect 14812 38836 14868 38846
rect 14812 38742 14868 38780
rect 14924 38500 14980 40126
rect 14924 38434 14980 38444
rect 14700 38052 14756 38062
rect 14700 38050 14868 38052
rect 14700 37998 14702 38050
rect 14754 37998 14868 38050
rect 14700 37996 14868 37998
rect 14700 37986 14756 37996
rect 14588 30706 14644 30716
rect 14700 37042 14756 37054
rect 14700 36990 14702 37042
rect 14754 36990 14756 37042
rect 14588 30212 14644 30222
rect 14364 29810 14420 29820
rect 14476 30210 14644 30212
rect 14476 30158 14590 30210
rect 14642 30158 14644 30210
rect 14476 30156 14644 30158
rect 14364 29316 14420 29326
rect 14476 29316 14532 30156
rect 14588 30146 14644 30156
rect 14700 29426 14756 36990
rect 14812 35586 14868 37996
rect 14812 35534 14814 35586
rect 14866 35534 14868 35586
rect 14812 32562 14868 35534
rect 14812 32510 14814 32562
rect 14866 32510 14868 32562
rect 14812 32498 14868 32510
rect 14700 29374 14702 29426
rect 14754 29374 14756 29426
rect 14700 29362 14756 29374
rect 14924 32228 14980 32238
rect 14364 29314 14532 29316
rect 14364 29262 14366 29314
rect 14418 29262 14532 29314
rect 14364 29260 14532 29262
rect 14364 29250 14420 29260
rect 14364 27860 14420 27870
rect 14252 27858 14420 27860
rect 14252 27806 14366 27858
rect 14418 27806 14420 27858
rect 14252 27804 14420 27806
rect 13916 27234 13972 27244
rect 14140 27188 14196 27198
rect 14140 27094 14196 27132
rect 13804 27022 13806 27074
rect 13858 27022 13860 27074
rect 13804 27010 13860 27022
rect 13916 27076 13972 27086
rect 13692 26126 13694 26178
rect 13746 26126 13748 26178
rect 13692 25172 13748 26126
rect 13692 25106 13748 25116
rect 13804 25956 13860 25966
rect 13692 24948 13748 24958
rect 13468 23846 13524 23884
rect 13580 24724 13636 24734
rect 13356 22754 13412 22764
rect 13468 23380 13524 23390
rect 13356 22596 13412 22606
rect 13356 22502 13412 22540
rect 13468 22372 13524 23324
rect 13468 22306 13524 22316
rect 13356 22036 13412 22046
rect 13356 20802 13412 21980
rect 13356 20750 13358 20802
rect 13410 20750 13412 20802
rect 13356 20738 13412 20750
rect 13468 21362 13524 21374
rect 13468 21310 13470 21362
rect 13522 21310 13524 21362
rect 13132 20290 13188 20300
rect 13132 20020 13188 20030
rect 13132 19926 13188 19964
rect 13468 19458 13524 21310
rect 13468 19406 13470 19458
rect 13522 19406 13524 19458
rect 13468 19394 13524 19406
rect 13580 20018 13636 24668
rect 13692 23380 13748 24892
rect 13804 23716 13860 25900
rect 13804 23650 13860 23660
rect 13692 23314 13748 23324
rect 13916 23156 13972 27020
rect 14252 26964 14308 26974
rect 13580 19966 13582 20018
rect 13634 19966 13636 20018
rect 13244 19236 13300 19246
rect 13244 19142 13300 19180
rect 13580 19236 13636 19966
rect 13692 23100 13972 23156
rect 14028 26740 14084 26750
rect 13692 19908 13748 23100
rect 13692 19842 13748 19852
rect 13804 22930 13860 22942
rect 13804 22878 13806 22930
rect 13858 22878 13860 22930
rect 13804 19906 13860 22878
rect 14028 21698 14084 26684
rect 14252 25956 14308 26908
rect 14252 25890 14308 25900
rect 14364 25732 14420 27804
rect 14140 25676 14420 25732
rect 14140 24724 14196 25676
rect 14476 25620 14532 29260
rect 14700 28642 14756 28654
rect 14700 28590 14702 28642
rect 14754 28590 14756 28642
rect 14588 27634 14644 27646
rect 14588 27582 14590 27634
rect 14642 27582 14644 27634
rect 14588 26292 14644 27582
rect 14700 26964 14756 28590
rect 14700 26898 14756 26908
rect 14924 26908 14980 32172
rect 15036 32116 15092 41356
rect 15484 40962 15540 40974
rect 15484 40910 15486 40962
rect 15538 40910 15540 40962
rect 15260 38836 15316 38846
rect 15148 38612 15204 38622
rect 15148 38274 15204 38556
rect 15148 38222 15150 38274
rect 15202 38222 15204 38274
rect 15148 38210 15204 38222
rect 15036 32050 15092 32060
rect 15148 37154 15204 37166
rect 15148 37102 15150 37154
rect 15202 37102 15204 37154
rect 15148 32004 15204 37102
rect 15148 31938 15204 31948
rect 15036 30884 15092 30894
rect 15036 30790 15092 30828
rect 15148 29428 15204 29438
rect 15148 29334 15204 29372
rect 15260 29204 15316 38780
rect 15484 37266 15540 40910
rect 15484 37214 15486 37266
rect 15538 37214 15540 37266
rect 15484 37202 15540 37214
rect 15596 39172 15652 39182
rect 15596 34804 15652 39116
rect 15708 38162 15764 45836
rect 15820 41748 15876 41758
rect 15820 41746 15988 41748
rect 15820 41694 15822 41746
rect 15874 41694 15988 41746
rect 15820 41692 15988 41694
rect 15820 41682 15876 41692
rect 15820 38836 15876 38846
rect 15820 38742 15876 38780
rect 15932 38668 15988 41692
rect 16044 40516 16100 50428
rect 16828 47012 16884 53676
rect 16828 46946 16884 46956
rect 17276 53620 17332 53630
rect 16940 46116 16996 46126
rect 16044 40450 16100 40460
rect 16716 41860 16772 41870
rect 16044 40180 16100 40190
rect 16044 40178 16660 40180
rect 16044 40126 16046 40178
rect 16098 40126 16660 40178
rect 16044 40124 16660 40126
rect 16044 40114 16100 40124
rect 15932 38612 16100 38668
rect 15708 38110 15710 38162
rect 15762 38110 15764 38162
rect 15708 38098 15764 38110
rect 15932 37268 15988 37278
rect 15932 37174 15988 37212
rect 15596 33234 15652 34748
rect 15596 33182 15598 33234
rect 15650 33182 15652 33234
rect 15596 33170 15652 33182
rect 15596 32676 15652 32686
rect 15596 32582 15652 32620
rect 15820 32340 15876 32350
rect 15708 30996 15764 31006
rect 15484 30882 15540 30894
rect 15484 30830 15486 30882
rect 15538 30830 15540 30882
rect 15484 29652 15540 30830
rect 15708 30436 15764 30940
rect 15820 30994 15876 32284
rect 15820 30942 15822 30994
rect 15874 30942 15876 30994
rect 15820 30930 15876 30942
rect 15932 32004 15988 32014
rect 15708 30380 15876 30436
rect 15484 29586 15540 29596
rect 15708 30210 15764 30222
rect 15708 30158 15710 30210
rect 15762 30158 15764 30210
rect 15484 29428 15540 29438
rect 15708 29428 15764 30158
rect 15540 29372 15652 29428
rect 15484 29362 15540 29372
rect 15148 29148 15316 29204
rect 15372 29204 15428 29214
rect 15372 29202 15540 29204
rect 15372 29150 15374 29202
rect 15426 29150 15540 29202
rect 15372 29148 15540 29150
rect 14924 26852 15092 26908
rect 14588 26226 14644 26236
rect 14364 25564 14532 25620
rect 14588 26068 14644 26078
rect 14364 24724 14420 25564
rect 14476 25396 14532 25406
rect 14588 25396 14644 26012
rect 14532 25340 14644 25396
rect 14812 26066 14868 26078
rect 14812 26014 14814 26066
rect 14866 26014 14868 26066
rect 14476 25302 14532 25340
rect 14812 24724 14868 26014
rect 14924 25732 14980 25742
rect 14924 25638 14980 25676
rect 14924 24724 14980 24734
rect 14364 24668 14532 24724
rect 14812 24722 14980 24724
rect 14812 24670 14926 24722
rect 14978 24670 14980 24722
rect 14812 24668 14980 24670
rect 14140 24658 14196 24668
rect 14364 24500 14420 24510
rect 14364 23938 14420 24444
rect 14364 23886 14366 23938
rect 14418 23886 14420 23938
rect 14364 23874 14420 23886
rect 14028 21646 14030 21698
rect 14082 21646 14084 21698
rect 14028 21634 14084 21646
rect 14364 22370 14420 22382
rect 14364 22318 14366 22370
rect 14418 22318 14420 22370
rect 14364 20804 14420 22318
rect 14476 21698 14532 24668
rect 14924 24658 14980 24668
rect 14476 21646 14478 21698
rect 14530 21646 14532 21698
rect 14476 21476 14532 21646
rect 14476 21410 14532 21420
rect 14588 24610 14644 24622
rect 14588 24558 14590 24610
rect 14642 24558 14644 24610
rect 14364 20710 14420 20748
rect 14588 20188 14644 24558
rect 13804 19854 13806 19906
rect 13858 19854 13860 19906
rect 13804 19842 13860 19854
rect 13916 20132 14644 20188
rect 14700 23156 14756 23166
rect 14700 20244 14756 23100
rect 14812 22484 14868 22494
rect 14812 22390 14868 22428
rect 14812 21588 14868 21598
rect 14812 21494 14868 21532
rect 14924 21028 14980 21038
rect 15036 21028 15092 26852
rect 15148 23716 15204 29148
rect 15372 29138 15428 29148
rect 15484 28866 15540 29148
rect 15484 28814 15486 28866
rect 15538 28814 15540 28866
rect 15484 28802 15540 28814
rect 15596 28196 15652 29372
rect 15708 29362 15764 29372
rect 15484 28140 15652 28196
rect 15708 28868 15764 28878
rect 15260 27858 15316 27870
rect 15260 27806 15262 27858
rect 15314 27806 15316 27858
rect 15260 27300 15316 27806
rect 15372 27300 15428 27310
rect 15260 27298 15428 27300
rect 15260 27246 15374 27298
rect 15426 27246 15428 27298
rect 15260 27244 15428 27246
rect 15372 27234 15428 27244
rect 15260 26292 15316 26302
rect 15260 26198 15316 26236
rect 15372 24724 15428 24734
rect 15372 24630 15428 24668
rect 15148 23650 15204 23660
rect 15260 24388 15316 24398
rect 15484 24388 15540 28140
rect 15596 26964 15652 26974
rect 15596 25172 15652 26908
rect 15596 25106 15652 25116
rect 15708 24948 15764 28812
rect 15820 27858 15876 30380
rect 15820 27806 15822 27858
rect 15874 27806 15876 27858
rect 15820 27794 15876 27806
rect 15820 26180 15876 26190
rect 15820 26086 15876 26124
rect 15596 24892 15764 24948
rect 15820 25060 15876 25070
rect 15596 24724 15652 24892
rect 15596 24668 15764 24724
rect 15316 24332 15540 24388
rect 15596 24498 15652 24510
rect 15596 24446 15598 24498
rect 15650 24446 15652 24498
rect 15148 23380 15204 23390
rect 15148 23042 15204 23324
rect 15148 22990 15150 23042
rect 15202 22990 15204 23042
rect 15148 22978 15204 22990
rect 15260 21588 15316 24332
rect 15596 24164 15652 24446
rect 15596 24098 15652 24108
rect 15484 23938 15540 23950
rect 15484 23886 15486 23938
rect 15538 23886 15540 23938
rect 15372 23716 15428 23726
rect 15372 22260 15428 23660
rect 15372 22036 15428 22204
rect 15372 21970 15428 21980
rect 14924 21026 15092 21028
rect 14924 20974 14926 21026
rect 14978 20974 15092 21026
rect 14924 20972 15092 20974
rect 15148 21586 15316 21588
rect 15148 21534 15262 21586
rect 15314 21534 15316 21586
rect 15148 21532 15316 21534
rect 14924 20962 14980 20972
rect 14700 20178 14756 20188
rect 14924 20804 14980 20814
rect 13916 19684 13972 20132
rect 14140 20020 14196 20030
rect 13580 19170 13636 19180
rect 13692 19628 13972 19684
rect 14028 19908 14084 19918
rect 14028 19684 14084 19852
rect 12684 18844 12964 18900
rect 12124 18788 12180 18798
rect 12124 18674 12180 18732
rect 12124 18622 12126 18674
rect 12178 18622 12180 18674
rect 12124 18610 12180 18622
rect 12684 17890 12740 18844
rect 13356 18676 13412 18686
rect 13020 18564 13076 18574
rect 13356 18564 13412 18620
rect 13020 18562 13524 18564
rect 13020 18510 13022 18562
rect 13074 18510 13524 18562
rect 13020 18508 13524 18510
rect 13020 18498 13076 18508
rect 12684 17838 12686 17890
rect 12738 17838 12740 17890
rect 12124 17666 12180 17678
rect 12124 17614 12126 17666
rect 12178 17614 12180 17666
rect 12124 17108 12180 17614
rect 12124 17042 12180 17052
rect 12012 16830 12014 16882
rect 12066 16830 12068 16882
rect 12012 14532 12068 16830
rect 12572 16660 12628 16670
rect 12124 16548 12180 16558
rect 12124 15538 12180 16492
rect 12124 15486 12126 15538
rect 12178 15486 12180 15538
rect 12124 15474 12180 15486
rect 12572 15540 12628 16604
rect 12460 15316 12516 15326
rect 12460 14754 12516 15260
rect 12460 14702 12462 14754
rect 12514 14702 12516 14754
rect 12460 14690 12516 14702
rect 12012 14466 12068 14476
rect 12460 14532 12516 14542
rect 12012 14196 12068 14206
rect 12012 13746 12068 14140
rect 12012 13694 12014 13746
rect 12066 13694 12068 13746
rect 12012 13682 12068 13694
rect 12236 12850 12292 12862
rect 12236 12798 12238 12850
rect 12290 12798 12292 12850
rect 12012 12516 12068 12526
rect 12012 12290 12068 12460
rect 12012 12238 12014 12290
rect 12066 12238 12068 12290
rect 12012 12226 12068 12238
rect 12236 12292 12292 12798
rect 12460 12628 12516 14476
rect 12572 12852 12628 15484
rect 12684 13412 12740 17838
rect 12908 18340 12964 18350
rect 12796 16884 12852 16894
rect 12796 16322 12852 16828
rect 12796 16270 12798 16322
rect 12850 16270 12852 16322
rect 12796 16258 12852 16270
rect 12796 13858 12852 13870
rect 12796 13806 12798 13858
rect 12850 13806 12852 13858
rect 12796 13524 12852 13806
rect 12908 13634 12964 18284
rect 13356 18340 13412 18350
rect 13356 18246 13412 18284
rect 13468 16098 13524 18508
rect 13468 16046 13470 16098
rect 13522 16046 13524 16098
rect 13468 16034 13524 16046
rect 13580 16772 13636 16782
rect 13468 15876 13524 15886
rect 13132 14420 13188 14430
rect 13132 14326 13188 14364
rect 12908 13582 12910 13634
rect 12962 13582 12964 13634
rect 12908 13570 12964 13582
rect 13132 13636 13188 13646
rect 13132 13634 13412 13636
rect 13132 13582 13134 13634
rect 13186 13582 13412 13634
rect 13132 13580 13412 13582
rect 13132 13570 13188 13580
rect 12796 13458 12852 13468
rect 12684 13346 12740 13356
rect 12908 13412 12964 13422
rect 12684 13076 12740 13086
rect 12684 12982 12740 13020
rect 12572 12786 12628 12796
rect 12460 12572 12628 12628
rect 12292 12236 12516 12292
rect 12236 12226 12292 12236
rect 11452 10558 11454 10610
rect 11506 10558 11508 10610
rect 11452 10276 11508 10558
rect 11452 10210 11508 10220
rect 11564 10668 11732 10724
rect 11788 10780 11956 10836
rect 12012 11394 12068 11406
rect 12012 11342 12014 11394
rect 12066 11342 12068 11394
rect 12012 10834 12068 11342
rect 12460 11394 12516 12236
rect 12460 11342 12462 11394
rect 12514 11342 12516 11394
rect 12460 11330 12516 11342
rect 12012 10782 12014 10834
rect 12066 10782 12068 10834
rect 11340 9774 11342 9826
rect 11394 9774 11396 9826
rect 11340 9156 11396 9774
rect 11340 9090 11396 9100
rect 11004 8988 11284 9044
rect 10892 8878 10894 8930
rect 10946 8878 10948 8930
rect 10892 8820 10948 8878
rect 10892 8754 10948 8764
rect 11116 8372 11172 8382
rect 10892 7700 10948 7710
rect 10780 7698 10948 7700
rect 10780 7646 10894 7698
rect 10946 7646 10948 7698
rect 10780 7644 10948 7646
rect 10892 7634 10948 7644
rect 10668 7298 10724 7308
rect 11004 7364 11060 7374
rect 11004 6804 11060 7308
rect 11004 6690 11060 6748
rect 11004 6638 11006 6690
rect 11058 6638 11060 6690
rect 11004 6626 11060 6638
rect 11116 5348 11172 8316
rect 11228 7252 11284 8988
rect 11564 8708 11620 10668
rect 11676 10498 11732 10510
rect 11676 10446 11678 10498
rect 11730 10446 11732 10498
rect 11676 10164 11732 10446
rect 11676 10098 11732 10108
rect 11564 8642 11620 8652
rect 11228 7186 11284 7196
rect 11564 6692 11620 6702
rect 11564 6598 11620 6636
rect 11116 5282 11172 5292
rect 11564 5682 11620 5694
rect 11564 5630 11566 5682
rect 11618 5630 11620 5682
rect 11564 5348 11620 5630
rect 11564 5282 11620 5292
rect 11564 4564 11620 4574
rect 11452 2100 11508 2110
rect 10332 2098 11508 2100
rect 10332 2046 11454 2098
rect 11506 2046 11508 2098
rect 10332 2044 11508 2046
rect 11452 2034 11508 2044
rect 11564 1092 11620 4508
rect 11788 3388 11844 10780
rect 12012 10770 12068 10782
rect 12124 10836 12180 10846
rect 11900 10610 11956 10622
rect 11900 10558 11902 10610
rect 11954 10558 11956 10610
rect 11900 9940 11956 10558
rect 12124 10610 12180 10780
rect 12124 10558 12126 10610
rect 12178 10558 12180 10610
rect 12124 10546 12180 10558
rect 12236 10612 12292 10622
rect 11900 9874 11956 9884
rect 12012 10500 12068 10510
rect 12012 6018 12068 10444
rect 12236 10386 12292 10556
rect 12236 10334 12238 10386
rect 12290 10334 12292 10386
rect 12236 10322 12292 10334
rect 12348 10276 12404 10286
rect 12124 9940 12180 9950
rect 12124 9268 12180 9884
rect 12236 9826 12292 9838
rect 12236 9774 12238 9826
rect 12290 9774 12292 9826
rect 12236 9492 12292 9774
rect 12236 9426 12292 9436
rect 12348 9604 12404 10220
rect 12124 9212 12292 9268
rect 12124 8932 12180 8942
rect 12124 7474 12180 8876
rect 12236 8482 12292 9212
rect 12348 8932 12404 9548
rect 12348 8866 12404 8876
rect 12460 9268 12516 9278
rect 12236 8430 12238 8482
rect 12290 8430 12292 8482
rect 12236 8418 12292 8430
rect 12460 8260 12516 9212
rect 12236 8204 12516 8260
rect 12236 7698 12292 8204
rect 12572 8148 12628 12572
rect 12796 12516 12852 12526
rect 12796 10836 12852 12460
rect 12796 10770 12852 10780
rect 12796 10610 12852 10622
rect 12796 10558 12798 10610
rect 12850 10558 12852 10610
rect 12684 10052 12740 10062
rect 12796 10052 12852 10558
rect 12684 10050 12852 10052
rect 12684 9998 12686 10050
rect 12738 9998 12852 10050
rect 12684 9996 12852 9998
rect 12684 9986 12740 9996
rect 12236 7646 12238 7698
rect 12290 7646 12292 7698
rect 12236 7634 12292 7646
rect 12348 8092 12628 8148
rect 12796 9044 12852 9054
rect 12348 7476 12404 8092
rect 12124 7422 12126 7474
rect 12178 7422 12180 7474
rect 12124 7410 12180 7422
rect 12236 7420 12404 7476
rect 12796 7476 12852 8988
rect 12908 8932 12964 13356
rect 13244 13412 13300 13422
rect 13020 12852 13076 12862
rect 13020 12402 13076 12796
rect 13020 12350 13022 12402
rect 13074 12350 13076 12402
rect 13020 12338 13076 12350
rect 13020 11506 13076 11518
rect 13020 11454 13022 11506
rect 13074 11454 13076 11506
rect 13020 11172 13076 11454
rect 13020 11106 13076 11116
rect 13244 11172 13300 13356
rect 13356 11732 13412 13580
rect 13356 11666 13412 11676
rect 13468 11508 13524 15820
rect 13580 14754 13636 16716
rect 13580 14702 13582 14754
rect 13634 14702 13636 14754
rect 13580 14690 13636 14702
rect 13244 11106 13300 11116
rect 13356 11452 13524 11508
rect 13692 13634 13748 19628
rect 14028 19618 14084 19628
rect 13916 19236 13972 19246
rect 13804 19234 13972 19236
rect 13804 19182 13918 19234
rect 13970 19182 13972 19234
rect 13804 19180 13972 19182
rect 13804 17890 13860 19180
rect 13916 19170 13972 19180
rect 13804 17838 13806 17890
rect 13858 17838 13860 17890
rect 13804 17826 13860 17838
rect 14140 16660 14196 19964
rect 14476 20020 14532 20030
rect 14812 20020 14868 20030
rect 14476 20018 14644 20020
rect 14476 19966 14478 20018
rect 14530 19966 14644 20018
rect 14476 19964 14644 19966
rect 14476 19954 14532 19964
rect 14476 19234 14532 19246
rect 14476 19182 14478 19234
rect 14530 19182 14532 19234
rect 14476 19012 14532 19182
rect 14476 18946 14532 18956
rect 14588 18674 14644 19964
rect 14700 20018 14868 20020
rect 14700 19966 14814 20018
rect 14866 19966 14868 20018
rect 14700 19964 14868 19966
rect 14700 19234 14756 19964
rect 14812 19954 14868 19964
rect 14924 20020 14980 20748
rect 15148 20356 15204 21532
rect 15260 21522 15316 21532
rect 15484 21474 15540 23886
rect 15484 21422 15486 21474
rect 15538 21422 15540 21474
rect 15484 21410 15540 21422
rect 15708 21252 15764 24668
rect 15148 20290 15204 20300
rect 15260 21196 15764 21252
rect 14924 19954 14980 19964
rect 15036 20018 15092 20030
rect 15036 19966 15038 20018
rect 15090 19966 15092 20018
rect 15036 19908 15092 19966
rect 15036 19842 15092 19852
rect 14700 19182 14702 19234
rect 14754 19182 14756 19234
rect 14700 19170 14756 19182
rect 14924 19684 14980 19694
rect 14588 18622 14590 18674
rect 14642 18622 14644 18674
rect 14588 18610 14644 18622
rect 14140 16594 14196 16604
rect 14700 16996 14756 17006
rect 14700 16770 14756 16940
rect 14700 16718 14702 16770
rect 14754 16718 14756 16770
rect 14476 16436 14532 16446
rect 13804 16210 13860 16222
rect 13804 16158 13806 16210
rect 13858 16158 13860 16210
rect 13804 16100 13860 16158
rect 13804 16034 13860 16044
rect 14364 15988 14420 15998
rect 14364 15314 14420 15932
rect 14364 15262 14366 15314
rect 14418 15262 14420 15314
rect 14364 15250 14420 15262
rect 14476 15540 14532 16380
rect 14476 15148 14532 15484
rect 14700 15204 14756 16718
rect 14028 15092 14084 15102
rect 14476 15092 14644 15148
rect 14700 15110 14756 15148
rect 14924 15148 14980 19628
rect 15260 17554 15316 21196
rect 15260 17502 15262 17554
rect 15314 17502 15316 17554
rect 15260 17490 15316 17502
rect 15372 21028 15428 21038
rect 15036 16884 15092 16894
rect 15036 16790 15092 16828
rect 15036 15876 15092 15886
rect 15036 15782 15092 15820
rect 15148 15316 15204 15326
rect 15148 15222 15204 15260
rect 14924 15092 15092 15148
rect 13916 15090 14084 15092
rect 13916 15038 14030 15090
rect 14082 15038 14084 15090
rect 13916 15036 14084 15038
rect 13692 13582 13694 13634
rect 13746 13582 13748 13634
rect 13692 12516 13748 13582
rect 13804 13636 13860 13646
rect 13804 13186 13860 13580
rect 13804 13134 13806 13186
rect 13858 13134 13860 13186
rect 13804 13122 13860 13134
rect 13916 12740 13972 15036
rect 14028 15026 14084 15036
rect 14364 14420 14420 14430
rect 14140 13746 14196 13758
rect 14140 13694 14142 13746
rect 14194 13694 14196 13746
rect 13916 12674 13972 12684
rect 14028 13524 14084 13534
rect 13244 10724 13300 10734
rect 13244 10630 13300 10668
rect 13020 10612 13076 10622
rect 13020 10518 13076 10556
rect 13132 9940 13188 9950
rect 13132 9846 13188 9884
rect 13244 9826 13300 9838
rect 13244 9774 13246 9826
rect 13298 9774 13300 9826
rect 13244 9268 13300 9774
rect 13244 9202 13300 9212
rect 12908 8876 13300 8932
rect 12908 8372 12964 8382
rect 12908 8148 12964 8316
rect 13244 8372 13300 8876
rect 13356 8596 13412 11452
rect 13692 11396 13748 12460
rect 14028 12178 14084 13468
rect 14028 12126 14030 12178
rect 14082 12126 14084 12178
rect 14028 12114 14084 12126
rect 14140 11618 14196 13694
rect 14364 13524 14420 14364
rect 14364 12962 14420 13468
rect 14364 12910 14366 12962
rect 14418 12910 14420 12962
rect 14364 12898 14420 12910
rect 14588 13746 14644 15092
rect 14700 14644 14756 14654
rect 14700 14550 14756 14588
rect 14588 13694 14590 13746
rect 14642 13694 14644 13746
rect 14140 11566 14142 11618
rect 14194 11566 14196 11618
rect 14140 11554 14196 11566
rect 13692 11340 14196 11396
rect 13468 10612 13524 10622
rect 14028 10612 14084 10622
rect 13468 10610 13972 10612
rect 13468 10558 13470 10610
rect 13522 10558 13972 10610
rect 13468 10556 13972 10558
rect 13468 10546 13524 10556
rect 13580 10386 13636 10398
rect 13580 10334 13582 10386
rect 13634 10334 13636 10386
rect 13356 8530 13412 8540
rect 13468 9826 13524 9838
rect 13468 9774 13470 9826
rect 13522 9774 13524 9826
rect 13468 8372 13524 9774
rect 13244 8370 13412 8372
rect 13244 8318 13246 8370
rect 13298 8318 13412 8370
rect 13244 8316 13412 8318
rect 13244 8306 13300 8316
rect 12908 8146 13076 8148
rect 12908 8094 12910 8146
rect 12962 8094 13076 8146
rect 12908 8092 13076 8094
rect 12908 8082 12964 8092
rect 12908 7476 12964 7486
rect 12796 7474 12964 7476
rect 12796 7422 12910 7474
rect 12962 7422 12964 7474
rect 12796 7420 12964 7422
rect 12012 5966 12014 6018
rect 12066 5966 12068 6018
rect 12012 5954 12068 5966
rect 12236 5908 12292 7420
rect 12796 7140 12852 7420
rect 12908 7410 12964 7420
rect 12348 7084 12852 7140
rect 12348 6690 12404 7084
rect 13020 7028 13076 8092
rect 13356 7364 13412 8316
rect 13468 8306 13524 8316
rect 13580 7476 13636 10334
rect 13692 10388 13748 10398
rect 13692 10294 13748 10332
rect 13916 10050 13972 10556
rect 13916 9998 13918 10050
rect 13970 9998 13972 10050
rect 13916 9986 13972 9998
rect 13804 9940 13860 9950
rect 13804 9826 13860 9884
rect 14028 9828 14084 10556
rect 13804 9774 13806 9826
rect 13858 9774 13860 9826
rect 13804 9762 13860 9774
rect 13916 9772 14084 9828
rect 13804 9268 13860 9278
rect 13916 9268 13972 9772
rect 14028 9604 14084 9614
rect 14028 9510 14084 9548
rect 13804 9266 13972 9268
rect 13804 9214 13806 9266
rect 13858 9214 13972 9266
rect 13804 9212 13972 9214
rect 13804 9202 13860 9212
rect 13580 7410 13636 7420
rect 13916 8484 13972 8494
rect 13020 6962 13076 6972
rect 13132 7362 13412 7364
rect 13132 7310 13358 7362
rect 13410 7310 13412 7362
rect 13132 7308 13412 7310
rect 12684 6804 12740 6814
rect 12684 6710 12740 6748
rect 12348 6638 12350 6690
rect 12402 6638 12404 6690
rect 12348 6626 12404 6638
rect 13132 6356 13188 7308
rect 13356 7298 13412 7308
rect 12236 5842 12292 5852
rect 12348 6300 13188 6356
rect 13244 7140 13300 7150
rect 12348 5122 12404 6300
rect 12796 5236 12852 5246
rect 13244 5236 13300 7084
rect 12796 5234 13300 5236
rect 12796 5182 12798 5234
rect 12850 5182 13300 5234
rect 12796 5180 13300 5182
rect 13356 7028 13412 7038
rect 12796 5170 12852 5180
rect 12348 5070 12350 5122
rect 12402 5070 12404 5122
rect 12348 5058 12404 5070
rect 13356 5122 13412 6972
rect 13916 6914 13972 8428
rect 13916 6862 13918 6914
rect 13970 6862 13972 6914
rect 13916 6850 13972 6862
rect 13804 6020 13860 6030
rect 14140 6020 14196 11340
rect 14588 10388 14644 13694
rect 14700 13972 14756 13982
rect 14700 13634 14756 13916
rect 14700 13582 14702 13634
rect 14754 13582 14756 13634
rect 14700 13570 14756 13582
rect 14812 13524 14868 13534
rect 14812 12178 14868 13468
rect 14924 13074 14980 13086
rect 14924 13022 14926 13074
rect 14978 13022 14980 13074
rect 14924 12404 14980 13022
rect 14924 12338 14980 12348
rect 14812 12126 14814 12178
rect 14866 12126 14868 12178
rect 14700 10724 14756 10734
rect 14812 10724 14868 12126
rect 14700 10722 14868 10724
rect 14700 10670 14702 10722
rect 14754 10670 14868 10722
rect 14700 10668 14868 10670
rect 14700 10658 14756 10668
rect 14812 10612 14868 10668
rect 14588 10332 14756 10388
rect 14588 10052 14644 10062
rect 14252 9602 14308 9614
rect 14252 9550 14254 9602
rect 14306 9550 14308 9602
rect 14252 8260 14308 9550
rect 14252 8194 14308 8204
rect 14476 8036 14532 8046
rect 13804 6018 14196 6020
rect 13804 5966 13806 6018
rect 13858 5966 14196 6018
rect 13804 5964 14196 5966
rect 14252 8034 14532 8036
rect 14252 7982 14478 8034
rect 14530 7982 14532 8034
rect 14252 7980 14532 7982
rect 13804 5954 13860 5964
rect 14252 5906 14308 7980
rect 14476 7970 14532 7980
rect 14588 7700 14644 9996
rect 14252 5854 14254 5906
rect 14306 5854 14308 5906
rect 14252 5842 14308 5854
rect 14476 7644 14644 7700
rect 13804 5348 13860 5358
rect 13804 5254 13860 5292
rect 14476 5348 14532 7644
rect 14588 7476 14644 7486
rect 14588 7382 14644 7420
rect 14700 5906 14756 10332
rect 14812 9042 14868 10556
rect 15036 10498 15092 15092
rect 15148 14530 15204 14542
rect 15148 14478 15150 14530
rect 15202 14478 15204 14530
rect 15148 13972 15204 14478
rect 15148 13906 15204 13916
rect 15260 13748 15316 13758
rect 15372 13748 15428 20972
rect 15596 20804 15652 20814
rect 15484 19236 15540 19246
rect 15484 19142 15540 19180
rect 15484 16884 15540 16894
rect 15596 16884 15652 20748
rect 15820 20018 15876 25004
rect 15932 21028 15988 31948
rect 16044 29426 16100 38612
rect 16380 38610 16436 38622
rect 16380 38558 16382 38610
rect 16434 38558 16436 38610
rect 16156 37042 16212 37054
rect 16156 36990 16158 37042
rect 16210 36990 16212 37042
rect 16156 36708 16212 36990
rect 16156 36642 16212 36652
rect 16044 29374 16046 29426
rect 16098 29374 16100 29426
rect 16044 29362 16100 29374
rect 16268 34916 16324 34926
rect 16268 33906 16324 34860
rect 16268 33854 16270 33906
rect 16322 33854 16324 33906
rect 16268 30994 16324 33854
rect 16380 32228 16436 38558
rect 16604 37266 16660 40124
rect 16604 37214 16606 37266
rect 16658 37214 16660 37266
rect 16604 37202 16660 37214
rect 16380 32162 16436 32172
rect 16492 37156 16548 37166
rect 16492 31892 16548 37100
rect 16716 36932 16772 41804
rect 16940 38946 16996 46060
rect 16940 38894 16942 38946
rect 16994 38894 16996 38946
rect 16940 38882 16996 38894
rect 17164 37380 17220 37390
rect 17164 37266 17220 37324
rect 17164 37214 17166 37266
rect 17218 37214 17220 37266
rect 17164 37202 17220 37214
rect 16604 36876 16772 36932
rect 16604 35252 16660 36876
rect 16716 36708 16772 36718
rect 16716 36614 16772 36652
rect 17276 36596 17332 53564
rect 16604 35186 16660 35196
rect 17164 36540 17332 36596
rect 17388 39060 17444 39070
rect 16268 30942 16270 30994
rect 16322 30942 16324 30994
rect 16044 28644 16100 28654
rect 16044 28550 16100 28588
rect 16268 26852 16324 30942
rect 16380 31836 16548 31892
rect 17052 34692 17108 34702
rect 16380 29652 16436 31836
rect 16716 31780 16772 31790
rect 16492 31778 16772 31780
rect 16492 31726 16718 31778
rect 16770 31726 16772 31778
rect 16492 31724 16772 31726
rect 16492 30882 16548 31724
rect 16716 31714 16772 31724
rect 16828 31780 16884 31790
rect 16492 30830 16494 30882
rect 16546 30830 16548 30882
rect 16492 30818 16548 30830
rect 16716 29652 16772 29662
rect 16380 29596 16548 29652
rect 16044 25282 16100 25294
rect 16044 25230 16046 25282
rect 16098 25230 16100 25282
rect 16044 24722 16100 25230
rect 16044 24670 16046 24722
rect 16098 24670 16100 24722
rect 16044 24658 16100 24670
rect 16044 24500 16100 24510
rect 16044 24050 16100 24444
rect 16044 23998 16046 24050
rect 16098 23998 16100 24050
rect 16044 23986 16100 23998
rect 16268 23604 16324 26796
rect 16156 23548 16324 23604
rect 16380 29428 16436 29438
rect 16156 23156 16212 23548
rect 16268 23380 16324 23390
rect 16268 23286 16324 23324
rect 16156 23100 16324 23156
rect 16044 22146 16100 22158
rect 16044 22094 16046 22146
rect 16098 22094 16100 22146
rect 16044 21924 16100 22094
rect 16044 21858 16100 21868
rect 16156 22148 16212 22158
rect 16156 21586 16212 22092
rect 16156 21534 16158 21586
rect 16210 21534 16212 21586
rect 16156 21522 16212 21534
rect 15932 20962 15988 20972
rect 16044 21252 16100 21262
rect 16044 20914 16100 21196
rect 16044 20862 16046 20914
rect 16098 20862 16100 20914
rect 16044 20850 16100 20862
rect 16268 20804 16324 23100
rect 16268 20738 16324 20748
rect 16380 21588 16436 29372
rect 16492 28868 16548 29596
rect 16492 28802 16548 28812
rect 16604 27860 16660 27870
rect 16604 27766 16660 27804
rect 16604 27524 16660 27534
rect 16604 24722 16660 27468
rect 16604 24670 16606 24722
rect 16658 24670 16660 24722
rect 16604 24658 16660 24670
rect 16716 27188 16772 29596
rect 16716 23828 16772 27132
rect 16828 26068 16884 31724
rect 16940 30884 16996 30894
rect 16940 30790 16996 30828
rect 17052 30436 17108 34636
rect 17164 31668 17220 36540
rect 17276 36370 17332 36382
rect 17276 36318 17278 36370
rect 17330 36318 17332 36370
rect 17276 35812 17332 36318
rect 17276 35746 17332 35756
rect 17388 35140 17444 39004
rect 17500 37380 17556 55918
rect 19516 55970 19572 55982
rect 19516 55918 19518 55970
rect 19570 55918 19572 55970
rect 18284 55300 18340 55310
rect 18284 55206 18340 55244
rect 19068 54290 19124 54302
rect 19068 54238 19070 54290
rect 19122 54238 19124 54290
rect 17500 37314 17556 37324
rect 17948 46564 18004 46574
rect 17276 35084 17444 35140
rect 17500 36596 17556 36606
rect 17500 35364 17556 36540
rect 17276 31890 17332 35084
rect 17500 34914 17556 35308
rect 17500 34862 17502 34914
rect 17554 34862 17556 34914
rect 17500 34850 17556 34862
rect 17724 36482 17780 36494
rect 17724 36430 17726 36482
rect 17778 36430 17780 36482
rect 17276 31838 17278 31890
rect 17330 31838 17332 31890
rect 17276 31826 17332 31838
rect 17388 34132 17444 34142
rect 17724 34132 17780 36430
rect 17948 35026 18004 46508
rect 19068 43708 19124 54238
rect 19516 43708 19572 55918
rect 19628 55972 19684 55982
rect 19628 54626 19684 55916
rect 21308 55972 21364 55982
rect 21308 55878 21364 55916
rect 21644 55860 21700 55870
rect 21644 55410 21700 55804
rect 21644 55358 21646 55410
rect 21698 55358 21700 55410
rect 21644 55346 21700 55358
rect 19628 54574 19630 54626
rect 19682 54574 19684 54626
rect 19628 54562 19684 54574
rect 19964 55298 20020 55310
rect 19964 55246 19966 55298
rect 20018 55246 20020 55298
rect 19964 48132 20020 55246
rect 20524 55300 20580 55310
rect 20524 55206 20580 55244
rect 20860 55298 20916 55310
rect 20860 55246 20862 55298
rect 20914 55246 20916 55298
rect 20636 54292 20692 54302
rect 20636 54198 20692 54236
rect 20860 53844 20916 55246
rect 21196 54516 21252 54526
rect 21196 54422 21252 54460
rect 20860 53778 20916 53788
rect 21532 54402 21588 54414
rect 21532 54350 21534 54402
rect 21586 54350 21588 54402
rect 21420 52164 21476 52174
rect 21420 52070 21476 52108
rect 19964 48066 20020 48076
rect 18620 43652 19124 43708
rect 19180 43652 19572 43708
rect 19740 47348 19796 47358
rect 18396 40180 18452 40190
rect 18172 37266 18228 37278
rect 18172 37214 18174 37266
rect 18226 37214 18228 37266
rect 17948 34974 17950 35026
rect 18002 34974 18004 35026
rect 17948 34962 18004 34974
rect 18060 35364 18116 35374
rect 17388 34130 17780 34132
rect 17388 34078 17390 34130
rect 17442 34078 17780 34130
rect 17388 34076 17780 34078
rect 17836 34244 17892 34254
rect 17164 31612 17332 31668
rect 17052 30380 17220 30436
rect 17052 30212 17108 30222
rect 16940 30156 17052 30212
rect 16940 29540 16996 30156
rect 17052 30118 17108 30156
rect 16940 29474 16996 29484
rect 17052 29876 17108 29886
rect 17052 26404 17108 29820
rect 17164 27636 17220 30380
rect 17276 29764 17332 31612
rect 17388 29988 17444 34076
rect 17836 34018 17892 34188
rect 17836 33966 17838 34018
rect 17890 33966 17892 34018
rect 17724 33796 17780 33806
rect 17500 33684 17556 33694
rect 17500 30548 17556 33628
rect 17500 30434 17556 30492
rect 17500 30382 17502 30434
rect 17554 30382 17556 30434
rect 17500 30370 17556 30382
rect 17724 30994 17780 33740
rect 17836 33684 17892 33966
rect 17836 33618 17892 33628
rect 18060 32004 18116 35308
rect 17724 30942 17726 30994
rect 17778 30942 17780 30994
rect 17724 30324 17780 30942
rect 17724 30258 17780 30268
rect 17948 31948 18060 32004
rect 17388 29922 17444 29932
rect 17724 29988 17780 29998
rect 17276 29708 17668 29764
rect 17500 29426 17556 29438
rect 17500 29374 17502 29426
rect 17554 29374 17556 29426
rect 17388 28532 17444 28542
rect 17388 28438 17444 28476
rect 17164 27570 17220 27580
rect 17388 27188 17444 27198
rect 17388 27094 17444 27132
rect 17052 26338 17108 26348
rect 17500 26740 17556 29374
rect 16828 26002 16884 26012
rect 17276 26066 17332 26078
rect 17276 26014 17278 26066
rect 17330 26014 17332 26066
rect 17276 25732 17332 26014
rect 17276 25666 17332 25676
rect 17388 26068 17444 26078
rect 16828 25506 16884 25518
rect 16828 25454 16830 25506
rect 16882 25454 16884 25506
rect 16828 24164 16884 25454
rect 17276 25508 17332 25518
rect 17388 25508 17444 26012
rect 17500 25620 17556 26684
rect 17612 26404 17668 29708
rect 17724 27074 17780 29932
rect 17836 28868 17892 28878
rect 17948 28868 18004 31948
rect 18060 31938 18116 31948
rect 18060 31780 18116 31790
rect 18060 31686 18116 31724
rect 17836 28866 17948 28868
rect 17836 28814 17838 28866
rect 17890 28814 17948 28866
rect 17836 28812 17948 28814
rect 17836 28802 17892 28812
rect 17948 28774 18004 28812
rect 18060 29426 18116 29438
rect 18060 29374 18062 29426
rect 18114 29374 18116 29426
rect 18060 29316 18116 29374
rect 17724 27022 17726 27074
rect 17778 27022 17780 27074
rect 17724 27010 17780 27022
rect 17836 27860 17892 27870
rect 17724 26404 17780 26414
rect 17612 26402 17780 26404
rect 17612 26350 17726 26402
rect 17778 26350 17780 26402
rect 17612 26348 17780 26350
rect 17724 26338 17780 26348
rect 17500 25554 17556 25564
rect 17276 25506 17444 25508
rect 17276 25454 17278 25506
rect 17330 25454 17444 25506
rect 17276 25452 17444 25454
rect 17276 25442 17332 25452
rect 17836 25396 17892 27804
rect 18060 27858 18116 29260
rect 18060 27806 18062 27858
rect 18114 27806 18116 27858
rect 18060 27794 18116 27806
rect 18172 27860 18228 37214
rect 18284 36596 18340 36606
rect 18284 36502 18340 36540
rect 18284 34804 18340 34814
rect 18284 33796 18340 34748
rect 18284 33730 18340 33740
rect 18396 33460 18452 40124
rect 18172 27794 18228 27804
rect 18284 33404 18452 33460
rect 17500 25340 17892 25396
rect 18060 27636 18116 27646
rect 17500 24717 17556 25340
rect 17500 24665 17502 24717
rect 17554 24665 17556 24717
rect 17500 24500 17556 24665
rect 18060 24612 18116 27580
rect 18172 27074 18228 27086
rect 18172 27022 18174 27074
rect 18226 27022 18228 27074
rect 18172 25396 18228 27022
rect 18284 26068 18340 33404
rect 18396 33234 18452 33246
rect 18396 33182 18398 33234
rect 18450 33182 18452 33234
rect 18396 31780 18452 33182
rect 18620 32116 18676 43652
rect 18732 34916 18788 34926
rect 19068 34916 19124 34926
rect 18732 34914 19012 34916
rect 18732 34862 18734 34914
rect 18786 34862 19012 34914
rect 18732 34860 19012 34862
rect 18732 34850 18788 34860
rect 18956 34354 19012 34860
rect 19068 34822 19124 34860
rect 18956 34302 18958 34354
rect 19010 34302 19012 34354
rect 18956 34290 19012 34302
rect 18732 33572 18788 33582
rect 19180 33572 19236 43652
rect 19404 36260 19460 36270
rect 19404 36166 19460 36204
rect 19292 35028 19348 35038
rect 19292 35026 19572 35028
rect 19292 34974 19294 35026
rect 19346 34974 19572 35026
rect 19292 34972 19572 34974
rect 19292 34962 19348 34972
rect 19516 34130 19572 34972
rect 19516 34078 19518 34130
rect 19570 34078 19572 34130
rect 19516 34066 19572 34078
rect 18732 33458 18788 33516
rect 18732 33406 18734 33458
rect 18786 33406 18788 33458
rect 18732 33394 18788 33406
rect 18844 33516 19236 33572
rect 19292 33572 19348 33582
rect 18620 32060 18788 32116
rect 18508 32004 18564 32014
rect 18508 31890 18564 31948
rect 18508 31838 18510 31890
rect 18562 31838 18564 31890
rect 18508 31826 18564 31838
rect 18396 31714 18452 31724
rect 18508 30996 18564 31006
rect 18508 30902 18564 30940
rect 18508 30548 18564 30558
rect 18508 29314 18564 30492
rect 18620 29988 18676 29998
rect 18620 29894 18676 29932
rect 18508 29262 18510 29314
rect 18562 29262 18564 29314
rect 18508 29250 18564 29262
rect 18508 28868 18564 28878
rect 18508 27746 18564 28812
rect 18732 28420 18788 32060
rect 18844 29204 18900 33516
rect 18956 33236 19012 33246
rect 18956 29988 19012 33180
rect 19292 32562 19348 33516
rect 19740 32674 19796 47292
rect 20188 44324 20244 44334
rect 19852 41972 19908 41982
rect 19852 36594 19908 41916
rect 20076 41300 20132 41310
rect 19852 36542 19854 36594
rect 19906 36542 19908 36594
rect 19852 36530 19908 36542
rect 19964 38724 20020 38734
rect 19852 36260 19908 36270
rect 19852 34914 19908 36204
rect 19852 34862 19854 34914
rect 19906 34862 19908 34914
rect 19852 34850 19908 34862
rect 19964 34468 20020 38668
rect 19964 34402 20020 34412
rect 20076 34244 20132 41244
rect 20188 35700 20244 44268
rect 21084 40068 21140 40078
rect 20748 38052 20804 38062
rect 20188 35634 20244 35644
rect 20412 36482 20468 36494
rect 20412 36430 20414 36482
rect 20466 36430 20468 36482
rect 19740 32622 19742 32674
rect 19794 32622 19796 32674
rect 19740 32610 19796 32622
rect 19852 34188 20132 34244
rect 19292 32510 19294 32562
rect 19346 32510 19348 32562
rect 19292 32498 19348 32510
rect 19740 31554 19796 31566
rect 19740 31502 19742 31554
rect 19794 31502 19796 31554
rect 19740 30996 19796 31502
rect 19740 30930 19796 30940
rect 19740 30436 19796 30446
rect 19852 30436 19908 34188
rect 20076 34018 20132 34030
rect 20076 33966 20078 34018
rect 20130 33966 20132 34018
rect 19964 33122 20020 33134
rect 19964 33070 19966 33122
rect 20018 33070 20020 33122
rect 19964 31108 20020 33070
rect 19964 31042 20020 31052
rect 19740 30434 19908 30436
rect 19740 30382 19742 30434
rect 19794 30382 19908 30434
rect 19740 30380 19908 30382
rect 19292 30212 19348 30222
rect 19292 30118 19348 30156
rect 18956 29922 19012 29932
rect 19068 30100 19124 30110
rect 18844 29138 18900 29148
rect 18732 28354 18788 28364
rect 18956 28418 19012 28430
rect 18956 28366 18958 28418
rect 19010 28366 19012 28418
rect 18508 27694 18510 27746
rect 18562 27694 18564 27746
rect 18508 27682 18564 27694
rect 18396 27188 18452 27198
rect 18396 27186 18676 27188
rect 18396 27134 18398 27186
rect 18450 27134 18676 27186
rect 18396 27132 18676 27134
rect 18396 27122 18452 27132
rect 18284 26002 18340 26012
rect 18396 26404 18452 26414
rect 18396 25396 18452 26348
rect 18620 25730 18676 27132
rect 18956 27074 19012 28366
rect 18956 27022 18958 27074
rect 19010 27022 19012 27074
rect 18956 27010 19012 27022
rect 18620 25678 18622 25730
rect 18674 25678 18676 25730
rect 18620 25666 18676 25678
rect 18732 26178 18788 26190
rect 18732 26126 18734 26178
rect 18786 26126 18788 26178
rect 18732 25732 18788 26126
rect 18956 25732 19012 25742
rect 18732 25666 18788 25676
rect 18844 25676 18956 25732
rect 18172 25340 18340 25396
rect 16828 24098 16884 24108
rect 17388 24444 17556 24500
rect 17612 24556 18116 24612
rect 17388 24388 17444 24444
rect 17164 24052 17220 24062
rect 16716 23734 16772 23772
rect 17052 23938 17108 23950
rect 17052 23886 17054 23938
rect 17106 23886 17108 23938
rect 17052 23380 17108 23886
rect 17052 23314 17108 23324
rect 16828 22148 16884 22158
rect 16828 22054 16884 22092
rect 16492 21588 16548 21598
rect 16380 21586 16548 21588
rect 16380 21534 16494 21586
rect 16546 21534 16548 21586
rect 16380 21532 16548 21534
rect 15820 19966 15822 20018
rect 15874 19966 15876 20018
rect 15820 19572 15876 19966
rect 15820 19236 15876 19516
rect 16268 20580 16324 20590
rect 15820 19170 15876 19180
rect 15932 19348 15988 19358
rect 15820 18450 15876 18462
rect 15820 18398 15822 18450
rect 15874 18398 15876 18450
rect 15484 16882 15652 16884
rect 15484 16830 15486 16882
rect 15538 16830 15652 16882
rect 15484 16828 15652 16830
rect 15708 17666 15764 17678
rect 15708 17614 15710 17666
rect 15762 17614 15764 17666
rect 15484 15314 15540 16828
rect 15708 16770 15764 17614
rect 15820 17332 15876 18398
rect 15820 17266 15876 17276
rect 15708 16718 15710 16770
rect 15762 16718 15764 16770
rect 15708 16706 15764 16718
rect 15820 17108 15876 17118
rect 15484 15262 15486 15314
rect 15538 15262 15540 15314
rect 15484 15250 15540 15262
rect 15596 16098 15652 16110
rect 15596 16046 15598 16098
rect 15650 16046 15652 16098
rect 15596 15204 15652 16046
rect 15708 15204 15764 15214
rect 15596 15202 15764 15204
rect 15596 15150 15710 15202
rect 15762 15150 15764 15202
rect 15596 15148 15764 15150
rect 15708 15138 15764 15148
rect 15708 14644 15764 14654
rect 15820 14644 15876 17052
rect 15708 14642 15876 14644
rect 15708 14590 15710 14642
rect 15762 14590 15876 14642
rect 15708 14588 15876 14590
rect 15708 14578 15764 14588
rect 15708 13748 15764 13758
rect 15372 13746 15764 13748
rect 15372 13694 15710 13746
rect 15762 13694 15764 13746
rect 15372 13692 15764 13694
rect 15148 13636 15204 13646
rect 15148 13542 15204 13580
rect 15260 12066 15316 13692
rect 15260 12014 15262 12066
rect 15314 12014 15316 12066
rect 15260 12002 15316 12014
rect 15596 11620 15652 11630
rect 15596 11526 15652 11564
rect 15708 11396 15764 13692
rect 15596 11340 15764 11396
rect 15036 10446 15038 10498
rect 15090 10446 15092 10498
rect 15036 10052 15092 10446
rect 15372 11170 15428 11182
rect 15372 11118 15374 11170
rect 15426 11118 15428 11170
rect 15036 9986 15092 9996
rect 15148 10164 15204 10174
rect 15148 9938 15204 10108
rect 15148 9886 15150 9938
rect 15202 9886 15204 9938
rect 15148 9874 15204 9886
rect 15260 10050 15316 10062
rect 15260 9998 15262 10050
rect 15314 9998 15316 10050
rect 14924 9828 14980 9838
rect 14924 9826 15092 9828
rect 14924 9774 14926 9826
rect 14978 9774 15092 9826
rect 14924 9772 15092 9774
rect 14924 9762 14980 9772
rect 14812 8990 14814 9042
rect 14866 8990 14868 9042
rect 14812 8978 14868 8990
rect 15036 9716 15092 9772
rect 15148 9716 15204 9726
rect 15036 9660 15148 9716
rect 14924 8484 14980 8494
rect 15036 8484 15092 9660
rect 15148 9650 15204 9660
rect 14980 8428 15092 8484
rect 14924 8370 14980 8428
rect 14924 8318 14926 8370
rect 14978 8318 14980 8370
rect 14812 8260 14868 8270
rect 14812 7924 14868 8204
rect 14812 7858 14868 7868
rect 14924 7364 14980 8318
rect 15260 8260 15316 9998
rect 15372 9716 15428 11118
rect 15372 9650 15428 9660
rect 15596 9716 15652 11340
rect 15708 11170 15764 11182
rect 15708 11118 15710 11170
rect 15762 11118 15764 11170
rect 15708 9826 15764 11118
rect 15932 10724 15988 19292
rect 16044 19234 16100 19246
rect 16044 19182 16046 19234
rect 16098 19182 16100 19234
rect 16044 19124 16100 19182
rect 16044 19058 16100 19068
rect 16156 19012 16212 19022
rect 16156 18918 16212 18956
rect 16044 18900 16100 18910
rect 16044 16210 16100 18844
rect 16156 17444 16212 17454
rect 16156 16882 16212 17388
rect 16268 17108 16324 20524
rect 16268 17042 16324 17052
rect 16156 16830 16158 16882
rect 16210 16830 16212 16882
rect 16156 16818 16212 16830
rect 16044 16158 16046 16210
rect 16098 16158 16100 16210
rect 16044 16146 16100 16158
rect 16156 15876 16212 15886
rect 16156 15314 16212 15820
rect 16156 15262 16158 15314
rect 16210 15262 16212 15314
rect 16156 15250 16212 15262
rect 16044 14530 16100 14542
rect 16044 14478 16046 14530
rect 16098 14478 16100 14530
rect 16044 13186 16100 14478
rect 16044 13134 16046 13186
rect 16098 13134 16100 13186
rect 16044 12964 16100 13134
rect 16044 12898 16100 12908
rect 16156 14306 16212 14318
rect 16156 14254 16158 14306
rect 16210 14254 16212 14306
rect 16156 12292 16212 14254
rect 16156 12226 16212 12236
rect 16380 11620 16436 21532
rect 16492 21522 16548 21532
rect 17052 21364 17108 21374
rect 17164 21364 17220 23996
rect 17388 22148 17444 24332
rect 17500 24276 17556 24286
rect 17500 23938 17556 24220
rect 17500 23886 17502 23938
rect 17554 23886 17556 23938
rect 17500 23716 17556 23886
rect 17500 23650 17556 23660
rect 17388 22082 17444 22092
rect 17500 21812 17556 21822
rect 17108 21308 17220 21364
rect 17388 21588 17444 21598
rect 16828 20914 16884 20926
rect 16828 20862 16830 20914
rect 16882 20862 16884 20914
rect 16492 20020 16548 20030
rect 16492 19926 16548 19964
rect 16604 18452 16660 18462
rect 16492 18450 16660 18452
rect 16492 18398 16606 18450
rect 16658 18398 16660 18450
rect 16492 18396 16660 18398
rect 16492 15204 16548 18396
rect 16604 18386 16660 18396
rect 16828 18450 16884 20862
rect 17052 19906 17108 21308
rect 17276 21252 17332 21262
rect 17276 20914 17332 21196
rect 17276 20862 17278 20914
rect 17330 20862 17332 20914
rect 17276 20850 17332 20862
rect 17052 19854 17054 19906
rect 17106 19854 17108 19906
rect 17052 19842 17108 19854
rect 17164 20802 17220 20814
rect 17164 20750 17166 20802
rect 17218 20750 17220 20802
rect 17164 19460 17220 20750
rect 17052 19404 17220 19460
rect 17388 19458 17444 21532
rect 17500 21586 17556 21756
rect 17500 21534 17502 21586
rect 17554 21534 17556 21586
rect 17500 21522 17556 21534
rect 17612 21364 17668 24556
rect 18172 24500 18228 24510
rect 17724 24498 18228 24500
rect 17724 24446 18174 24498
rect 18226 24446 18228 24498
rect 17724 24444 18228 24446
rect 17724 24162 17780 24444
rect 18172 24434 18228 24444
rect 17724 24110 17726 24162
rect 17778 24110 17780 24162
rect 17724 24098 17780 24110
rect 18172 23940 18228 23950
rect 18060 23938 18228 23940
rect 18060 23886 18174 23938
rect 18226 23886 18228 23938
rect 18060 23884 18228 23886
rect 18060 22596 18116 23884
rect 18172 23874 18228 23884
rect 18284 23716 18340 25340
rect 18396 25330 18452 25340
rect 18732 24836 18788 24846
rect 18844 24836 18900 25676
rect 18956 25666 19012 25676
rect 18732 24834 18900 24836
rect 18732 24782 18734 24834
rect 18786 24782 18900 24834
rect 18732 24780 18900 24782
rect 18732 24770 18788 24780
rect 19068 24052 19124 30044
rect 19740 30100 19796 30380
rect 19740 30034 19796 30044
rect 20076 30100 20132 33966
rect 20188 31666 20244 31678
rect 20188 31614 20190 31666
rect 20242 31614 20244 31666
rect 20188 30884 20244 31614
rect 20188 30818 20244 30828
rect 20412 30212 20468 36430
rect 20524 34914 20580 34926
rect 20524 34862 20526 34914
rect 20578 34862 20580 34914
rect 20524 31556 20580 34862
rect 20748 32674 20804 37996
rect 20748 32622 20750 32674
rect 20802 32622 20804 32674
rect 20748 32610 20804 32622
rect 20636 31780 20692 31790
rect 20972 31780 21028 31790
rect 20636 31778 20916 31780
rect 20636 31726 20638 31778
rect 20690 31726 20916 31778
rect 20636 31724 20916 31726
rect 20636 31714 20692 31724
rect 20524 31490 20580 31500
rect 20636 30884 20692 30894
rect 20692 30828 20804 30884
rect 20636 30790 20692 30828
rect 20412 30146 20468 30156
rect 20076 30034 20132 30044
rect 19292 29988 19348 29998
rect 19180 28532 19236 28542
rect 19180 25618 19236 28476
rect 19180 25566 19182 25618
rect 19234 25566 19236 25618
rect 19180 25554 19236 25566
rect 19068 23986 19124 23996
rect 18284 23650 18340 23660
rect 18732 23938 18788 23950
rect 18732 23886 18734 23938
rect 18786 23886 18788 23938
rect 18060 22530 18116 22540
rect 18396 23156 18452 23166
rect 17948 22484 18004 22494
rect 17948 22390 18004 22428
rect 18396 22370 18452 23100
rect 18396 22318 18398 22370
rect 18450 22318 18452 22370
rect 18396 22306 18452 22318
rect 18396 22148 18452 22158
rect 18284 21812 18340 21822
rect 18172 21700 18228 21710
rect 17388 19406 17390 19458
rect 17442 19406 17444 19458
rect 16940 19236 16996 19246
rect 17052 19236 17108 19404
rect 17388 19394 17444 19406
rect 17500 21308 17668 21364
rect 17724 21698 18228 21700
rect 17724 21646 18174 21698
rect 18226 21646 18228 21698
rect 17724 21644 18228 21646
rect 16940 19234 17108 19236
rect 16940 19182 16942 19234
rect 16994 19182 17108 19234
rect 16940 19180 17108 19182
rect 17164 19234 17220 19246
rect 17164 19182 17166 19234
rect 17218 19182 17220 19234
rect 16940 19170 16996 19180
rect 16828 18398 16830 18450
rect 16882 18398 16884 18450
rect 16828 18386 16884 18398
rect 17164 19012 17220 19182
rect 17388 19236 17444 19246
rect 17388 19142 17444 19180
rect 16828 17892 16884 17902
rect 16828 17798 16884 17836
rect 16716 17668 16772 17678
rect 16716 17574 16772 17612
rect 16940 17332 16996 17342
rect 16940 16884 16996 17276
rect 16828 16882 16996 16884
rect 16828 16830 16942 16882
rect 16994 16830 16996 16882
rect 16828 16828 16996 16830
rect 16716 16100 16772 16110
rect 16492 15138 16548 15148
rect 16604 16098 16772 16100
rect 16604 16046 16718 16098
rect 16770 16046 16772 16098
rect 16604 16044 16772 16046
rect 16604 13972 16660 16044
rect 16716 16034 16772 16044
rect 16828 15540 16884 16828
rect 16940 16818 16996 16828
rect 17052 16322 17108 16334
rect 17052 16270 17054 16322
rect 17106 16270 17108 16322
rect 16716 15484 16884 15540
rect 16940 16100 16996 16110
rect 16940 15540 16996 16044
rect 17052 15652 17108 16270
rect 17164 15876 17220 18956
rect 17500 18900 17556 21308
rect 17500 18834 17556 18844
rect 17612 20578 17668 20590
rect 17612 20526 17614 20578
rect 17666 20526 17668 20578
rect 17612 19908 17668 20526
rect 17388 18340 17444 18350
rect 17388 18246 17444 18284
rect 17612 18116 17668 19852
rect 17724 19234 17780 21644
rect 18172 21634 18228 21644
rect 18284 21364 18340 21756
rect 18060 21362 18340 21364
rect 18060 21310 18286 21362
rect 18338 21310 18340 21362
rect 18060 21308 18340 21310
rect 17948 21028 18004 21038
rect 17948 20934 18004 20972
rect 17724 19182 17726 19234
rect 17778 19182 17780 19234
rect 17724 19170 17780 19182
rect 17836 19908 17892 19918
rect 17836 18338 17892 19852
rect 17836 18286 17838 18338
rect 17890 18286 17892 18338
rect 17836 18274 17892 18286
rect 17948 18450 18004 18462
rect 17948 18398 17950 18450
rect 18002 18398 18004 18450
rect 17948 18116 18004 18398
rect 17612 18060 18004 18116
rect 17276 17778 17332 17790
rect 17276 17726 17278 17778
rect 17330 17726 17332 17778
rect 17276 17668 17332 17726
rect 17500 17780 17556 17790
rect 17500 17686 17556 17724
rect 17276 16884 17332 17612
rect 17388 17554 17444 17566
rect 17388 17502 17390 17554
rect 17442 17502 17444 17554
rect 17388 17108 17444 17502
rect 17388 17042 17444 17052
rect 17276 16818 17332 16828
rect 17388 16436 17444 16446
rect 17276 16212 17332 16222
rect 17276 16098 17332 16156
rect 17276 16046 17278 16098
rect 17330 16046 17332 16098
rect 17276 16034 17332 16046
rect 17164 15810 17220 15820
rect 17276 15876 17332 15886
rect 17388 15876 17444 16380
rect 17276 15874 17444 15876
rect 17276 15822 17278 15874
rect 17330 15822 17444 15874
rect 17276 15820 17444 15822
rect 17276 15810 17332 15820
rect 17052 15596 17220 15652
rect 16940 15484 17108 15540
rect 16716 15314 16772 15484
rect 16716 15262 16718 15314
rect 16770 15262 16772 15314
rect 16716 15250 16772 15262
rect 16828 15316 16884 15326
rect 16828 14754 16884 15260
rect 16828 14702 16830 14754
rect 16882 14702 16884 14754
rect 16828 14690 16884 14702
rect 16940 15314 16996 15326
rect 16940 15262 16942 15314
rect 16994 15262 16996 15314
rect 16940 14754 16996 15262
rect 17052 14980 17108 15484
rect 17052 14914 17108 14924
rect 16940 14702 16942 14754
rect 16994 14702 16996 14754
rect 16940 14690 16996 14702
rect 17052 14644 17108 14654
rect 16716 14532 16772 14542
rect 16716 14438 16772 14476
rect 16604 13906 16660 13916
rect 16828 14420 16884 14430
rect 16716 13748 16772 13758
rect 16828 13748 16884 14364
rect 16716 13746 16884 13748
rect 16716 13694 16718 13746
rect 16770 13694 16884 13746
rect 16716 13692 16884 13694
rect 16716 13682 16772 13692
rect 16828 12738 16884 12750
rect 16828 12686 16830 12738
rect 16882 12686 16884 12738
rect 16492 12180 16548 12190
rect 16828 12180 16884 12686
rect 16940 12180 16996 12190
rect 16828 12178 16996 12180
rect 16828 12126 16942 12178
rect 16994 12126 16996 12178
rect 16828 12124 16996 12126
rect 17052 12180 17108 14588
rect 17164 14084 17220 15596
rect 17500 15092 17556 15102
rect 17164 14018 17220 14028
rect 17276 14980 17332 14990
rect 17164 12740 17220 12750
rect 17164 12646 17220 12684
rect 17164 12180 17220 12190
rect 17052 12178 17220 12180
rect 17052 12126 17166 12178
rect 17218 12126 17220 12178
rect 17052 12124 17220 12126
rect 16492 12086 16548 12124
rect 16940 12114 16996 12124
rect 16380 11554 16436 11564
rect 17052 11956 17108 11966
rect 15708 9774 15710 9826
rect 15762 9774 15764 9826
rect 15708 9762 15764 9774
rect 15820 10668 15988 10724
rect 16716 11506 16772 11518
rect 16716 11454 16718 11506
rect 16770 11454 16772 11506
rect 15596 9650 15652 9660
rect 15484 9604 15540 9614
rect 15484 9510 15540 9548
rect 15708 9604 15764 9614
rect 15372 8820 15428 8830
rect 15372 8726 15428 8764
rect 15596 8372 15652 8382
rect 15596 8278 15652 8316
rect 15708 8370 15764 9548
rect 15708 8318 15710 8370
rect 15762 8318 15764 8370
rect 15260 8194 15316 8204
rect 15372 8258 15428 8270
rect 15372 8206 15374 8258
rect 15426 8206 15428 8258
rect 15036 8036 15092 8046
rect 15036 7942 15092 7980
rect 15372 8036 15428 8206
rect 15372 7970 15428 7980
rect 15708 7812 15764 8318
rect 15484 7756 15764 7812
rect 15484 7476 15540 7756
rect 15484 7410 15540 7420
rect 14924 7298 14980 7308
rect 15596 7364 15652 7374
rect 15596 7270 15652 7308
rect 15708 7252 15764 7262
rect 15708 7158 15764 7196
rect 15820 6132 15876 10668
rect 16604 10612 16660 10622
rect 15932 10610 16660 10612
rect 15932 10558 16606 10610
rect 16658 10558 16660 10610
rect 15932 10556 16660 10558
rect 15932 7474 15988 10556
rect 16604 10546 16660 10556
rect 16268 10386 16324 10398
rect 16268 10334 16270 10386
rect 16322 10334 16324 10386
rect 16044 10164 16100 10174
rect 16044 10050 16100 10108
rect 16268 10164 16324 10334
rect 16268 10098 16324 10108
rect 16044 9998 16046 10050
rect 16098 9998 16100 10050
rect 16044 9986 16100 9998
rect 16492 10052 16548 10062
rect 16156 9826 16212 9838
rect 16156 9774 16158 9826
rect 16210 9774 16212 9826
rect 15932 7422 15934 7474
rect 15986 7422 15988 7474
rect 15932 7410 15988 7422
rect 16044 9716 16100 9726
rect 14700 5854 14702 5906
rect 14754 5854 14756 5906
rect 14700 5842 14756 5854
rect 15708 6076 15876 6132
rect 15260 5796 15316 5806
rect 14924 5794 15316 5796
rect 14924 5742 15262 5794
rect 15314 5742 15316 5794
rect 14924 5740 15316 5742
rect 14812 5684 14868 5694
rect 14812 5590 14868 5628
rect 14476 5282 14532 5292
rect 14924 5346 14980 5740
rect 15260 5730 15316 5740
rect 14924 5294 14926 5346
rect 14978 5294 14980 5346
rect 14924 5282 14980 5294
rect 15372 5684 15428 5694
rect 15372 5346 15428 5628
rect 15372 5294 15374 5346
rect 15426 5294 15428 5346
rect 15372 5282 15428 5294
rect 13356 5070 13358 5122
rect 13410 5070 13412 5122
rect 13356 5058 13412 5070
rect 15708 5124 15764 6076
rect 16044 5906 16100 9660
rect 16156 9492 16212 9774
rect 16156 9426 16212 9436
rect 16492 9266 16548 9996
rect 16604 9826 16660 9838
rect 16604 9774 16606 9826
rect 16658 9774 16660 9826
rect 16604 9604 16660 9774
rect 16604 9538 16660 9548
rect 16492 9214 16494 9266
rect 16546 9214 16548 9266
rect 16492 9202 16548 9214
rect 16716 8260 16772 11454
rect 17052 11506 17108 11900
rect 17052 11454 17054 11506
rect 17106 11454 17108 11506
rect 17052 11442 17108 11454
rect 17164 11508 17220 12124
rect 17164 11442 17220 11452
rect 16828 11284 16884 11294
rect 16828 10276 16884 11228
rect 17276 10836 17332 14924
rect 17388 13972 17444 13982
rect 17388 13878 17444 13916
rect 17276 10770 17332 10780
rect 17388 12964 17444 12974
rect 17388 10612 17444 12908
rect 17500 12402 17556 15036
rect 17612 13748 17668 18060
rect 17836 17556 17892 17566
rect 17724 17554 17892 17556
rect 17724 17502 17838 17554
rect 17890 17502 17892 17554
rect 17724 17500 17892 17502
rect 17724 16882 17780 17500
rect 17836 17490 17892 17500
rect 18060 17444 18116 21308
rect 18284 21298 18340 21308
rect 18172 19796 18228 19806
rect 18172 19794 18340 19796
rect 18172 19742 18174 19794
rect 18226 19742 18340 19794
rect 18172 19740 18340 19742
rect 18172 19730 18228 19740
rect 18172 19234 18228 19246
rect 18172 19182 18174 19234
rect 18226 19182 18228 19234
rect 18172 18676 18228 19182
rect 18172 18610 18228 18620
rect 18060 17378 18116 17388
rect 18284 18340 18340 19740
rect 18284 17666 18340 18284
rect 18284 17614 18286 17666
rect 18338 17614 18340 17666
rect 18284 17444 18340 17614
rect 18284 17378 18340 17388
rect 18284 17108 18340 17118
rect 18284 17014 18340 17052
rect 17724 16830 17726 16882
rect 17778 16830 17780 16882
rect 17724 15652 17780 16830
rect 17948 16436 18004 16446
rect 17948 16322 18004 16380
rect 17948 16270 17950 16322
rect 18002 16270 18004 16322
rect 17948 16258 18004 16270
rect 17836 16100 17892 16110
rect 17836 16098 18004 16100
rect 17836 16046 17838 16098
rect 17890 16046 18004 16098
rect 17836 16044 18004 16046
rect 17836 16034 17892 16044
rect 17724 15314 17780 15596
rect 17724 15262 17726 15314
rect 17778 15262 17780 15314
rect 17724 14642 17780 15262
rect 17724 14590 17726 14642
rect 17778 14590 17780 14642
rect 17724 14578 17780 14590
rect 17836 15204 17892 15214
rect 17724 13748 17780 13758
rect 17612 13746 17780 13748
rect 17612 13694 17726 13746
rect 17778 13694 17780 13746
rect 17612 13692 17780 13694
rect 17724 12740 17780 13692
rect 17836 13076 17892 15148
rect 17948 14308 18004 16044
rect 18172 16098 18228 16110
rect 18172 16046 18174 16098
rect 18226 16046 18228 16098
rect 18172 15876 18228 16046
rect 18284 16100 18340 16110
rect 18284 16006 18340 16044
rect 18396 15876 18452 22092
rect 18508 21474 18564 21486
rect 18508 21422 18510 21474
rect 18562 21422 18564 21474
rect 18508 21252 18564 21422
rect 18508 21186 18564 21196
rect 18732 21028 18788 23886
rect 18956 23940 19012 23950
rect 18956 23846 19012 23884
rect 19292 23548 19348 29932
rect 19740 29204 19796 29214
rect 19516 29202 19796 29204
rect 19516 29150 19742 29202
rect 19794 29150 19796 29202
rect 19516 29148 19796 29150
rect 19404 28530 19460 28542
rect 19404 28478 19406 28530
rect 19458 28478 19460 28530
rect 19404 27074 19460 28478
rect 19404 27022 19406 27074
rect 19458 27022 19460 27074
rect 19404 23940 19460 27022
rect 19404 23874 19460 23884
rect 19516 23548 19572 29148
rect 19740 29138 19796 29148
rect 20412 28756 20468 28766
rect 20412 28754 20692 28756
rect 20412 28702 20414 28754
rect 20466 28702 20692 28754
rect 20412 28700 20692 28702
rect 20412 28690 20468 28700
rect 19852 28642 19908 28654
rect 19852 28590 19854 28642
rect 19906 28590 19908 28642
rect 19740 27634 19796 27646
rect 19740 27582 19742 27634
rect 19794 27582 19796 27634
rect 19740 25620 19796 27582
rect 19852 26516 19908 28590
rect 20300 28642 20356 28654
rect 20300 28590 20302 28642
rect 20354 28590 20356 28642
rect 20300 26908 20356 28590
rect 20636 27858 20692 28700
rect 20636 27806 20638 27858
rect 20690 27806 20692 27858
rect 20636 27794 20692 27806
rect 20188 26852 20356 26908
rect 20524 27074 20580 27086
rect 20524 27022 20526 27074
rect 20578 27022 20580 27074
rect 19964 26516 20020 26526
rect 19852 26514 20020 26516
rect 19852 26462 19966 26514
rect 20018 26462 20020 26514
rect 19852 26460 20020 26462
rect 19964 26450 20020 26460
rect 19180 23492 19348 23548
rect 19404 23492 19572 23548
rect 19628 25564 19796 25620
rect 20076 25618 20132 25630
rect 20076 25566 20078 25618
rect 20130 25566 20132 25618
rect 19068 22372 19124 22382
rect 19068 21924 19124 22316
rect 19068 21586 19124 21868
rect 19068 21534 19070 21586
rect 19122 21534 19124 21586
rect 19068 21522 19124 21534
rect 18508 20972 18788 21028
rect 18844 21474 18900 21486
rect 18844 21422 18846 21474
rect 18898 21422 18900 21474
rect 18844 21028 18900 21422
rect 18508 19012 18564 20972
rect 18844 20962 18900 20972
rect 19068 21252 19124 21262
rect 19068 20808 19124 21196
rect 19068 20756 19070 20808
rect 19122 20756 19124 20808
rect 19068 20744 19124 20756
rect 18732 20690 18788 20702
rect 18732 20638 18734 20690
rect 18786 20638 18788 20690
rect 18732 20020 18788 20638
rect 18732 19954 18788 19964
rect 18620 19908 18676 19918
rect 18620 19814 18676 19852
rect 18732 19794 18788 19806
rect 18732 19742 18734 19794
rect 18786 19742 18788 19794
rect 18508 18946 18564 18956
rect 18620 19572 18676 19582
rect 18508 18450 18564 18462
rect 18508 18398 18510 18450
rect 18562 18398 18564 18450
rect 18508 17668 18564 18398
rect 18508 17602 18564 17612
rect 18620 17666 18676 19516
rect 18620 17614 18622 17666
rect 18674 17614 18676 17666
rect 18508 17108 18564 17118
rect 18508 17014 18564 17052
rect 18620 16884 18676 17614
rect 18732 17108 18788 19742
rect 18844 19794 18900 19806
rect 18844 19742 18846 19794
rect 18898 19742 18900 19794
rect 18844 19684 18900 19742
rect 18844 19618 18900 19628
rect 19180 19012 19236 23492
rect 19292 22258 19348 22270
rect 19292 22206 19294 22258
rect 19346 22206 19348 22258
rect 19292 22148 19348 22206
rect 19292 22082 19348 22092
rect 19292 21588 19348 21598
rect 19292 21494 19348 21532
rect 19292 21140 19348 21150
rect 19292 19460 19348 21084
rect 19404 21028 19460 23492
rect 19628 23044 19684 25564
rect 19740 25396 19796 25406
rect 19740 25302 19796 25340
rect 20076 24052 20132 25566
rect 20188 25284 20244 26796
rect 20524 25956 20580 27022
rect 20748 26908 20804 30828
rect 20860 30434 20916 31724
rect 20972 31686 21028 31724
rect 20972 31108 21028 31118
rect 20972 30994 21028 31052
rect 20972 30942 20974 30994
rect 21026 30942 21028 30994
rect 20972 30930 21028 30942
rect 20860 30382 20862 30434
rect 20914 30382 20916 30434
rect 20860 30370 20916 30382
rect 21084 29092 21140 40012
rect 21308 34914 21364 34926
rect 21308 34862 21310 34914
rect 21362 34862 21364 34914
rect 21308 34132 21364 34862
rect 21308 34066 21364 34076
rect 21532 33124 21588 54350
rect 21756 52276 21812 56030
rect 22428 55300 22484 55310
rect 22428 55206 22484 55244
rect 22540 54738 22596 56140
rect 22988 55522 23044 57372
rect 23520 57344 23632 57456
rect 24864 57344 24976 57456
rect 25564 57372 25956 57428
rect 23548 56308 23604 57344
rect 24332 56644 24388 56654
rect 23804 56476 24068 56486
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 23804 56410 24068 56420
rect 23548 56242 23604 56252
rect 22988 55470 22990 55522
rect 23042 55470 23044 55522
rect 22988 55458 23044 55470
rect 23884 55970 23940 55982
rect 23884 55918 23886 55970
rect 23938 55918 23940 55970
rect 23884 55468 23940 55918
rect 22540 54686 22542 54738
rect 22594 54686 22596 54738
rect 22540 54674 22596 54686
rect 23548 55412 23604 55422
rect 21980 54068 22036 54078
rect 21980 53618 22036 54012
rect 21980 53566 21982 53618
rect 22034 53566 22036 53618
rect 21980 53554 22036 53566
rect 22428 53730 22484 53742
rect 22428 53678 22430 53730
rect 22482 53678 22484 53730
rect 21980 52276 22036 52286
rect 21756 52274 22036 52276
rect 21756 52222 21982 52274
rect 22034 52222 22036 52274
rect 21756 52220 22036 52222
rect 21980 52210 22036 52220
rect 22428 50820 22484 53678
rect 22764 53732 22820 53742
rect 22764 53638 22820 53676
rect 23548 53730 23604 55356
rect 23660 55412 23940 55468
rect 24220 55972 24276 55982
rect 23660 54068 23716 55412
rect 23804 54908 24068 54918
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 23804 54842 24068 54852
rect 23772 54740 23828 54750
rect 23772 54646 23828 54684
rect 24108 54516 24164 54526
rect 24108 54422 24164 54460
rect 23660 54002 23716 54012
rect 23548 53678 23550 53730
rect 23602 53678 23604 53730
rect 23548 53666 23604 53678
rect 23804 53340 24068 53350
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 23804 53274 24068 53284
rect 24220 53060 24276 55916
rect 23548 53004 24276 53060
rect 23212 52946 23268 52958
rect 23212 52894 23214 52946
rect 23266 52894 23268 52946
rect 22764 52164 22820 52174
rect 22764 52070 22820 52108
rect 22428 50754 22484 50764
rect 23212 43708 23268 52894
rect 23548 50482 23604 53004
rect 24332 52948 24388 56588
rect 24444 56308 24500 56318
rect 24444 56214 24500 56252
rect 24892 56308 24948 57344
rect 24892 56242 24948 56252
rect 25004 57204 25060 57214
rect 24464 55692 24728 55702
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24464 55626 24728 55636
rect 24892 55300 24948 55310
rect 24892 55206 24948 55244
rect 24892 54514 24948 54526
rect 24892 54462 24894 54514
rect 24946 54462 24948 54514
rect 24464 54124 24728 54134
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24464 54058 24728 54068
rect 24892 53956 24948 54462
rect 24892 53890 24948 53900
rect 24668 53730 24724 53742
rect 24668 53678 24670 53730
rect 24722 53678 24724 53730
rect 24668 53620 24724 53678
rect 24668 53554 24724 53564
rect 23772 52892 24388 52948
rect 23660 52724 23716 52734
rect 23660 52630 23716 52668
rect 23772 52050 23828 52892
rect 24668 52836 24724 52846
rect 24668 52742 24724 52780
rect 25004 52724 25060 57148
rect 25452 55972 25508 55982
rect 25452 55878 25508 55916
rect 25004 52658 25060 52668
rect 25340 55300 25396 55310
rect 24464 52556 24728 52566
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24464 52490 24728 52500
rect 24892 52164 24948 52174
rect 24892 52070 24948 52108
rect 23772 51998 23774 52050
rect 23826 51998 23828 52050
rect 23772 51986 23828 51998
rect 23804 51772 24068 51782
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 23804 51706 24068 51716
rect 24668 51268 24724 51278
rect 24668 51174 24724 51212
rect 24464 50988 24728 50998
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24464 50922 24728 50932
rect 23884 50596 23940 50606
rect 23884 50502 23940 50540
rect 24668 50594 24724 50606
rect 24668 50542 24670 50594
rect 24722 50542 24724 50594
rect 23548 50430 23550 50482
rect 23602 50430 23604 50482
rect 23548 50418 23604 50430
rect 24668 50484 24724 50542
rect 24668 50418 24724 50428
rect 23804 50204 24068 50214
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 23804 50138 24068 50148
rect 24668 49700 24724 49710
rect 24668 49606 24724 49644
rect 24464 49420 24728 49430
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24464 49354 24728 49364
rect 24668 49028 24724 49038
rect 24668 48934 24724 48972
rect 23804 48636 24068 48646
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 23804 48570 24068 48580
rect 24464 47852 24728 47862
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24464 47786 24728 47796
rect 24668 47460 24724 47470
rect 24668 47366 24724 47404
rect 23804 47068 24068 47078
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 23804 47002 24068 47012
rect 24668 46564 24724 46574
rect 24668 46470 24724 46508
rect 24464 46284 24728 46294
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24464 46218 24728 46228
rect 24668 45892 24724 45902
rect 24668 45798 24724 45836
rect 23804 45500 24068 45510
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 23804 45434 24068 45444
rect 24464 44716 24728 44726
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24464 44650 24728 44660
rect 24668 44324 24724 44334
rect 24668 44230 24724 44268
rect 23804 43932 24068 43942
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 23804 43866 24068 43876
rect 23212 43652 23492 43708
rect 23324 42868 23380 42878
rect 22316 39620 22372 39630
rect 22316 38668 22372 39564
rect 22204 38612 22372 38668
rect 21532 33058 21588 33068
rect 21868 34580 21924 34590
rect 21196 32564 21252 32574
rect 21196 32562 21700 32564
rect 21196 32510 21198 32562
rect 21250 32510 21700 32562
rect 21196 32508 21700 32510
rect 21196 32498 21252 32508
rect 21532 32340 21588 32350
rect 21308 32338 21588 32340
rect 21308 32286 21534 32338
rect 21586 32286 21588 32338
rect 21308 32284 21588 32286
rect 21196 32004 21252 32014
rect 21308 32004 21364 32284
rect 21532 32274 21588 32284
rect 21196 32002 21364 32004
rect 21196 31950 21198 32002
rect 21250 31950 21364 32002
rect 21196 31948 21364 31950
rect 21420 32004 21476 32014
rect 21196 31938 21252 31948
rect 21420 31780 21476 31948
rect 20972 29036 21140 29092
rect 21196 31724 21476 31780
rect 21532 31780 21588 31790
rect 20748 26852 20916 26908
rect 20524 25890 20580 25900
rect 20748 26290 20804 26302
rect 20748 26238 20750 26290
rect 20802 26238 20804 26290
rect 20748 25732 20804 26238
rect 20188 25218 20244 25228
rect 20524 25676 20804 25732
rect 20524 25396 20580 25676
rect 20076 23996 20244 24052
rect 19852 23940 19908 23950
rect 19852 23938 20132 23940
rect 19852 23886 19854 23938
rect 19906 23886 20132 23938
rect 19852 23884 20132 23886
rect 19852 23874 19908 23884
rect 19964 23156 20020 23166
rect 19516 23042 19684 23044
rect 19516 22990 19630 23042
rect 19682 22990 19684 23042
rect 19516 22988 19684 22990
rect 19516 21588 19572 22988
rect 19628 22978 19684 22988
rect 19740 23154 20020 23156
rect 19740 23102 19966 23154
rect 20018 23102 20020 23154
rect 19740 23100 20020 23102
rect 19628 22372 19684 22382
rect 19628 22278 19684 22316
rect 19740 22036 19796 23100
rect 19964 23090 20020 23100
rect 20076 23156 20132 23884
rect 20188 23492 20244 23996
rect 20524 23938 20580 25340
rect 20748 25396 20804 25406
rect 20636 24836 20692 24846
rect 20748 24836 20804 25340
rect 20636 24834 20804 24836
rect 20636 24782 20638 24834
rect 20690 24782 20804 24834
rect 20636 24780 20804 24782
rect 20636 24770 20692 24780
rect 20524 23886 20526 23938
rect 20578 23886 20580 23938
rect 20524 23874 20580 23886
rect 20188 23426 20244 23436
rect 20860 23380 20916 26852
rect 20972 24948 21028 29036
rect 21084 28642 21140 28654
rect 21084 28590 21086 28642
rect 21138 28590 21140 28642
rect 21084 26908 21140 28590
rect 21196 27970 21252 31724
rect 21196 27918 21198 27970
rect 21250 27918 21252 27970
rect 21196 27906 21252 27918
rect 21308 31556 21364 31566
rect 21308 27188 21364 31500
rect 21532 30994 21588 31724
rect 21532 30942 21534 30994
rect 21586 30942 21588 30994
rect 21420 30212 21476 30222
rect 21420 30118 21476 30156
rect 21308 27122 21364 27132
rect 21420 28642 21476 28654
rect 21420 28590 21422 28642
rect 21474 28590 21476 28642
rect 21084 26852 21252 26908
rect 21084 25956 21140 25966
rect 21084 25060 21140 25900
rect 21196 25732 21252 26852
rect 21308 26068 21364 26078
rect 21308 25974 21364 26012
rect 21308 25732 21364 25742
rect 21196 25730 21364 25732
rect 21196 25678 21310 25730
rect 21362 25678 21364 25730
rect 21196 25676 21364 25678
rect 21308 25666 21364 25676
rect 21420 25508 21476 28590
rect 21532 27524 21588 30942
rect 21644 30882 21700 32508
rect 21644 30830 21646 30882
rect 21698 30830 21700 30882
rect 21644 30818 21700 30830
rect 21756 31778 21812 31790
rect 21756 31726 21758 31778
rect 21810 31726 21812 31778
rect 21644 30324 21700 30334
rect 21644 28642 21700 30268
rect 21756 30212 21812 31726
rect 21756 30146 21812 30156
rect 21868 30322 21924 34524
rect 22092 32676 22148 32686
rect 22092 32582 22148 32620
rect 22092 30996 22148 31006
rect 22092 30902 22148 30940
rect 21868 30270 21870 30322
rect 21922 30270 21924 30322
rect 21644 28590 21646 28642
rect 21698 28590 21700 28642
rect 21644 28578 21700 28590
rect 21532 27458 21588 27468
rect 21308 25452 21476 25508
rect 21532 27188 21588 27198
rect 21308 25396 21364 25452
rect 21308 25330 21364 25340
rect 21420 25284 21476 25294
rect 21084 25004 21364 25060
rect 20972 24892 21252 24948
rect 21084 24722 21140 24734
rect 21084 24670 21086 24722
rect 21138 24670 21140 24722
rect 21084 24164 21140 24670
rect 21084 24098 21140 24108
rect 20972 24052 21028 24062
rect 20972 23958 21028 23996
rect 20860 23324 21028 23380
rect 20076 23090 20132 23100
rect 19740 21970 19796 21980
rect 19852 22930 19908 22942
rect 20076 22932 20132 22942
rect 19852 22878 19854 22930
rect 19906 22878 19908 22930
rect 19852 22148 19908 22878
rect 19852 21812 19908 22092
rect 19516 21522 19572 21532
rect 19628 21756 19908 21812
rect 19964 22930 20132 22932
rect 19964 22878 20078 22930
rect 20130 22878 20132 22930
rect 19964 22876 20132 22878
rect 19628 21586 19684 21756
rect 19964 21700 20020 22876
rect 20076 22866 20132 22876
rect 20300 22482 20356 22494
rect 20300 22430 20302 22482
rect 20354 22430 20356 22482
rect 20076 22370 20132 22382
rect 20076 22318 20078 22370
rect 20130 22318 20132 22370
rect 20076 22260 20132 22318
rect 20076 22194 20132 22204
rect 20188 22372 20244 22382
rect 19628 21534 19630 21586
rect 19682 21534 19684 21586
rect 19628 21522 19684 21534
rect 19740 21644 20020 21700
rect 19628 21364 19684 21374
rect 19628 21270 19684 21308
rect 19404 20244 19460 20972
rect 19516 21140 19572 21150
rect 19516 20802 19572 21084
rect 19740 21026 19796 21644
rect 20076 21474 20132 21486
rect 20076 21422 20078 21474
rect 20130 21422 20132 21474
rect 19964 21362 20020 21374
rect 19964 21310 19966 21362
rect 20018 21310 20020 21362
rect 19964 21140 20020 21310
rect 19964 21074 20020 21084
rect 19740 20974 19742 21026
rect 19794 20974 19796 21026
rect 19740 20962 19796 20974
rect 20076 21028 20132 21422
rect 20076 20962 20132 20972
rect 19516 20750 19518 20802
rect 19570 20750 19572 20802
rect 19516 20738 19572 20750
rect 20188 20914 20244 22316
rect 20188 20862 20190 20914
rect 20242 20862 20244 20914
rect 19404 20178 19460 20188
rect 19740 20244 19796 20254
rect 19740 20018 19796 20188
rect 19964 20244 20020 20254
rect 19964 20130 20020 20188
rect 19964 20078 19966 20130
rect 20018 20078 20020 20130
rect 19964 20066 20020 20078
rect 20188 20132 20244 20862
rect 20300 20244 20356 22430
rect 20748 22370 20804 22382
rect 20748 22318 20750 22370
rect 20802 22318 20804 22370
rect 20636 21586 20692 21598
rect 20636 21534 20638 21586
rect 20690 21534 20692 21586
rect 20636 21364 20692 21534
rect 20636 21298 20692 21308
rect 20748 21252 20804 22318
rect 20300 20188 20692 20244
rect 20188 20066 20244 20076
rect 20636 20130 20692 20188
rect 20636 20078 20638 20130
rect 20690 20078 20692 20130
rect 20636 20066 20692 20078
rect 19740 19966 19742 20018
rect 19794 19966 19796 20018
rect 19740 19908 19796 19966
rect 19740 19842 19796 19852
rect 19852 20020 19908 20030
rect 19516 19684 19572 19694
rect 19292 19404 19460 19460
rect 19180 18946 19236 18956
rect 19292 19234 19348 19246
rect 19292 19182 19294 19234
rect 19346 19182 19348 19234
rect 18844 18900 18900 18910
rect 18844 18338 18900 18844
rect 19292 18900 19348 19182
rect 19292 18834 19348 18844
rect 18844 18286 18846 18338
rect 18898 18286 18900 18338
rect 18844 18228 18900 18286
rect 18844 18162 18900 18172
rect 19068 18450 19124 18462
rect 19068 18398 19070 18450
rect 19122 18398 19124 18450
rect 19068 18116 19124 18398
rect 19068 18050 19124 18060
rect 19292 18228 19348 18238
rect 18844 17780 18900 17790
rect 18844 17686 18900 17724
rect 19292 17668 19348 18172
rect 19292 17574 19348 17612
rect 19404 17220 19460 19404
rect 19516 18226 19572 19628
rect 19852 19346 19908 19964
rect 20076 19908 20132 19918
rect 20076 19906 20356 19908
rect 20076 19854 20078 19906
rect 20130 19854 20356 19906
rect 20076 19852 20356 19854
rect 20076 19842 20132 19852
rect 20300 19458 20356 19852
rect 20300 19406 20302 19458
rect 20354 19406 20356 19458
rect 20300 19394 20356 19406
rect 20412 19572 20468 19582
rect 19852 19294 19854 19346
rect 19906 19294 19908 19346
rect 19852 19236 19908 19294
rect 19852 19170 19908 19180
rect 20412 19234 20468 19516
rect 20412 19182 20414 19234
rect 20466 19182 20468 19234
rect 20412 19170 20468 19182
rect 20748 19236 20804 21196
rect 20860 21586 20916 21598
rect 20860 21534 20862 21586
rect 20914 21534 20916 21586
rect 20860 20244 20916 21534
rect 20972 21364 21028 23324
rect 21084 21588 21140 21598
rect 21084 21494 21140 21532
rect 21196 21364 21252 24892
rect 20972 21308 21140 21364
rect 20972 20802 21028 20814
rect 20972 20750 20974 20802
rect 21026 20750 21028 20802
rect 20972 20468 21028 20750
rect 20972 20402 21028 20412
rect 20860 20178 20916 20188
rect 20972 20132 21028 20142
rect 20972 20038 21028 20076
rect 20860 19908 20916 19918
rect 20860 19814 20916 19852
rect 21084 19908 21140 21308
rect 21196 21298 21252 21308
rect 21308 22370 21364 25004
rect 21420 24722 21476 25228
rect 21420 24670 21422 24722
rect 21474 24670 21476 24722
rect 21420 24658 21476 24670
rect 21532 24164 21588 27132
rect 21868 26068 21924 30270
rect 22204 28756 22260 38612
rect 22428 31778 22484 31790
rect 22428 31726 22430 31778
rect 22482 31726 22484 31778
rect 22428 30996 22484 31726
rect 23212 31778 23268 31790
rect 23212 31726 23214 31778
rect 23266 31726 23268 31778
rect 23212 31444 23268 31726
rect 23212 31378 23268 31388
rect 22652 30996 22708 31006
rect 22428 30994 22708 30996
rect 22428 30942 22654 30994
rect 22706 30942 22708 30994
rect 22428 30940 22708 30942
rect 22092 28700 22260 28756
rect 22428 30772 22484 30782
rect 22092 26964 22148 28700
rect 22428 28642 22484 30716
rect 22428 28590 22430 28642
rect 22482 28590 22484 28642
rect 22428 28420 22484 28590
rect 22092 26898 22148 26908
rect 22204 28364 22484 28420
rect 21756 25508 21812 25518
rect 21644 25506 21812 25508
rect 21644 25454 21758 25506
rect 21810 25454 21812 25506
rect 21644 25452 21812 25454
rect 21644 24610 21700 25452
rect 21756 25442 21812 25452
rect 21644 24558 21646 24610
rect 21698 24558 21700 24610
rect 21644 24546 21700 24558
rect 21756 25284 21812 25294
rect 21532 24108 21700 24164
rect 21308 22318 21310 22370
rect 21362 22318 21364 22370
rect 21084 19842 21140 19852
rect 21196 20468 21252 20478
rect 20860 19236 20916 19246
rect 20748 19234 20916 19236
rect 20748 19182 20862 19234
rect 20914 19182 20916 19234
rect 20748 19180 20916 19182
rect 20860 19170 20916 19180
rect 20076 18900 20132 18910
rect 19516 18174 19518 18226
rect 19570 18174 19572 18226
rect 19516 17892 19572 18174
rect 19516 17826 19572 17836
rect 19628 18226 19684 18238
rect 19628 18174 19630 18226
rect 19682 18174 19684 18226
rect 19628 17220 19684 18174
rect 19740 18228 19796 18238
rect 19740 18226 19908 18228
rect 19740 18174 19742 18226
rect 19794 18174 19908 18226
rect 19740 18172 19908 18174
rect 19740 18162 19796 18172
rect 19404 17154 19460 17164
rect 19516 17164 19684 17220
rect 18732 17042 18788 17052
rect 18172 15810 18228 15820
rect 18284 15820 18452 15876
rect 18508 16828 18676 16884
rect 18732 16882 18788 16894
rect 18732 16830 18734 16882
rect 18786 16830 18788 16882
rect 18284 15148 18340 15820
rect 18508 15764 18564 16828
rect 18620 16660 18676 16670
rect 18620 16098 18676 16604
rect 18732 16548 18788 16830
rect 19180 16884 19236 16894
rect 19516 16884 19572 17164
rect 19180 16882 19572 16884
rect 19180 16830 19182 16882
rect 19234 16830 19572 16882
rect 19180 16828 19572 16830
rect 19628 16994 19684 17006
rect 19628 16942 19630 16994
rect 19682 16942 19684 16994
rect 19180 16818 19236 16828
rect 18732 16482 18788 16492
rect 18956 16770 19012 16782
rect 18956 16718 18958 16770
rect 19010 16718 19012 16770
rect 18956 16436 19012 16718
rect 19068 16770 19124 16782
rect 19068 16718 19070 16770
rect 19122 16718 19124 16770
rect 19068 16660 19124 16718
rect 19068 16604 19236 16660
rect 18956 16370 19012 16380
rect 18620 16046 18622 16098
rect 18674 16046 18676 16098
rect 18620 16034 18676 16046
rect 18732 16100 18788 16110
rect 18956 16100 19012 16110
rect 18788 16098 19012 16100
rect 18788 16046 18958 16098
rect 19010 16046 19012 16098
rect 18788 16044 19012 16046
rect 18732 16034 18788 16044
rect 18396 15316 18452 15326
rect 18396 15222 18452 15260
rect 18172 15092 18340 15148
rect 18396 15092 18452 15102
rect 17948 14242 18004 14252
rect 18060 14532 18116 14542
rect 17836 12982 17892 13020
rect 17948 12964 18004 12974
rect 18060 12964 18116 14476
rect 17948 12962 18116 12964
rect 17948 12910 17950 12962
rect 18002 12910 18116 12962
rect 17948 12908 18116 12910
rect 17948 12898 18004 12908
rect 18060 12852 18116 12908
rect 18060 12786 18116 12796
rect 17724 12674 17780 12684
rect 17500 12350 17502 12402
rect 17554 12350 17556 12402
rect 17500 12338 17556 12350
rect 17612 12292 17668 12302
rect 17612 12178 17668 12236
rect 18060 12180 18116 12190
rect 17612 12126 17614 12178
rect 17666 12126 17668 12178
rect 17612 12114 17668 12126
rect 18004 12178 18116 12180
rect 18004 12126 18062 12178
rect 18114 12126 18116 12178
rect 18004 12114 18116 12126
rect 18004 12068 18060 12114
rect 17724 12012 18060 12068
rect 17724 11954 17780 12012
rect 17724 11902 17726 11954
rect 17778 11902 17780 11954
rect 17724 11890 17780 11902
rect 17836 11844 17892 11854
rect 18060 11844 18116 11854
rect 17836 11732 18004 11788
rect 17724 11284 17780 11294
rect 17612 11282 17780 11284
rect 17612 11230 17726 11282
rect 17778 11230 17780 11282
rect 17612 11228 17780 11230
rect 17500 10612 17556 10622
rect 17388 10610 17556 10612
rect 17388 10558 17502 10610
rect 17554 10558 17556 10610
rect 17388 10556 17556 10558
rect 17500 10546 17556 10556
rect 16940 10388 16996 10398
rect 16940 10386 17108 10388
rect 16940 10334 16942 10386
rect 16994 10334 17108 10386
rect 16940 10332 17108 10334
rect 16940 10322 16996 10332
rect 16828 10210 16884 10220
rect 17052 10052 17108 10332
rect 17164 10386 17220 10398
rect 17164 10334 17166 10386
rect 17218 10334 17220 10386
rect 17164 10164 17220 10334
rect 17276 10388 17332 10398
rect 17276 10386 17556 10388
rect 17276 10334 17278 10386
rect 17330 10334 17556 10386
rect 17276 10332 17556 10334
rect 17276 10322 17332 10332
rect 17164 10108 17332 10164
rect 17276 10052 17332 10108
rect 17052 9996 17220 10052
rect 16940 9940 16996 9950
rect 16940 9268 16996 9884
rect 17164 9938 17220 9996
rect 17332 9996 17444 10052
rect 17276 9986 17332 9996
rect 17164 9886 17166 9938
rect 17218 9886 17220 9938
rect 17164 9874 17220 9886
rect 17052 9828 17108 9838
rect 17052 9734 17108 9772
rect 17276 9828 17332 9838
rect 17276 9734 17332 9772
rect 17052 9268 17108 9278
rect 16940 9266 17108 9268
rect 16940 9214 17054 9266
rect 17106 9214 17108 9266
rect 16940 9212 17108 9214
rect 17052 9202 17108 9212
rect 17388 9156 17444 9996
rect 17276 9100 17444 9156
rect 16492 8204 16772 8260
rect 16940 8260 16996 8270
rect 16156 8036 16212 8046
rect 16156 7942 16212 7980
rect 16156 7476 16212 7486
rect 16156 7382 16212 7420
rect 16380 7474 16436 7486
rect 16380 7422 16382 7474
rect 16434 7422 16436 7474
rect 16380 7364 16436 7422
rect 16380 7298 16436 7308
rect 16492 6580 16548 8204
rect 16940 8166 16996 8204
rect 17276 8258 17332 9100
rect 17500 8372 17556 10332
rect 17612 9940 17668 11228
rect 17724 11218 17780 11228
rect 17724 10724 17780 10734
rect 17724 10630 17780 10668
rect 17836 10498 17892 10510
rect 17836 10446 17838 10498
rect 17890 10446 17892 10498
rect 17612 9380 17668 9884
rect 17724 10276 17780 10286
rect 17724 9828 17780 10220
rect 17836 10052 17892 10446
rect 17836 9986 17892 9996
rect 17948 9940 18004 11732
rect 18060 11394 18116 11788
rect 18060 11342 18062 11394
rect 18114 11342 18116 11394
rect 18060 10164 18116 11342
rect 18060 10098 18116 10108
rect 17948 9884 18116 9940
rect 17724 9762 17780 9772
rect 17948 9716 18004 9726
rect 17612 9314 17668 9324
rect 17836 9714 18004 9716
rect 17836 9662 17950 9714
rect 18002 9662 18004 9714
rect 17836 9660 18004 9662
rect 17836 9492 17892 9660
rect 17948 9650 18004 9660
rect 18060 9492 18116 9884
rect 17836 8484 17892 9436
rect 17836 8418 17892 8428
rect 17948 9436 18116 9492
rect 17612 8372 17668 8382
rect 17500 8370 17668 8372
rect 17500 8318 17614 8370
rect 17666 8318 17668 8370
rect 17500 8316 17668 8318
rect 17612 8306 17668 8316
rect 17276 8206 17278 8258
rect 17330 8206 17332 8258
rect 17276 8194 17332 8206
rect 17388 8258 17444 8270
rect 17388 8206 17390 8258
rect 17442 8206 17444 8258
rect 16716 8036 16772 8046
rect 16716 7942 16772 7980
rect 16604 7812 16660 7822
rect 16604 7698 16660 7756
rect 17052 7812 17108 7822
rect 16604 7646 16606 7698
rect 16658 7646 16660 7698
rect 16604 7634 16660 7646
rect 16716 7700 16772 7710
rect 16716 7606 16772 7644
rect 17052 7586 17108 7756
rect 17388 7700 17444 8206
rect 17388 7634 17444 7644
rect 17500 8146 17556 8158
rect 17500 8094 17502 8146
rect 17554 8094 17556 8146
rect 17052 7534 17054 7586
rect 17106 7534 17108 7586
rect 17052 7522 17108 7534
rect 16492 6514 16548 6524
rect 16940 7476 16996 7486
rect 16044 5854 16046 5906
rect 16098 5854 16100 5906
rect 16044 5842 16100 5854
rect 16940 5906 16996 7420
rect 17388 7476 17444 7486
rect 17388 7382 17444 7420
rect 16940 5854 16942 5906
rect 16994 5854 16996 5906
rect 16940 5842 16996 5854
rect 15932 5348 15988 5358
rect 15932 5234 15988 5292
rect 15932 5182 15934 5234
rect 15986 5182 15988 5234
rect 15932 5170 15988 5182
rect 15708 5058 15764 5068
rect 15484 4900 15540 4910
rect 11788 3332 11956 3388
rect 11452 1036 11620 1092
rect 10108 980 10164 990
rect 10108 112 10164 924
rect 11452 112 11508 1036
rect 11900 980 11956 3332
rect 13244 2100 13300 2110
rect 13244 2006 13300 2044
rect 11900 914 11956 924
rect 12012 1986 12068 1998
rect 12012 1934 12014 1986
rect 12066 1934 12068 1986
rect 12012 644 12068 1934
rect 13804 1988 13860 1998
rect 13804 1894 13860 1932
rect 12012 578 12068 588
rect 12796 1316 12852 1326
rect 12796 112 12852 1260
rect 14140 980 14196 990
rect 14140 112 14196 924
rect 15484 112 15540 4844
rect 17500 4228 17556 8094
rect 17948 5236 18004 9436
rect 18172 9268 18228 15092
rect 18396 14998 18452 15036
rect 18508 14530 18564 15708
rect 18844 15876 18900 15886
rect 18620 15538 18676 15550
rect 18620 15486 18622 15538
rect 18674 15486 18676 15538
rect 18620 14644 18676 15486
rect 18844 15314 18900 15820
rect 18844 15262 18846 15314
rect 18898 15262 18900 15314
rect 18844 15250 18900 15262
rect 18620 14578 18676 14588
rect 18732 14642 18788 14654
rect 18732 14590 18734 14642
rect 18786 14590 18788 14642
rect 18508 14478 18510 14530
rect 18562 14478 18564 14530
rect 18508 14466 18564 14478
rect 18396 14308 18452 14318
rect 18396 13746 18452 14252
rect 18396 13694 18398 13746
rect 18450 13694 18452 13746
rect 18396 13682 18452 13694
rect 18284 13634 18340 13646
rect 18284 13582 18286 13634
rect 18338 13582 18340 13634
rect 18284 13076 18340 13582
rect 18284 13010 18340 13020
rect 18732 13074 18788 14590
rect 18732 13022 18734 13074
rect 18786 13022 18788 13074
rect 18732 13010 18788 13022
rect 18956 13076 19012 16044
rect 19180 15988 19236 16604
rect 19404 16436 19460 16446
rect 19404 16098 19460 16380
rect 19404 16046 19406 16098
rect 19458 16046 19460 16098
rect 19404 16034 19460 16046
rect 19628 16100 19684 16942
rect 19740 16884 19796 16894
rect 19852 16884 19908 18172
rect 19964 17892 20020 17902
rect 19964 17106 20020 17836
rect 19964 17054 19966 17106
rect 20018 17054 20020 17106
rect 19964 17042 20020 17054
rect 20076 17666 20132 18844
rect 20860 18676 20916 18686
rect 20636 18338 20692 18350
rect 20636 18286 20638 18338
rect 20690 18286 20692 18338
rect 20524 18228 20580 18238
rect 20076 17614 20078 17666
rect 20130 17614 20132 17666
rect 19852 16828 20020 16884
rect 19740 16770 19796 16828
rect 19740 16718 19742 16770
rect 19794 16718 19796 16770
rect 19740 16706 19796 16718
rect 19628 16034 19684 16044
rect 19740 16436 19796 16446
rect 19740 16100 19796 16380
rect 19964 16322 20020 16828
rect 19964 16270 19966 16322
rect 20018 16270 20020 16322
rect 19964 16258 20020 16270
rect 19740 16098 19908 16100
rect 19740 16046 19742 16098
rect 19794 16046 19908 16098
rect 19740 16044 19908 16046
rect 19740 16034 19796 16044
rect 19180 15922 19236 15932
rect 19740 15316 19796 15326
rect 19740 15222 19796 15260
rect 19180 15202 19236 15214
rect 19180 15150 19182 15202
rect 19234 15150 19236 15202
rect 19180 14532 19236 15150
rect 19180 14466 19236 14476
rect 19292 14644 19348 14654
rect 19292 14530 19348 14588
rect 19292 14478 19294 14530
rect 19346 14478 19348 14530
rect 19292 14466 19348 14478
rect 19740 14644 19796 14654
rect 19740 14530 19796 14588
rect 19740 14478 19742 14530
rect 19794 14478 19796 14530
rect 19740 14466 19796 14478
rect 19068 14084 19124 14094
rect 19068 13970 19124 14028
rect 19068 13918 19070 13970
rect 19122 13918 19124 13970
rect 19068 13906 19124 13918
rect 19292 13972 19348 13982
rect 19292 13878 19348 13916
rect 19740 13860 19796 13898
rect 19740 13794 19796 13804
rect 19516 13746 19572 13758
rect 19516 13694 19518 13746
rect 19570 13694 19572 13746
rect 19516 13300 19572 13694
rect 19740 13524 19796 13534
rect 19740 13430 19796 13468
rect 19572 13244 19796 13300
rect 19516 13234 19572 13244
rect 19180 13076 19236 13086
rect 18956 13020 19180 13076
rect 19180 12982 19236 13020
rect 18396 12964 18452 12974
rect 18396 12870 18452 12908
rect 19628 12962 19684 12974
rect 19628 12910 19630 12962
rect 19682 12910 19684 12962
rect 19628 12852 19684 12910
rect 19628 12786 19684 12796
rect 18396 12738 18452 12750
rect 18396 12686 18398 12738
rect 18450 12686 18452 12738
rect 18284 12404 18340 12414
rect 18396 12404 18452 12686
rect 18284 12402 18452 12404
rect 18284 12350 18286 12402
rect 18338 12350 18452 12402
rect 18284 12348 18452 12350
rect 18284 12338 18340 12348
rect 19628 12292 19684 12302
rect 18508 12180 18564 12190
rect 18508 12086 18564 12124
rect 18956 12180 19012 12190
rect 19516 12180 19572 12190
rect 18956 12178 19572 12180
rect 18956 12126 18958 12178
rect 19010 12126 19518 12178
rect 19570 12126 19572 12178
rect 18956 12124 19572 12126
rect 18956 12114 19012 12124
rect 19516 12114 19572 12124
rect 19628 12178 19684 12236
rect 19628 12126 19630 12178
rect 19682 12126 19684 12178
rect 19628 12114 19684 12126
rect 19180 12012 19460 12068
rect 18732 11956 18788 11966
rect 18620 11954 18788 11956
rect 18620 11902 18734 11954
rect 18786 11902 18788 11954
rect 18620 11900 18788 11902
rect 18396 11508 18452 11518
rect 18284 10836 18340 10846
rect 18284 10742 18340 10780
rect 18396 9826 18452 11452
rect 18508 11396 18564 11406
rect 18508 11302 18564 11340
rect 18396 9774 18398 9826
rect 18450 9774 18452 9826
rect 18396 9762 18452 9774
rect 18508 11060 18564 11070
rect 17948 5170 18004 5180
rect 18060 9212 18228 9268
rect 17500 4162 17556 4172
rect 18060 2772 18116 9212
rect 18508 9156 18564 11004
rect 18620 10724 18676 11900
rect 18732 11890 18788 11900
rect 18844 11956 18900 11966
rect 18844 11862 18900 11900
rect 19180 11732 19236 12012
rect 19404 11954 19460 12012
rect 19404 11902 19406 11954
rect 19458 11902 19460 11954
rect 19404 11890 19460 11902
rect 19516 11956 19572 11966
rect 18732 11676 19236 11732
rect 19292 11844 19348 11854
rect 18732 11618 18788 11676
rect 18732 11566 18734 11618
rect 18786 11566 18788 11618
rect 18732 11554 18788 11566
rect 19180 11508 19236 11518
rect 19180 11414 19236 11452
rect 18620 10658 18676 10668
rect 18956 10052 19012 10062
rect 18956 9958 19012 9996
rect 19292 9940 19348 11788
rect 19404 11172 19460 11182
rect 19404 10498 19460 11116
rect 19404 10446 19406 10498
rect 19458 10446 19460 10498
rect 19404 10434 19460 10446
rect 19292 9874 19348 9884
rect 19404 10164 19460 10174
rect 19404 9938 19460 10108
rect 19404 9886 19406 9938
rect 19458 9886 19460 9938
rect 19404 9874 19460 9886
rect 18844 9826 18900 9838
rect 18844 9774 18846 9826
rect 18898 9774 18900 9826
rect 18620 9156 18676 9166
rect 18508 9154 18676 9156
rect 18508 9102 18622 9154
rect 18674 9102 18676 9154
rect 18508 9100 18676 9102
rect 18620 9090 18676 9100
rect 18172 9044 18228 9054
rect 18172 8930 18228 8988
rect 18172 8878 18174 8930
rect 18226 8878 18228 8930
rect 18172 8866 18228 8878
rect 18844 8372 18900 9774
rect 18844 8306 18900 8316
rect 19516 8484 19572 11900
rect 19740 11956 19796 13244
rect 19852 13188 19908 16044
rect 20076 15428 20132 17614
rect 20076 15362 20132 15372
rect 20300 18116 20356 18126
rect 20076 15204 20132 15242
rect 20076 15138 20132 15148
rect 19964 15090 20020 15102
rect 19964 15038 19966 15090
rect 20018 15038 20020 15090
rect 19964 13972 20020 15038
rect 19964 13906 20020 13916
rect 20076 14308 20132 14318
rect 19964 13636 20020 13646
rect 19964 13542 20020 13580
rect 19852 13132 20020 13188
rect 19740 11890 19796 11900
rect 19852 12964 19908 12974
rect 19852 11394 19908 12908
rect 19964 12962 20020 13132
rect 19964 12910 19966 12962
rect 20018 12910 20020 12962
rect 19964 12404 20020 12910
rect 20076 12852 20132 14252
rect 20076 12786 20132 12796
rect 20188 13074 20244 13086
rect 20188 13022 20190 13074
rect 20242 13022 20244 13074
rect 19964 12348 20132 12404
rect 19964 12180 20020 12190
rect 19964 12086 20020 12124
rect 19852 11342 19854 11394
rect 19906 11342 19908 11394
rect 19852 11330 19908 11342
rect 20076 11396 20132 12348
rect 20188 11844 20244 13022
rect 20188 11778 20244 11788
rect 20076 11330 20132 11340
rect 19964 10836 20020 10846
rect 19852 10612 19908 10622
rect 19852 10518 19908 10556
rect 19516 8370 19572 8428
rect 19516 8318 19518 8370
rect 19570 8318 19572 8370
rect 19516 8306 19572 8318
rect 19964 8258 20020 10780
rect 19964 8206 19966 8258
rect 20018 8206 20020 8258
rect 19964 8194 20020 8206
rect 20076 9826 20132 9838
rect 20076 9774 20078 9826
rect 20130 9774 20132 9826
rect 20076 8260 20132 9774
rect 19068 8036 19124 8046
rect 18060 2706 18116 2716
rect 18508 6580 18564 6590
rect 18508 2100 18564 6524
rect 19068 5460 19124 7980
rect 20076 7252 20132 8204
rect 20300 8372 20356 18060
rect 20412 16212 20468 16222
rect 20412 13076 20468 16156
rect 20524 16098 20580 18172
rect 20636 17668 20692 18286
rect 20636 17602 20692 17612
rect 20860 17668 20916 18620
rect 20972 18450 21028 18462
rect 20972 18398 20974 18450
rect 21026 18398 21028 18450
rect 20972 18228 21028 18398
rect 20972 18162 21028 18172
rect 20860 17666 21140 17668
rect 20860 17614 20862 17666
rect 20914 17614 21140 17666
rect 20860 17612 21140 17614
rect 20860 17602 20916 17612
rect 20972 17332 21028 17342
rect 20972 16884 21028 17276
rect 20972 16790 21028 16828
rect 20748 16658 20804 16670
rect 20748 16606 20750 16658
rect 20802 16606 20804 16658
rect 20524 16046 20526 16098
rect 20578 16046 20580 16098
rect 20524 16034 20580 16046
rect 20636 16548 20692 16558
rect 20636 15652 20692 16492
rect 20748 15652 20804 16606
rect 20860 16660 20916 16670
rect 20860 16566 20916 16604
rect 20748 15596 21028 15652
rect 20636 15428 20692 15596
rect 20636 15334 20692 15372
rect 20524 15316 20580 15326
rect 20524 15148 20580 15260
rect 20972 15314 21028 15596
rect 20972 15262 20974 15314
rect 21026 15262 21028 15314
rect 20524 15092 20916 15148
rect 20524 14980 20580 14990
rect 20524 13412 20580 14924
rect 20748 14532 20804 14542
rect 20748 14438 20804 14476
rect 20860 13748 20916 15092
rect 20972 14308 21028 15262
rect 21084 15092 21140 17612
rect 21196 16100 21252 20412
rect 21308 20356 21364 22318
rect 21308 20290 21364 20300
rect 21420 22260 21476 22270
rect 21308 20020 21364 20030
rect 21308 19122 21364 19964
rect 21308 19070 21310 19122
rect 21362 19070 21364 19122
rect 21308 16548 21364 19070
rect 21420 18450 21476 22204
rect 21644 20580 21700 24108
rect 21756 20804 21812 25228
rect 21868 22484 21924 26012
rect 22092 24164 22148 24174
rect 22092 24070 22148 24108
rect 21868 22418 21924 22428
rect 22204 22148 22260 28364
rect 22316 26964 22372 26974
rect 22316 25618 22372 26908
rect 22316 25566 22318 25618
rect 22370 25566 22372 25618
rect 22316 25554 22372 25566
rect 22428 26066 22484 26078
rect 22428 26014 22430 26066
rect 22482 26014 22484 26066
rect 22316 24724 22372 24734
rect 22428 24724 22484 26014
rect 22652 24948 22708 30940
rect 23100 30212 23156 30222
rect 23100 30118 23156 30156
rect 22988 28980 23044 28990
rect 22652 24892 22820 24948
rect 22316 24722 22484 24724
rect 22316 24670 22318 24722
rect 22370 24670 22484 24722
rect 22316 24668 22484 24670
rect 22652 24722 22708 24734
rect 22652 24670 22654 24722
rect 22706 24670 22708 24722
rect 22316 24658 22372 24668
rect 22540 24052 22596 24062
rect 22540 23958 22596 23996
rect 22428 22372 22484 22382
rect 22428 22370 22596 22372
rect 22428 22318 22430 22370
rect 22482 22318 22596 22370
rect 22428 22316 22596 22318
rect 22428 22306 22484 22316
rect 22204 22092 22484 22148
rect 21980 21812 22036 21822
rect 21980 21586 22036 21756
rect 21980 21534 21982 21586
rect 22034 21534 22036 21586
rect 21980 21522 22036 21534
rect 22204 21586 22260 21598
rect 22204 21534 22206 21586
rect 22258 21534 22260 21586
rect 21756 20710 21812 20748
rect 21868 21474 21924 21486
rect 21868 21422 21870 21474
rect 21922 21422 21924 21474
rect 21644 20524 21812 20580
rect 21420 18398 21422 18450
rect 21474 18398 21476 18450
rect 21420 18116 21476 18398
rect 21644 20356 21700 20366
rect 21644 18452 21700 20300
rect 21644 18386 21700 18396
rect 21420 18050 21476 18060
rect 21532 18228 21588 18238
rect 21532 17890 21588 18172
rect 21644 18226 21700 18238
rect 21644 18174 21646 18226
rect 21698 18174 21700 18226
rect 21644 18004 21700 18174
rect 21644 17938 21700 17948
rect 21532 17838 21534 17890
rect 21586 17838 21588 17890
rect 21532 17826 21588 17838
rect 21308 16482 21364 16492
rect 21532 17668 21588 17678
rect 21196 16098 21364 16100
rect 21196 16046 21198 16098
rect 21250 16046 21364 16098
rect 21196 16044 21364 16046
rect 21196 16034 21252 16044
rect 21084 14532 21140 15036
rect 21196 15316 21252 15326
rect 21196 14980 21252 15260
rect 21196 14914 21252 14924
rect 21084 14466 21140 14476
rect 20972 14242 21028 14252
rect 21308 13748 21364 16044
rect 21420 15988 21476 15998
rect 21420 15764 21476 15932
rect 21420 15314 21476 15708
rect 21420 15262 21422 15314
rect 21474 15262 21476 15314
rect 21420 15250 21476 15262
rect 21420 14308 21476 14318
rect 21420 14214 21476 14252
rect 20524 13346 20580 13356
rect 20636 13634 20692 13646
rect 20636 13582 20638 13634
rect 20690 13582 20692 13634
rect 20412 13020 20580 13076
rect 20300 8258 20356 8316
rect 20300 8206 20302 8258
rect 20354 8206 20356 8258
rect 20300 7700 20356 8206
rect 20412 12852 20468 12862
rect 20412 8148 20468 12796
rect 20524 12516 20580 13020
rect 20524 12450 20580 12460
rect 20636 12180 20692 13582
rect 20860 13634 20916 13692
rect 21084 13692 21364 13748
rect 21420 13748 21476 13758
rect 20860 13582 20862 13634
rect 20914 13582 20916 13634
rect 20860 13570 20916 13582
rect 20972 13636 21028 13646
rect 20748 13524 20804 13534
rect 20748 13430 20804 13468
rect 20860 13412 20916 13422
rect 20860 12962 20916 13356
rect 20860 12910 20862 12962
rect 20914 12910 20916 12962
rect 20860 12898 20916 12910
rect 20972 12740 21028 13580
rect 21084 13300 21140 13692
rect 21420 13654 21476 13692
rect 21532 13524 21588 17612
rect 21644 15204 21700 15214
rect 21644 15090 21700 15148
rect 21644 15038 21646 15090
rect 21698 15038 21700 15090
rect 21644 15026 21700 15038
rect 21084 13234 21140 13244
rect 21308 13468 21588 13524
rect 21644 13748 21700 13758
rect 20748 12684 21028 12740
rect 20748 12290 20804 12684
rect 20748 12238 20750 12290
rect 20802 12238 20804 12290
rect 20748 12226 20804 12238
rect 20860 12516 20916 12526
rect 20524 12124 20692 12180
rect 20860 12178 20916 12460
rect 20860 12126 20862 12178
rect 20914 12126 20916 12178
rect 20524 8370 20580 12124
rect 20860 12114 20916 12126
rect 20636 11954 20692 11966
rect 20636 11902 20638 11954
rect 20690 11902 20692 11954
rect 20636 11844 20692 11902
rect 21084 11956 21140 11966
rect 21084 11862 21140 11900
rect 20636 11778 20692 11788
rect 20860 11508 20916 11518
rect 20860 11394 20916 11452
rect 20860 11342 20862 11394
rect 20914 11342 20916 11394
rect 20860 10276 20916 11342
rect 20860 9044 20916 10220
rect 21084 9828 21140 9838
rect 21084 9734 21140 9772
rect 20860 8978 20916 8988
rect 20524 8318 20526 8370
rect 20578 8318 20580 8370
rect 20524 8306 20580 8318
rect 20972 8260 21028 8270
rect 20636 8258 21028 8260
rect 20636 8206 20974 8258
rect 21026 8206 21028 8258
rect 20636 8204 21028 8206
rect 20636 8148 20692 8204
rect 20972 8194 21028 8204
rect 21308 8260 21364 13468
rect 21420 13300 21476 13310
rect 21420 12964 21476 13244
rect 21420 12870 21476 12908
rect 21532 12516 21588 12526
rect 21532 12402 21588 12460
rect 21532 12350 21534 12402
rect 21586 12350 21588 12402
rect 21532 12338 21588 12350
rect 21644 12178 21700 13692
rect 21644 12126 21646 12178
rect 21698 12126 21700 12178
rect 21644 12114 21700 12126
rect 21308 8194 21364 8204
rect 21420 11956 21476 11966
rect 20412 8092 20692 8148
rect 20300 7634 20356 7644
rect 20076 7186 20132 7196
rect 19068 5394 19124 5404
rect 18508 2034 18564 2044
rect 16828 1652 16884 1662
rect 16828 112 16884 1596
rect 20860 1652 20916 1662
rect 18172 1316 18228 1326
rect 18172 112 18228 1260
rect 19516 196 19572 206
rect 19516 112 19572 140
rect 20860 112 20916 1596
rect 21420 980 21476 11900
rect 21644 8260 21700 8270
rect 21644 6804 21700 8204
rect 21644 6738 21700 6748
rect 21756 3388 21812 20524
rect 21868 14532 21924 21422
rect 21980 21252 22036 21262
rect 21980 18340 22036 21196
rect 22092 20804 22148 20814
rect 22092 18564 22148 20748
rect 22204 20132 22260 21534
rect 22204 20066 22260 20076
rect 22092 18508 22260 18564
rect 21980 17556 22036 18284
rect 21980 17490 22036 17500
rect 22092 18338 22148 18350
rect 22092 18286 22094 18338
rect 22146 18286 22148 18338
rect 22092 17444 22148 18286
rect 22092 17378 22148 17388
rect 22204 16996 22260 18508
rect 22092 16940 22260 16996
rect 22092 16100 22148 16940
rect 21980 16098 22148 16100
rect 21980 16046 22094 16098
rect 22146 16046 22148 16098
rect 21980 16044 22148 16046
rect 21980 15148 22036 16044
rect 22092 16034 22148 16044
rect 22204 16658 22260 16670
rect 22204 16606 22206 16658
rect 22258 16606 22260 16658
rect 22092 15316 22148 15326
rect 22092 15222 22148 15260
rect 21980 15092 22148 15148
rect 21868 14476 22036 14532
rect 21868 14308 21924 14318
rect 21868 11732 21924 14252
rect 21868 11666 21924 11676
rect 21868 10052 21924 10062
rect 21868 8148 21924 9996
rect 21868 8082 21924 8092
rect 21980 3556 22036 14476
rect 22092 12964 22148 15092
rect 22204 14196 22260 16606
rect 22204 14130 22260 14140
rect 22204 12964 22260 12974
rect 22092 12962 22260 12964
rect 22092 12910 22206 12962
rect 22258 12910 22260 12962
rect 22092 12908 22260 12910
rect 22204 11508 22260 12908
rect 22204 11442 22260 11452
rect 21980 3490 22036 3500
rect 21644 3332 21812 3388
rect 21644 1876 21700 3332
rect 21644 1810 21700 1820
rect 22204 1988 22260 1998
rect 21420 914 21476 924
rect 22204 112 22260 1932
rect 22428 1428 22484 22092
rect 22540 18452 22596 22316
rect 22652 21252 22708 24670
rect 22652 21186 22708 21196
rect 22764 20020 22820 24892
rect 22764 19954 22820 19964
rect 22876 22484 22932 22494
rect 22876 22370 22932 22428
rect 22876 22318 22878 22370
rect 22930 22318 22932 22370
rect 22876 19796 22932 22318
rect 22764 19740 22932 19796
rect 22540 18386 22596 18396
rect 22652 18450 22708 18462
rect 22652 18398 22654 18450
rect 22706 18398 22708 18450
rect 22652 18340 22708 18398
rect 22652 17668 22708 18284
rect 22764 17778 22820 19740
rect 22764 17726 22766 17778
rect 22818 17726 22820 17778
rect 22764 17714 22820 17726
rect 22876 18452 22932 18462
rect 22652 17602 22708 17612
rect 22540 16324 22596 16334
rect 22540 14754 22596 16268
rect 22540 14702 22542 14754
rect 22594 14702 22596 14754
rect 22540 14690 22596 14702
rect 22764 15314 22820 15326
rect 22764 15262 22766 15314
rect 22818 15262 22820 15314
rect 22652 14642 22708 14654
rect 22652 14590 22654 14642
rect 22706 14590 22708 14642
rect 22540 13522 22596 13534
rect 22540 13470 22542 13522
rect 22594 13470 22596 13522
rect 22540 13188 22596 13470
rect 22540 13122 22596 13132
rect 22540 11954 22596 11966
rect 22540 11902 22542 11954
rect 22594 11902 22596 11954
rect 22540 8428 22596 11902
rect 22652 11844 22708 14590
rect 22764 14644 22820 15262
rect 22764 13860 22820 14588
rect 22764 13794 22820 13804
rect 22652 11778 22708 11788
rect 22876 9828 22932 18396
rect 22988 15316 23044 28924
rect 23100 24612 23156 24622
rect 23100 24050 23156 24556
rect 23100 23998 23102 24050
rect 23154 23998 23156 24050
rect 23100 23986 23156 23998
rect 23324 17780 23380 42812
rect 23436 22932 23492 43652
rect 24892 43538 24948 43550
rect 24892 43486 24894 43538
rect 24946 43486 24948 43538
rect 24464 43148 24728 43158
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24464 43082 24728 43092
rect 24668 42754 24724 42766
rect 24668 42702 24670 42754
rect 24722 42702 24724 42754
rect 24668 42644 24724 42702
rect 24668 42578 24724 42588
rect 23804 42364 24068 42374
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 23804 42298 24068 42308
rect 24464 41580 24728 41590
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24464 41514 24728 41524
rect 24780 41186 24836 41198
rect 24780 41134 24782 41186
rect 24834 41134 24836 41186
rect 23804 40796 24068 40806
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 23804 40730 24068 40740
rect 24668 40292 24724 40302
rect 24220 40290 24724 40292
rect 24220 40238 24670 40290
rect 24722 40238 24724 40290
rect 24220 40236 24724 40238
rect 23804 39228 24068 39238
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 23804 39162 24068 39172
rect 23660 37940 23716 37950
rect 23660 31780 23716 37884
rect 23804 37660 24068 37670
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 23804 37594 24068 37604
rect 23804 36092 24068 36102
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 23804 36026 24068 36036
rect 23804 34524 24068 34534
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 23804 34458 24068 34468
rect 23804 32956 24068 32966
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 23804 32890 24068 32900
rect 24220 32004 24276 40236
rect 24668 40226 24724 40236
rect 24780 40180 24836 41134
rect 24780 40114 24836 40124
rect 24464 40012 24728 40022
rect 24332 39956 24388 39966
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24464 39946 24728 39956
rect 24332 36596 24388 39900
rect 24668 39620 24724 39630
rect 24668 39526 24724 39564
rect 24464 38444 24728 38454
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24464 38378 24728 38388
rect 24892 38276 24948 43486
rect 24892 38210 24948 38220
rect 24892 38050 24948 38062
rect 24892 37998 24894 38050
rect 24946 37998 24948 38050
rect 24668 37156 24724 37166
rect 24668 37062 24724 37100
rect 24464 36876 24728 36886
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24464 36810 24728 36820
rect 24668 36596 24724 36606
rect 24332 36594 24724 36596
rect 24332 36542 24670 36594
rect 24722 36542 24724 36594
rect 24332 36540 24724 36542
rect 24668 36530 24724 36540
rect 24892 36260 24948 37998
rect 24892 36194 24948 36204
rect 24464 35308 24728 35318
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24464 35242 24728 35252
rect 24668 34914 24724 34926
rect 24668 34862 24670 34914
rect 24722 34862 24724 34914
rect 24668 33908 24724 34862
rect 24892 34132 24948 34142
rect 24892 34130 25172 34132
rect 24892 34078 24894 34130
rect 24946 34078 25172 34130
rect 24892 34076 25172 34078
rect 24892 34066 24948 34076
rect 24668 33842 24724 33852
rect 24464 33740 24728 33750
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24464 33674 24728 33684
rect 24892 33346 24948 33358
rect 24892 33294 24894 33346
rect 24946 33294 24948 33346
rect 24464 32172 24728 32182
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24464 32106 24728 32116
rect 24220 31938 24276 31948
rect 24780 31892 24836 31902
rect 24668 31780 24724 31790
rect 23660 31778 24724 31780
rect 23660 31726 24670 31778
rect 24722 31726 24724 31778
rect 23660 31724 24724 31726
rect 24668 31714 24724 31724
rect 23660 31444 23716 31454
rect 23660 30996 23716 31388
rect 23804 31388 24068 31398
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 23804 31322 24068 31332
rect 23660 30902 23716 30940
rect 24780 30994 24836 31836
rect 24892 31220 24948 33294
rect 24892 31154 24948 31164
rect 24780 30942 24782 30994
rect 24834 30942 24836 30994
rect 24780 30930 24836 30942
rect 24464 30604 24728 30614
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24464 30538 24728 30548
rect 23804 29820 24068 29830
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 23804 29754 24068 29764
rect 24464 29036 24728 29046
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24464 28970 24728 28980
rect 23804 28252 24068 28262
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 23804 28186 24068 28196
rect 25004 28084 25060 28094
rect 24892 27858 24948 27870
rect 24892 27806 24894 27858
rect 24946 27806 24948 27858
rect 24464 27468 24728 27478
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24464 27402 24728 27412
rect 24892 27300 24948 27806
rect 24892 27234 24948 27244
rect 24668 27074 24724 27086
rect 24668 27022 24670 27074
rect 24722 27022 24724 27074
rect 24668 26908 24724 27022
rect 24220 26852 24724 26908
rect 23804 26684 24068 26694
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 23804 26618 24068 26628
rect 23804 25116 24068 25126
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 23804 25050 24068 25060
rect 23660 24722 23716 24734
rect 23660 24670 23662 24722
rect 23714 24670 23716 24722
rect 23436 22866 23492 22876
rect 23548 23492 23604 23502
rect 23436 22484 23492 22494
rect 23436 22390 23492 22428
rect 23548 22148 23604 23436
rect 23548 21586 23604 22092
rect 23548 21534 23550 21586
rect 23602 21534 23604 21586
rect 23548 21522 23604 21534
rect 23660 18676 23716 24670
rect 23804 23548 24068 23558
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 23804 23482 24068 23492
rect 23804 21980 24068 21990
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 23804 21914 24068 21924
rect 23996 21700 24052 21710
rect 23996 21606 24052 21644
rect 23804 20412 24068 20422
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 23804 20346 24068 20356
rect 24220 19460 24276 26852
rect 24332 26180 24388 26190
rect 24332 24164 24388 26124
rect 24464 25900 24728 25910
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24464 25834 24728 25844
rect 24668 25506 24724 25518
rect 24668 25454 24670 25506
rect 24722 25454 24724 25506
rect 24668 24500 24724 25454
rect 24668 24434 24724 24444
rect 24892 24722 24948 24734
rect 24892 24670 24894 24722
rect 24946 24670 24948 24722
rect 24464 24332 24728 24342
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24464 24266 24728 24276
rect 24332 24108 24724 24164
rect 24668 24050 24724 24108
rect 24668 23998 24670 24050
rect 24722 23998 24724 24050
rect 24668 23986 24724 23998
rect 24892 23268 24948 24670
rect 24892 23202 24948 23212
rect 24464 22764 24728 22774
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24464 22698 24728 22708
rect 24892 22372 24948 22382
rect 25004 22372 25060 28028
rect 25116 26516 25172 34076
rect 25340 26908 25396 55244
rect 25564 54626 25620 57372
rect 25900 57316 25956 57372
rect 26208 57344 26320 57456
rect 27552 57344 27664 57456
rect 25900 57250 25956 57260
rect 26236 57316 26292 57344
rect 26236 57250 26292 57260
rect 25788 56756 25844 56766
rect 25564 54574 25566 54626
rect 25618 54574 25620 54626
rect 25564 54562 25620 54574
rect 25676 55074 25732 55086
rect 25676 55022 25678 55074
rect 25730 55022 25732 55074
rect 25676 54516 25732 55022
rect 25676 54450 25732 54460
rect 25676 53620 25732 53630
rect 25676 53526 25732 53564
rect 25452 52834 25508 52846
rect 25452 52782 25454 52834
rect 25506 52782 25508 52834
rect 25452 52724 25508 52782
rect 25452 52658 25508 52668
rect 25676 51938 25732 51950
rect 25676 51886 25678 51938
rect 25730 51886 25732 51938
rect 25676 51828 25732 51886
rect 25676 51762 25732 51772
rect 25676 51604 25732 51614
rect 25788 51604 25844 56700
rect 27580 56644 27636 57344
rect 27580 56578 27636 56588
rect 26012 56308 26068 56318
rect 26012 56214 26068 56252
rect 26236 55300 26292 55310
rect 26236 55206 26292 55244
rect 27244 55074 27300 55086
rect 27244 55022 27246 55074
rect 27298 55022 27300 55074
rect 26348 54514 26404 54526
rect 26348 54462 26350 54514
rect 26402 54462 26404 54514
rect 26236 53730 26292 53742
rect 26236 53678 26238 53730
rect 26290 53678 26292 53730
rect 26236 53172 26292 53678
rect 26236 53106 26292 53116
rect 26236 52388 26292 52398
rect 26236 52274 26292 52332
rect 26236 52222 26238 52274
rect 26290 52222 26292 52274
rect 26236 52210 26292 52222
rect 25676 51602 25844 51604
rect 25676 51550 25678 51602
rect 25730 51550 25844 51602
rect 25676 51548 25844 51550
rect 25676 51538 25732 51548
rect 26236 51266 26292 51278
rect 26236 51214 26238 51266
rect 26290 51214 26292 51266
rect 26236 51156 26292 51214
rect 26236 51090 26292 51100
rect 26236 50708 26292 50718
rect 26236 50614 26292 50652
rect 25676 50484 25732 50494
rect 25676 50390 25732 50428
rect 25676 49922 25732 49934
rect 25676 49870 25678 49922
rect 25730 49870 25732 49922
rect 25676 49588 25732 49870
rect 25676 49522 25732 49532
rect 26236 49698 26292 49710
rect 26236 49646 26238 49698
rect 26290 49646 26292 49698
rect 26236 49252 26292 49646
rect 26236 49186 26292 49196
rect 26236 49026 26292 49038
rect 26236 48974 26238 49026
rect 26290 48974 26292 49026
rect 26236 48916 26292 48974
rect 26236 48850 26292 48860
rect 25676 48802 25732 48814
rect 25676 48750 25678 48802
rect 25730 48750 25732 48802
rect 25676 48692 25732 48750
rect 25676 48626 25732 48636
rect 26236 47460 26292 47470
rect 26236 47366 26292 47404
rect 25676 47348 25732 47358
rect 25676 47254 25732 47292
rect 25676 46786 25732 46798
rect 25676 46734 25678 46786
rect 25730 46734 25732 46786
rect 25676 46452 25732 46734
rect 25676 46386 25732 46396
rect 26236 46562 26292 46574
rect 26236 46510 26238 46562
rect 26290 46510 26292 46562
rect 26236 46116 26292 46510
rect 26236 46050 26292 46060
rect 26236 45892 26292 45902
rect 25788 45890 26292 45892
rect 25788 45838 26238 45890
rect 26290 45838 26292 45890
rect 25788 45836 26292 45838
rect 25676 45666 25732 45678
rect 25676 45614 25678 45666
rect 25730 45614 25732 45666
rect 25676 45556 25732 45614
rect 25676 45490 25732 45500
rect 25564 44324 25620 44334
rect 25452 37154 25508 37166
rect 25452 37102 25454 37154
rect 25506 37102 25508 37154
rect 25452 37044 25508 37102
rect 25452 36978 25508 36988
rect 25564 35812 25620 44268
rect 25676 44212 25732 44222
rect 25676 44118 25732 44156
rect 25676 43650 25732 43662
rect 25676 43598 25678 43650
rect 25730 43598 25732 43650
rect 25676 43316 25732 43598
rect 25676 43250 25732 43260
rect 25676 42530 25732 42542
rect 25676 42478 25678 42530
rect 25730 42478 25732 42530
rect 25676 42420 25732 42478
rect 25676 42354 25732 42364
rect 25676 41076 25732 41086
rect 25676 40982 25732 41020
rect 25676 40514 25732 40526
rect 25676 40462 25678 40514
rect 25730 40462 25732 40514
rect 25676 40180 25732 40462
rect 25788 40292 25844 45836
rect 26236 45826 26292 45836
rect 26236 44996 26292 45006
rect 26236 44902 26292 44940
rect 26236 44324 26292 44334
rect 26236 44230 26292 44268
rect 26348 43876 26404 54462
rect 27020 54402 27076 54414
rect 27020 54350 27022 54402
rect 27074 54350 27076 54402
rect 27020 53172 27076 54350
rect 27244 54068 27300 55022
rect 27244 54002 27300 54012
rect 27020 53106 27076 53116
rect 27244 53506 27300 53518
rect 27244 53454 27246 53506
rect 27298 53454 27300 53506
rect 27132 53058 27188 53070
rect 27132 53006 27134 53058
rect 27186 53006 27188 53058
rect 26460 52946 26516 52958
rect 26460 52894 26462 52946
rect 26514 52894 26516 52946
rect 26460 48468 26516 52894
rect 26460 48402 26516 48412
rect 26572 52164 26628 52174
rect 26236 43820 26404 43876
rect 26460 48242 26516 48254
rect 26460 48190 26462 48242
rect 26514 48190 26516 48242
rect 26236 43708 26292 43820
rect 26460 43708 26516 48190
rect 25788 40226 25844 40236
rect 25900 43652 26292 43708
rect 26348 43652 26516 43708
rect 25676 40114 25732 40124
rect 25676 39394 25732 39406
rect 25676 39342 25678 39394
rect 25730 39342 25732 39394
rect 25676 39284 25732 39342
rect 25676 39218 25732 39228
rect 25676 37940 25732 37950
rect 25676 37846 25732 37884
rect 25676 36258 25732 36270
rect 25676 36206 25678 36258
rect 25730 36206 25732 36258
rect 25676 36148 25732 36206
rect 25676 36082 25732 36092
rect 25564 35746 25620 35756
rect 25788 35140 25844 35150
rect 25676 34804 25732 34814
rect 25676 34710 25732 34748
rect 25676 34242 25732 34254
rect 25676 34190 25678 34242
rect 25730 34190 25732 34242
rect 25676 33908 25732 34190
rect 25676 33842 25732 33852
rect 25676 33122 25732 33134
rect 25676 33070 25678 33122
rect 25730 33070 25732 33122
rect 25676 33012 25732 33070
rect 25676 32946 25732 32956
rect 25676 31668 25732 31678
rect 25676 31574 25732 31612
rect 25452 30882 25508 30894
rect 25452 30830 25454 30882
rect 25506 30830 25508 30882
rect 25452 30772 25508 30830
rect 25452 30706 25508 30716
rect 25788 29428 25844 35084
rect 25788 29362 25844 29372
rect 25788 29204 25844 29214
rect 25676 27970 25732 27982
rect 25676 27918 25678 27970
rect 25730 27918 25732 27970
rect 25676 27188 25732 27918
rect 25676 27122 25732 27132
rect 25340 26852 25508 26908
rect 25116 26450 25172 26460
rect 24892 22370 25060 22372
rect 24892 22318 24894 22370
rect 24946 22318 25060 22370
rect 24892 22316 25060 22318
rect 25228 26292 25284 26302
rect 24892 22306 24948 22316
rect 24220 19394 24276 19404
rect 24332 22148 24388 22158
rect 23804 18844 24068 18854
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 23804 18778 24068 18788
rect 23324 17714 23380 17724
rect 23548 18620 23716 18676
rect 22988 15250 23044 15260
rect 23100 17554 23156 17566
rect 23100 17502 23102 17554
rect 23154 17502 23156 17554
rect 23100 15148 23156 17502
rect 23548 17108 23604 18620
rect 23660 18452 23716 18462
rect 23660 18358 23716 18396
rect 23804 17276 24068 17286
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 23804 17210 24068 17220
rect 23548 17042 23604 17052
rect 23884 16884 23940 16894
rect 23884 16882 24276 16884
rect 23884 16830 23886 16882
rect 23938 16830 24276 16882
rect 23884 16828 24276 16830
rect 23884 16818 23940 16828
rect 22988 15092 23156 15148
rect 23324 16658 23380 16670
rect 23324 16606 23326 16658
rect 23378 16606 23380 16658
rect 22988 14418 23044 15092
rect 22988 14366 22990 14418
rect 23042 14366 23044 14418
rect 22988 13746 23044 14366
rect 22988 13694 22990 13746
rect 23042 13694 23044 13746
rect 22988 10612 23044 13694
rect 23324 13188 23380 16606
rect 23804 15708 24068 15718
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 23804 15642 24068 15652
rect 23772 15314 23828 15326
rect 23772 15262 23774 15314
rect 23826 15262 23828 15314
rect 23772 15148 23828 15262
rect 23660 15092 23828 15148
rect 23660 13972 23716 15036
rect 23804 14140 24068 14150
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 23804 14074 24068 14084
rect 23660 13916 23828 13972
rect 23324 13122 23380 13132
rect 23660 13522 23716 13534
rect 23660 13470 23662 13522
rect 23714 13470 23716 13522
rect 23660 12628 23716 13470
rect 23772 13524 23828 13916
rect 23772 13458 23828 13468
rect 24220 13748 24276 16828
rect 24332 13860 24388 22092
rect 25004 21812 25060 21822
rect 24464 21196 24728 21206
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24464 21130 24728 21140
rect 25004 20914 25060 21756
rect 25004 20862 25006 20914
rect 25058 20862 25060 20914
rect 25004 20850 25060 20862
rect 24464 19628 24728 19638
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24464 19562 24728 19572
rect 24464 18060 24728 18070
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24464 17994 24728 18004
rect 24556 17780 24612 17790
rect 24556 17686 24612 17724
rect 25228 17780 25284 26236
rect 25340 21362 25396 21374
rect 25340 21310 25342 21362
rect 25394 21310 25396 21362
rect 25340 20580 25396 21310
rect 25340 20514 25396 20524
rect 25228 17714 25284 17724
rect 25340 19124 25396 19134
rect 25116 17666 25172 17678
rect 25116 17614 25118 17666
rect 25170 17614 25172 17666
rect 24464 16492 24728 16502
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24464 16426 24728 16436
rect 25116 15148 25172 17614
rect 24892 15092 25172 15148
rect 24464 14924 24728 14934
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24464 14858 24728 14868
rect 24780 14420 24836 14430
rect 24892 14420 24948 15092
rect 24780 14418 24948 14420
rect 24780 14366 24782 14418
rect 24834 14366 24948 14418
rect 24780 14364 24948 14366
rect 24780 14354 24836 14364
rect 24332 13804 24836 13860
rect 24220 12740 24276 13692
rect 24332 13636 24388 13646
rect 24332 13076 24388 13580
rect 24780 13634 24836 13804
rect 24892 13748 24948 14364
rect 24892 13682 24948 13692
rect 25116 14642 25172 14654
rect 25116 14590 25118 14642
rect 25170 14590 25172 14642
rect 24780 13582 24782 13634
rect 24834 13582 24836 13634
rect 24780 13570 24836 13582
rect 24464 13356 24728 13366
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24464 13290 24728 13300
rect 25116 13186 25172 14590
rect 25228 13748 25284 13786
rect 25228 13682 25284 13692
rect 25116 13134 25118 13186
rect 25170 13134 25172 13186
rect 25116 13122 25172 13134
rect 25228 13524 25284 13534
rect 24556 13076 24612 13086
rect 24332 13074 24612 13076
rect 24332 13022 24558 13074
rect 24610 13022 24612 13074
rect 24332 13020 24612 13022
rect 24556 13010 24612 13020
rect 23660 12562 23716 12572
rect 23804 12572 24068 12582
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 23804 12506 24068 12516
rect 24220 12178 24276 12684
rect 24220 12126 24222 12178
rect 24274 12126 24276 12178
rect 24220 12114 24276 12126
rect 25004 12962 25060 12974
rect 25004 12910 25006 12962
rect 25058 12910 25060 12962
rect 23660 11954 23716 11966
rect 23660 11902 23662 11954
rect 23714 11902 23716 11954
rect 23212 11844 23268 11854
rect 23212 11618 23268 11788
rect 23660 11844 23716 11902
rect 23660 11778 23716 11788
rect 24464 11788 24728 11798
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24464 11722 24728 11732
rect 23212 11566 23214 11618
rect 23266 11566 23268 11618
rect 23212 11554 23268 11566
rect 23772 11508 23828 11518
rect 23772 11414 23828 11452
rect 25004 11172 25060 12910
rect 25004 11106 25060 11116
rect 23804 11004 24068 11014
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 23804 10938 24068 10948
rect 22988 10546 23044 10556
rect 24464 10220 24728 10230
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24464 10154 24728 10164
rect 22540 8372 22708 8428
rect 22540 8260 22596 8270
rect 22540 7476 22596 8204
rect 22652 7588 22708 8372
rect 22876 8260 22932 9772
rect 25116 9716 25172 9726
rect 25116 9622 25172 9660
rect 23804 9436 24068 9446
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 23804 9370 24068 9380
rect 24464 8652 24728 8662
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24464 8586 24728 8596
rect 22876 8194 22932 8204
rect 23804 7868 24068 7878
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 23804 7802 24068 7812
rect 22652 7522 22708 7532
rect 22540 7410 22596 7420
rect 24464 7084 24728 7094
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24464 7018 24728 7028
rect 23324 6692 23380 6702
rect 23324 2212 23380 6636
rect 23804 6300 24068 6310
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 23804 6234 24068 6244
rect 24892 5908 24948 5918
rect 24464 5516 24728 5526
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24464 5450 24728 5460
rect 23804 4732 24068 4742
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 23804 4666 24068 4676
rect 24464 3948 24728 3958
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24464 3882 24728 3892
rect 23804 3164 24068 3174
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 23804 3098 24068 3108
rect 24464 2380 24728 2390
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24464 2314 24728 2324
rect 23324 2146 23380 2156
rect 23804 1596 24068 1606
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 23804 1530 24068 1540
rect 22428 1362 22484 1372
rect 24892 1314 24948 5852
rect 25228 2882 25284 13468
rect 25340 11732 25396 19068
rect 25340 11666 25396 11676
rect 25452 11508 25508 26852
rect 25676 26850 25732 26862
rect 25676 26798 25678 26850
rect 25730 26798 25732 26850
rect 25676 26292 25732 26798
rect 25676 26226 25732 26236
rect 25676 25282 25732 25294
rect 25676 25230 25678 25282
rect 25730 25230 25732 25282
rect 25676 24948 25732 25230
rect 25676 24882 25732 24892
rect 25564 24834 25620 24846
rect 25564 24782 25566 24834
rect 25618 24782 25620 24834
rect 25564 24052 25620 24782
rect 25564 23986 25620 23996
rect 25676 23714 25732 23726
rect 25676 23662 25678 23714
rect 25730 23662 25732 23714
rect 25676 23156 25732 23662
rect 25676 23090 25732 23100
rect 25564 22932 25620 22942
rect 25564 21588 25620 22876
rect 25676 22146 25732 22158
rect 25676 22094 25678 22146
rect 25730 22094 25732 22146
rect 25676 21812 25732 22094
rect 25676 21746 25732 21756
rect 25564 21532 25732 21588
rect 25564 20802 25620 20814
rect 25564 20750 25566 20802
rect 25618 20750 25620 20802
rect 25564 20132 25620 20750
rect 25564 20066 25620 20076
rect 25676 19908 25732 21532
rect 25452 11442 25508 11452
rect 25564 19852 25732 19908
rect 25340 11396 25396 11406
rect 25340 9154 25396 11340
rect 25340 9102 25342 9154
rect 25394 9102 25396 9154
rect 25340 9090 25396 9102
rect 25340 7476 25396 7486
rect 25340 6018 25396 7420
rect 25340 5966 25342 6018
rect 25394 5966 25396 6018
rect 25340 5954 25396 5966
rect 25564 5796 25620 19852
rect 25676 14532 25732 14542
rect 25676 10052 25732 14476
rect 25676 9986 25732 9996
rect 25676 9826 25732 9838
rect 25676 9774 25678 9826
rect 25730 9774 25732 9826
rect 25676 9268 25732 9774
rect 25676 9202 25732 9212
rect 25564 5730 25620 5740
rect 25788 3388 25844 29148
rect 25900 21700 25956 43652
rect 26236 43428 26292 43438
rect 26124 43426 26292 43428
rect 26124 43374 26238 43426
rect 26290 43374 26292 43426
rect 26124 43372 26292 43374
rect 26012 41748 26068 41758
rect 26012 31108 26068 41692
rect 26124 41412 26180 43372
rect 26236 43362 26292 43372
rect 26236 42756 26292 42766
rect 26236 42662 26292 42700
rect 26236 41860 26292 41870
rect 26236 41766 26292 41804
rect 26124 41346 26180 41356
rect 26236 40404 26292 40414
rect 26236 40310 26292 40348
rect 26236 39618 26292 39630
rect 26236 39566 26238 39618
rect 26290 39566 26292 39618
rect 26236 39060 26292 39566
rect 26236 38994 26292 39004
rect 26236 38724 26292 38734
rect 26236 38630 26292 38668
rect 26236 38052 26292 38062
rect 26236 37958 26292 37996
rect 26236 37156 26292 37166
rect 26124 37154 26292 37156
rect 26124 37102 26238 37154
rect 26290 37102 26292 37154
rect 26124 37100 26292 37102
rect 26124 36372 26180 37100
rect 26236 37090 26292 37100
rect 26124 36306 26180 36316
rect 26236 36482 26292 36494
rect 26236 36430 26238 36482
rect 26290 36430 26292 36482
rect 26236 35924 26292 36430
rect 26236 35858 26292 35868
rect 26236 35588 26292 35598
rect 26124 35586 26292 35588
rect 26124 35534 26238 35586
rect 26290 35534 26292 35586
rect 26124 35532 26292 35534
rect 26124 34356 26180 35532
rect 26236 35522 26292 35532
rect 26236 34914 26292 34926
rect 26236 34862 26238 34914
rect 26290 34862 26292 34914
rect 26236 34692 26292 34862
rect 26236 34626 26292 34636
rect 26124 34290 26180 34300
rect 26236 34020 26292 34030
rect 26124 34018 26292 34020
rect 26124 33966 26238 34018
rect 26290 33966 26292 34018
rect 26124 33964 26292 33966
rect 26124 32788 26180 33964
rect 26236 33954 26292 33964
rect 26124 32722 26180 32732
rect 26236 33346 26292 33358
rect 26236 33294 26238 33346
rect 26290 33294 26292 33346
rect 26236 32676 26292 33294
rect 26236 32610 26292 32620
rect 26348 31444 26404 43652
rect 26460 41186 26516 41198
rect 26460 41134 26462 41186
rect 26514 41134 26516 41186
rect 26460 35028 26516 41134
rect 26460 34962 26516 34972
rect 26460 32564 26516 32574
rect 26460 32470 26516 32508
rect 26460 31780 26516 31790
rect 26460 31686 26516 31724
rect 26348 31378 26404 31388
rect 26012 31052 26516 31108
rect 26236 30882 26292 30894
rect 26236 30830 26238 30882
rect 26290 30830 26292 30882
rect 26236 30436 26292 30830
rect 26236 30370 26292 30380
rect 26236 30212 26292 30222
rect 26124 30210 26292 30212
rect 26124 30158 26238 30210
rect 26290 30158 26292 30210
rect 26124 30156 26292 30158
rect 26124 28532 26180 30156
rect 26236 30146 26292 30156
rect 26236 29428 26292 29438
rect 26236 29334 26292 29372
rect 26348 29316 26404 29326
rect 26236 28644 26292 28654
rect 26236 28550 26292 28588
rect 26124 28466 26180 28476
rect 26124 27972 26180 27982
rect 26124 24724 26180 27916
rect 26236 27748 26292 27758
rect 26236 27654 26292 27692
rect 26236 27076 26292 27086
rect 26236 26982 26292 27020
rect 26236 26180 26292 26190
rect 26236 26086 26292 26124
rect 26236 25732 26292 25742
rect 26236 25618 26292 25676
rect 26236 25566 26238 25618
rect 26290 25566 26292 25618
rect 26236 25554 26292 25566
rect 26236 24724 26292 24734
rect 26124 24722 26292 24724
rect 26124 24670 26238 24722
rect 26290 24670 26292 24722
rect 26124 24668 26292 24670
rect 26236 24658 26292 24668
rect 26236 23940 26292 23950
rect 26236 23846 26292 23884
rect 25900 21634 25956 21644
rect 26124 23828 26180 23838
rect 25900 21474 25956 21486
rect 25900 21422 25902 21474
rect 25954 21422 25956 21474
rect 25900 21364 25956 21422
rect 26124 21364 26180 23772
rect 26236 23044 26292 23054
rect 26236 22950 26292 22988
rect 26236 22596 26292 22606
rect 26236 22482 26292 22540
rect 26236 22430 26238 22482
rect 26290 22430 26292 22482
rect 26236 22418 26292 22430
rect 26236 21588 26292 21598
rect 26236 21494 26292 21532
rect 26124 21308 26292 21364
rect 25900 21298 25956 21308
rect 25900 20804 25956 20814
rect 25900 20710 25956 20748
rect 26012 20020 26068 20030
rect 26012 19926 26068 19964
rect 26012 19796 26068 19806
rect 25900 19348 25956 19358
rect 25900 19254 25956 19292
rect 25900 18676 25956 18686
rect 25900 16212 25956 18620
rect 26012 18450 26068 19740
rect 26012 18398 26014 18450
rect 26066 18398 26068 18450
rect 26012 18386 26068 18398
rect 26012 17780 26068 17790
rect 26012 17686 26068 17724
rect 26012 16996 26068 17006
rect 26012 16902 26068 16940
rect 26012 16212 26068 16222
rect 25900 16210 26068 16212
rect 25900 16158 26014 16210
rect 26066 16158 26068 16210
rect 25900 16156 26068 16158
rect 26012 16146 26068 16156
rect 26012 15876 26068 15886
rect 26012 15426 26068 15820
rect 26012 15374 26014 15426
rect 26066 15374 26068 15426
rect 26012 15362 26068 15374
rect 26012 15204 26068 15214
rect 26012 13858 26068 15148
rect 26236 15204 26292 21308
rect 26236 15138 26292 15148
rect 26348 14532 26404 29260
rect 26460 20914 26516 31052
rect 26572 22484 26628 52108
rect 27132 51380 27188 53006
rect 27244 52276 27300 53454
rect 27244 52210 27300 52220
rect 27132 51314 27188 51324
rect 27244 51938 27300 51950
rect 27244 51886 27246 51938
rect 27298 51886 27300 51938
rect 27020 51266 27076 51278
rect 27020 51214 27022 51266
rect 27074 51214 27076 51266
rect 27020 50036 27076 51214
rect 27244 50932 27300 51886
rect 27244 50866 27300 50876
rect 27020 49970 27076 49980
rect 27244 50370 27300 50382
rect 27244 50318 27246 50370
rect 27298 50318 27300 50370
rect 27132 49922 27188 49934
rect 27132 49870 27134 49922
rect 27186 49870 27188 49922
rect 27132 48244 27188 49870
rect 27244 49140 27300 50318
rect 27244 49074 27300 49084
rect 27132 48178 27188 48188
rect 27244 48802 27300 48814
rect 27244 48750 27246 48802
rect 27298 48750 27300 48802
rect 27020 48130 27076 48142
rect 27020 48078 27022 48130
rect 27074 48078 27076 48130
rect 27020 46900 27076 48078
rect 27244 47796 27300 48750
rect 27244 47730 27300 47740
rect 27356 48468 27412 48478
rect 27020 46834 27076 46844
rect 27244 47234 27300 47246
rect 27244 47182 27246 47234
rect 27298 47182 27300 47234
rect 27132 46786 27188 46798
rect 27132 46734 27134 46786
rect 27186 46734 27188 46786
rect 27132 45108 27188 46734
rect 27244 46004 27300 47182
rect 27244 45938 27300 45948
rect 27132 45042 27188 45052
rect 27244 45666 27300 45678
rect 27244 45614 27246 45666
rect 27298 45614 27300 45666
rect 27020 44994 27076 45006
rect 27020 44942 27022 44994
rect 27074 44942 27076 44994
rect 27020 43764 27076 44942
rect 27244 44660 27300 45614
rect 27244 44594 27300 44604
rect 27356 44436 27412 48412
rect 27020 43698 27076 43708
rect 27132 44380 27412 44436
rect 26908 43650 26964 43662
rect 26908 43598 26910 43650
rect 26962 43598 26964 43650
rect 26908 41972 26964 43598
rect 26908 41906 26964 41916
rect 27020 41858 27076 41870
rect 27020 41806 27022 41858
rect 27074 41806 27076 41858
rect 27020 40628 27076 41806
rect 27020 40562 27076 40572
rect 27020 40290 27076 40302
rect 27020 40238 27022 40290
rect 27074 40238 27076 40290
rect 27020 38948 27076 40238
rect 27020 38882 27076 38892
rect 27020 38722 27076 38734
rect 27020 38670 27022 38722
rect 27074 38670 27076 38722
rect 26908 37938 26964 37950
rect 26908 37886 26910 37938
rect 26962 37886 26964 37938
rect 26572 22418 26628 22428
rect 26684 37380 26740 37390
rect 26460 20862 26462 20914
rect 26514 20862 26516 20914
rect 26460 20850 26516 20862
rect 26684 20916 26740 37324
rect 26908 36596 26964 37886
rect 27020 37492 27076 38670
rect 27132 37828 27188 44380
rect 27244 44098 27300 44110
rect 27244 44046 27246 44098
rect 27298 44046 27300 44098
rect 27244 42868 27300 44046
rect 27244 42802 27300 42812
rect 27244 42530 27300 42542
rect 27244 42478 27246 42530
rect 27298 42478 27300 42530
rect 27244 41524 27300 42478
rect 27244 41458 27300 41468
rect 27468 41188 27524 41198
rect 27244 40962 27300 40974
rect 27244 40910 27246 40962
rect 27298 40910 27300 40962
rect 27244 39732 27300 40910
rect 27244 39666 27300 39676
rect 27244 39394 27300 39406
rect 27244 39342 27246 39394
rect 27298 39342 27300 39394
rect 27244 38388 27300 39342
rect 27244 38322 27300 38332
rect 27132 37772 27412 37828
rect 27020 37426 27076 37436
rect 26908 36530 26964 36540
rect 27132 37378 27188 37390
rect 27132 37326 27134 37378
rect 27186 37326 27188 37378
rect 27132 35700 27188 37326
rect 27132 35634 27188 35644
rect 27244 36258 27300 36270
rect 27244 36206 27246 36258
rect 27298 36206 27300 36258
rect 27020 35586 27076 35598
rect 27020 35534 27022 35586
rect 27074 35534 27076 35586
rect 27020 34356 27076 35534
rect 27244 35252 27300 36206
rect 27244 35186 27300 35196
rect 27020 34290 27076 34300
rect 27244 34690 27300 34702
rect 27244 34638 27246 34690
rect 27298 34638 27300 34690
rect 27132 34242 27188 34254
rect 27132 34190 27134 34242
rect 27186 34190 27188 34242
rect 27132 32564 27188 34190
rect 27244 33460 27300 34638
rect 27244 33394 27300 33404
rect 27132 32498 27188 32508
rect 27244 33122 27300 33134
rect 27244 33070 27246 33122
rect 27298 33070 27300 33122
rect 27020 32450 27076 32462
rect 27020 32398 27022 32450
rect 27074 32398 27076 32450
rect 27020 31220 27076 32398
rect 27132 32340 27188 32350
rect 27132 31948 27188 32284
rect 27244 32116 27300 33070
rect 27244 32050 27300 32060
rect 27132 31892 27300 31948
rect 27020 31154 27076 31164
rect 27132 31666 27188 31678
rect 27132 31614 27134 31666
rect 27186 31614 27188 31666
rect 27020 30882 27076 30894
rect 27020 30830 27022 30882
rect 27074 30830 27076 30882
rect 27020 29876 27076 30830
rect 27132 30324 27188 31614
rect 27132 30258 27188 30268
rect 27020 29810 27076 29820
rect 27132 30098 27188 30110
rect 27132 30046 27134 30098
rect 27186 30046 27188 30098
rect 26908 29540 26964 29550
rect 26908 21028 26964 29484
rect 27132 29428 27188 30046
rect 27132 29362 27188 29372
rect 27020 29314 27076 29326
rect 27020 29262 27022 29314
rect 27074 29262 27076 29314
rect 27020 28980 27076 29262
rect 27020 28914 27076 28924
rect 27132 28532 27188 28542
rect 27132 28438 27188 28476
rect 27132 28084 27188 28094
rect 27132 27970 27188 28028
rect 27132 27918 27134 27970
rect 27186 27918 27188 27970
rect 27132 27906 27188 27918
rect 27020 27636 27076 27646
rect 27020 27186 27076 27580
rect 27020 27134 27022 27186
rect 27074 27134 27076 27186
rect 27020 27122 27076 27134
rect 27244 26908 27300 31892
rect 27132 26852 27300 26908
rect 27132 25620 27188 26852
rect 27244 26740 27300 26750
rect 27244 26514 27300 26684
rect 27244 26462 27246 26514
rect 27298 26462 27300 26514
rect 27244 26450 27300 26462
rect 27132 25554 27188 25564
rect 27244 25844 27300 25854
rect 27132 25396 27188 25406
rect 27132 24834 27188 25340
rect 27244 25394 27300 25788
rect 27244 25342 27246 25394
rect 27298 25342 27300 25394
rect 27244 25330 27300 25342
rect 27132 24782 27134 24834
rect 27186 24782 27188 24834
rect 27132 24770 27188 24782
rect 27356 24612 27412 37772
rect 27468 32340 27524 41132
rect 27468 32274 27524 32284
rect 27356 24546 27412 24556
rect 27468 31780 27524 31790
rect 27244 24500 27300 24510
rect 27244 23826 27300 24444
rect 27244 23774 27246 23826
rect 27298 23774 27300 23826
rect 27244 23762 27300 23774
rect 27132 23604 27188 23614
rect 27132 23266 27188 23548
rect 27132 23214 27134 23266
rect 27186 23214 27188 23266
rect 27132 23202 27188 23214
rect 27244 22708 27300 22718
rect 27132 22260 27188 22270
rect 27132 21698 27188 22204
rect 27244 22258 27300 22652
rect 27244 22206 27246 22258
rect 27298 22206 27300 22258
rect 27244 22194 27300 22206
rect 27132 21646 27134 21698
rect 27186 21646 27188 21698
rect 27132 21634 27188 21646
rect 27468 21588 27524 31724
rect 27244 21532 27524 21588
rect 27692 30996 27748 31006
rect 26908 20972 27188 21028
rect 26684 20850 26740 20860
rect 26908 20804 26964 20814
rect 26908 20710 26964 20748
rect 26572 20468 26628 20478
rect 26572 20018 26628 20412
rect 26572 19966 26574 20018
rect 26626 19966 26628 20018
rect 26572 19954 26628 19966
rect 26796 20244 26852 20254
rect 26460 19348 26516 19358
rect 26460 19254 26516 19292
rect 26796 18788 26852 20188
rect 26908 19908 26964 19918
rect 26908 19814 26964 19852
rect 26908 19122 26964 19134
rect 26908 19070 26910 19122
rect 26962 19070 26964 19122
rect 26908 19012 26964 19070
rect 26908 18946 26964 18956
rect 26796 18732 27076 18788
rect 26572 18452 26628 18462
rect 26572 18358 26628 18396
rect 26908 18340 26964 18350
rect 26908 18246 26964 18284
rect 26908 17892 26964 17902
rect 26572 17780 26628 17790
rect 26572 17686 26628 17724
rect 26908 17778 26964 17836
rect 26908 17726 26910 17778
rect 26962 17726 26964 17778
rect 26908 17714 26964 17726
rect 26908 17556 26964 17566
rect 26572 16884 26628 16894
rect 26572 16790 26628 16828
rect 26908 16772 26964 17500
rect 27020 16994 27076 18732
rect 27020 16942 27022 16994
rect 27074 16942 27076 16994
rect 27020 16930 27076 16942
rect 26908 16716 27076 16772
rect 26908 16212 26964 16222
rect 26908 16118 26964 16156
rect 26572 16098 26628 16110
rect 26572 16046 26574 16098
rect 26626 16046 26628 16098
rect 26572 15988 26628 16046
rect 26572 15922 26628 15932
rect 26908 15540 26964 15550
rect 26684 15428 26740 15438
rect 26572 15092 26628 15102
rect 26572 14998 26628 15036
rect 26348 14466 26404 14476
rect 26348 14308 26404 14318
rect 26348 14214 26404 14252
rect 26012 13806 26014 13858
rect 26066 13806 26068 13858
rect 26012 13794 26068 13806
rect 26572 13748 26628 13758
rect 26572 13654 26628 13692
rect 26572 13524 26628 13534
rect 26460 13468 26572 13524
rect 26012 12850 26068 12862
rect 26012 12798 26014 12850
rect 26066 12798 26068 12850
rect 26012 12404 26068 12798
rect 26012 12338 26068 12348
rect 26012 12180 26068 12190
rect 26012 12086 26068 12124
rect 25900 11732 25956 11742
rect 25900 10724 25956 11676
rect 26012 11620 26068 11630
rect 26012 11506 26068 11564
rect 26012 11454 26014 11506
rect 26066 11454 26068 11506
rect 26012 11442 26068 11454
rect 26236 11284 26292 11294
rect 26012 10724 26068 10734
rect 25900 10722 26068 10724
rect 25900 10670 26014 10722
rect 26066 10670 26068 10722
rect 25900 10668 26068 10670
rect 26012 10658 26068 10668
rect 26012 9714 26068 9726
rect 26012 9662 26014 9714
rect 26066 9662 26068 9714
rect 26012 9156 26068 9662
rect 26012 9090 26068 9100
rect 25900 8820 25956 8830
rect 25900 8726 25956 8764
rect 26012 8484 26068 8494
rect 26012 7586 26068 8428
rect 26012 7534 26014 7586
rect 26066 7534 26068 7586
rect 26012 7522 26068 7534
rect 26124 7476 26180 7486
rect 26012 6804 26068 6814
rect 26012 6710 26068 6748
rect 25900 5684 25956 5694
rect 25900 5590 25956 5628
rect 26124 3442 26180 7420
rect 26236 6132 26292 11228
rect 26348 9940 26404 9950
rect 26348 9268 26404 9884
rect 26460 9492 26516 13468
rect 26572 13458 26628 13468
rect 26572 12962 26628 12974
rect 26572 12910 26574 12962
rect 26626 12910 26628 12962
rect 26572 12852 26628 12910
rect 26572 12786 26628 12796
rect 26572 11956 26628 11966
rect 26572 11862 26628 11900
rect 26572 11394 26628 11406
rect 26572 11342 26574 11394
rect 26626 11342 26628 11394
rect 26572 11060 26628 11342
rect 26572 10994 26628 11004
rect 26572 10386 26628 10398
rect 26572 10334 26574 10386
rect 26626 10334 26628 10386
rect 26572 10164 26628 10334
rect 26572 10098 26628 10108
rect 26572 9826 26628 9838
rect 26572 9774 26574 9826
rect 26626 9774 26628 9826
rect 26572 9716 26628 9774
rect 26572 9650 26628 9660
rect 26460 9436 26628 9492
rect 26460 9268 26516 9278
rect 26348 9266 26516 9268
rect 26348 9214 26462 9266
rect 26514 9214 26516 9266
rect 26348 9212 26516 9214
rect 26460 9202 26516 9212
rect 26460 9044 26516 9054
rect 26460 8146 26516 8988
rect 26460 8094 26462 8146
rect 26514 8094 26516 8146
rect 26460 8082 26516 8094
rect 26572 7924 26628 9436
rect 26460 7868 26628 7924
rect 26460 6356 26516 7868
rect 26684 7476 26740 15372
rect 26908 15426 26964 15484
rect 26908 15374 26910 15426
rect 26962 15374 26964 15426
rect 26908 15362 26964 15374
rect 27020 15148 27076 16716
rect 26908 15092 27076 15148
rect 26908 14642 26964 15092
rect 26908 14590 26910 14642
rect 26962 14590 26964 14642
rect 26908 14578 26964 14590
rect 27020 14532 27076 14542
rect 27020 14084 27076 14476
rect 26908 14028 27076 14084
rect 26908 12628 26964 14028
rect 27020 13860 27076 13870
rect 27020 13766 27076 13804
rect 27020 12852 27076 12862
rect 27132 12852 27188 20972
rect 27020 12850 27188 12852
rect 27020 12798 27022 12850
rect 27074 12798 27188 12850
rect 27020 12796 27188 12798
rect 27020 12786 27076 12796
rect 27132 12628 27188 12638
rect 26908 12572 27076 12628
rect 26908 12068 26964 12078
rect 26908 11974 26964 12012
rect 26908 11508 26964 11518
rect 26908 11414 26964 11452
rect 26908 10948 26964 10958
rect 26908 9938 26964 10892
rect 27020 10722 27076 12572
rect 27020 10670 27022 10722
rect 27074 10670 27076 10722
rect 27020 10658 27076 10670
rect 26908 9886 26910 9938
rect 26962 9886 26964 9938
rect 26908 9874 26964 9886
rect 26684 7410 26740 7420
rect 26908 7700 26964 7710
rect 26572 7252 26628 7262
rect 26572 7250 26740 7252
rect 26572 7198 26574 7250
rect 26626 7198 26740 7250
rect 26572 7196 26740 7198
rect 26572 7186 26628 7196
rect 26572 6690 26628 6702
rect 26572 6638 26574 6690
rect 26626 6638 26628 6690
rect 26572 6580 26628 6638
rect 26572 6514 26628 6524
rect 26460 6300 26628 6356
rect 26460 6132 26516 6142
rect 26236 6130 26516 6132
rect 26236 6078 26462 6130
rect 26514 6078 26516 6130
rect 26236 6076 26516 6078
rect 26460 6066 26516 6076
rect 26572 5908 26628 6300
rect 26684 6132 26740 7196
rect 26908 6802 26964 7644
rect 27020 7588 27076 7598
rect 27020 7494 27076 7532
rect 26908 6750 26910 6802
rect 26962 6750 26964 6802
rect 26908 6738 26964 6750
rect 26684 6066 26740 6076
rect 26124 3390 26126 3442
rect 26178 3390 26180 3442
rect 25788 3332 26068 3388
rect 26124 3378 26180 3390
rect 26460 5852 26628 5908
rect 25228 2830 25230 2882
rect 25282 2830 25284 2882
rect 25228 2818 25284 2830
rect 25564 2772 25620 2782
rect 25564 2212 25620 2716
rect 26012 2660 26068 3332
rect 26460 3220 26516 5852
rect 26684 5236 26740 5246
rect 26684 5142 26740 5180
rect 26908 4228 26964 4238
rect 26908 4134 26964 4172
rect 26908 3668 26964 3678
rect 26908 3574 26964 3612
rect 26124 3164 26516 3220
rect 26572 3554 26628 3566
rect 26572 3502 26574 3554
rect 26626 3502 26628 3554
rect 26124 2882 26180 3164
rect 26572 2996 26628 3502
rect 26572 2930 26628 2940
rect 26124 2830 26126 2882
rect 26178 2830 26180 2882
rect 26124 2818 26180 2830
rect 27020 2884 27076 2894
rect 27132 2884 27188 12572
rect 27244 9380 27300 21532
rect 27468 21364 27524 21374
rect 27356 20916 27412 20926
rect 27356 20822 27412 20860
rect 27468 20018 27524 21308
rect 27468 19966 27470 20018
rect 27522 19966 27524 20018
rect 27468 19954 27524 19966
rect 27580 20916 27636 20926
rect 27356 19572 27412 19582
rect 27356 18450 27412 19516
rect 27468 19460 27524 19470
rect 27580 19460 27636 20860
rect 27468 19458 27636 19460
rect 27468 19406 27470 19458
rect 27522 19406 27636 19458
rect 27468 19404 27636 19406
rect 27468 19394 27524 19404
rect 27356 18398 27358 18450
rect 27410 18398 27412 18450
rect 27356 18386 27412 18398
rect 27580 19124 27636 19134
rect 27356 18228 27412 18238
rect 27356 16882 27412 18172
rect 27468 17892 27524 17902
rect 27580 17892 27636 19068
rect 27692 18340 27748 30940
rect 27692 18274 27748 18284
rect 27804 25620 27860 25630
rect 27468 17890 27636 17892
rect 27468 17838 27470 17890
rect 27522 17838 27636 17890
rect 27468 17836 27636 17838
rect 27468 17826 27524 17836
rect 27356 16830 27358 16882
rect 27410 16830 27412 16882
rect 27356 16818 27412 16830
rect 27580 17332 27636 17342
rect 27356 16436 27412 16446
rect 27356 15314 27412 16380
rect 27468 16324 27524 16334
rect 27580 16324 27636 17276
rect 27468 16322 27636 16324
rect 27468 16270 27470 16322
rect 27522 16270 27636 16322
rect 27468 16268 27636 16270
rect 27468 16258 27524 16268
rect 27356 15262 27358 15314
rect 27410 15262 27412 15314
rect 27356 15250 27412 15262
rect 27580 15540 27636 15550
rect 27468 14756 27524 14766
rect 27580 14756 27636 15484
rect 27468 14754 27636 14756
rect 27468 14702 27470 14754
rect 27522 14702 27636 14754
rect 27468 14700 27636 14702
rect 27692 15316 27748 15326
rect 27468 14690 27524 14700
rect 27356 14644 27412 14654
rect 27356 13746 27412 14588
rect 27356 13694 27358 13746
rect 27410 13694 27412 13746
rect 27356 13682 27412 13694
rect 27468 14196 27524 14206
rect 27356 13300 27412 13310
rect 27356 12178 27412 13244
rect 27468 13186 27524 14140
rect 27468 13134 27470 13186
rect 27522 13134 27524 13186
rect 27468 13122 27524 13134
rect 27468 12964 27524 12974
rect 27468 12292 27524 12908
rect 27468 12226 27524 12236
rect 27580 12404 27636 12414
rect 27356 12126 27358 12178
rect 27410 12126 27412 12178
rect 27356 12114 27412 12126
rect 27468 11620 27524 11630
rect 27580 11620 27636 12348
rect 27468 11618 27636 11620
rect 27468 11566 27470 11618
rect 27522 11566 27636 11618
rect 27468 11564 27636 11566
rect 27468 11554 27524 11564
rect 27356 11508 27412 11518
rect 27356 10610 27412 11452
rect 27692 10948 27748 15260
rect 27692 10882 27748 10892
rect 27356 10558 27358 10610
rect 27410 10558 27412 10610
rect 27356 10546 27412 10558
rect 27580 10612 27636 10622
rect 27468 10052 27524 10062
rect 27580 10052 27636 10556
rect 27468 10050 27636 10052
rect 27468 9998 27470 10050
rect 27522 9998 27636 10050
rect 27468 9996 27636 9998
rect 27468 9986 27524 9996
rect 27804 9940 27860 25564
rect 28028 23716 28084 23726
rect 27580 9884 27860 9940
rect 27916 20804 27972 20814
rect 27244 9314 27300 9324
rect 27468 9604 27524 9614
rect 27244 9042 27300 9054
rect 27244 8990 27246 9042
rect 27298 8990 27300 9042
rect 27244 8372 27300 8990
rect 27244 8306 27300 8316
rect 27356 8258 27412 8270
rect 27356 8206 27358 8258
rect 27410 8206 27412 8258
rect 27244 8148 27300 8158
rect 27244 4340 27300 8092
rect 27356 7476 27412 8206
rect 27468 7812 27524 9548
rect 27580 8260 27636 9884
rect 27580 8194 27636 8204
rect 27692 9380 27748 9390
rect 27468 7756 27636 7812
rect 27356 7410 27412 7420
rect 27468 7364 27524 7374
rect 27468 7270 27524 7308
rect 27468 7028 27524 7038
rect 27468 6914 27524 6972
rect 27468 6862 27470 6914
rect 27522 6862 27524 6914
rect 27468 6850 27524 6862
rect 27356 5906 27412 5918
rect 27356 5854 27358 5906
rect 27410 5854 27412 5906
rect 27356 5236 27412 5854
rect 27356 5170 27412 5180
rect 27468 5122 27524 5134
rect 27468 5070 27470 5122
rect 27522 5070 27524 5122
rect 27468 4788 27524 5070
rect 27468 4722 27524 4732
rect 27244 4274 27300 4284
rect 27468 4340 27524 4350
rect 27468 4246 27524 4284
rect 27468 3892 27524 3902
rect 27468 3778 27524 3836
rect 27468 3726 27470 3778
rect 27522 3726 27524 3778
rect 27468 3714 27524 3726
rect 27580 3668 27636 7756
rect 27692 5348 27748 9324
rect 27916 8428 27972 20748
rect 28028 16212 28084 23660
rect 28252 20580 28308 20590
rect 28028 16146 28084 16156
rect 28140 16996 28196 17006
rect 28028 15876 28084 15886
rect 28028 12628 28084 15820
rect 28028 12562 28084 12572
rect 27692 5282 27748 5292
rect 27804 8372 27972 8428
rect 28028 12292 28084 12302
rect 28028 8428 28084 12236
rect 28140 9604 28196 16940
rect 28140 9538 28196 9548
rect 28028 8372 28196 8428
rect 27804 4900 27860 8372
rect 28140 7588 28196 8372
rect 28140 7522 28196 7532
rect 27804 4834 27860 4844
rect 28252 4564 28308 20524
rect 28252 4498 28308 4508
rect 27580 3602 27636 3612
rect 27692 4452 27748 4462
rect 27020 2882 27188 2884
rect 27020 2830 27022 2882
rect 27074 2830 27188 2882
rect 27020 2828 27188 2830
rect 27468 3444 27524 3454
rect 27020 2818 27076 2828
rect 27468 2770 27524 3388
rect 27468 2718 27470 2770
rect 27522 2718 27524 2770
rect 27468 2706 27524 2718
rect 26012 2604 26516 2660
rect 25676 2548 25732 2558
rect 25676 2546 25844 2548
rect 25676 2494 25678 2546
rect 25730 2494 25844 2546
rect 25676 2492 25844 2494
rect 25676 2482 25732 2492
rect 25564 2156 25732 2212
rect 25564 1986 25620 1998
rect 25564 1934 25566 1986
rect 25618 1934 25620 1986
rect 25228 1876 25284 1886
rect 25228 1782 25284 1820
rect 24892 1262 24894 1314
rect 24946 1262 24948 1314
rect 24892 1250 24948 1262
rect 25564 1204 25620 1934
rect 25676 1314 25732 2156
rect 25788 2100 25844 2492
rect 25788 2034 25844 2044
rect 25676 1262 25678 1314
rect 25730 1262 25732 1314
rect 25676 1250 25732 1262
rect 26012 1986 26068 1998
rect 26012 1934 26014 1986
rect 26066 1934 26068 1986
rect 26012 1316 26068 1934
rect 26460 1874 26516 2604
rect 26572 2548 26628 2558
rect 26572 2454 26628 2492
rect 27468 2212 27524 2222
rect 27692 2212 27748 4396
rect 27468 2098 27524 2156
rect 27468 2046 27470 2098
rect 27522 2046 27524 2098
rect 27468 2034 27524 2046
rect 27580 2156 27748 2212
rect 26460 1822 26462 1874
rect 26514 1822 26516 1874
rect 26460 1810 26516 1822
rect 26908 1986 26964 1998
rect 26908 1934 26910 1986
rect 26962 1934 26964 1986
rect 26012 1250 26068 1260
rect 26572 1428 26628 1438
rect 26572 1314 26628 1372
rect 26572 1262 26574 1314
rect 26626 1262 26628 1314
rect 26572 1250 26628 1262
rect 25564 1138 25620 1148
rect 23548 1092 23604 1102
rect 23548 112 23604 1036
rect 25340 978 25396 990
rect 25340 926 25342 978
rect 25394 926 25396 978
rect 24464 812 24728 822
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24464 746 24728 756
rect 25340 756 25396 926
rect 26236 980 26292 990
rect 26236 978 26404 980
rect 26236 926 26238 978
rect 26290 926 26404 978
rect 26236 924 26404 926
rect 26236 914 26292 924
rect 25340 690 25396 700
rect 26236 644 26292 654
rect 24892 420 24948 430
rect 24892 112 24948 364
rect 26236 112 26292 588
rect 26348 308 26404 924
rect 26348 242 26404 252
rect 26908 196 26964 1934
rect 27132 1652 27188 1662
rect 27132 1202 27188 1596
rect 27132 1150 27134 1202
rect 27186 1150 27188 1202
rect 27132 1138 27188 1150
rect 26908 130 26964 140
rect 27580 112 27636 2156
rect 672 0 784 112
rect 2016 0 2128 112
rect 3360 0 3472 112
rect 4704 0 4816 112
rect 6048 0 6160 112
rect 7392 0 7504 112
rect 8736 0 8848 112
rect 10080 0 10192 112
rect 11424 0 11536 112
rect 12768 0 12880 112
rect 14112 0 14224 112
rect 15456 0 15568 112
rect 16800 0 16912 112
rect 18144 0 18256 112
rect 19488 0 19600 112
rect 20832 0 20944 112
rect 22176 0 22288 112
rect 23520 0 23632 112
rect 24864 0 24976 112
rect 26208 0 26320 112
rect 27552 0 27664 112
<< via2 >>
rect 3804 56474 3860 56476
rect 3804 56422 3806 56474
rect 3806 56422 3858 56474
rect 3858 56422 3860 56474
rect 3804 56420 3860 56422
rect 3908 56474 3964 56476
rect 3908 56422 3910 56474
rect 3910 56422 3962 56474
rect 3962 56422 3964 56474
rect 3908 56420 3964 56422
rect 4012 56474 4068 56476
rect 4012 56422 4014 56474
rect 4014 56422 4066 56474
rect 4066 56422 4068 56474
rect 4012 56420 4068 56422
rect 3052 55970 3108 55972
rect 3052 55918 3054 55970
rect 3054 55918 3106 55970
rect 3106 55918 3108 55970
rect 3052 55916 3108 55918
rect 4464 55690 4520 55692
rect 4464 55638 4466 55690
rect 4466 55638 4518 55690
rect 4518 55638 4520 55690
rect 4464 55636 4520 55638
rect 4568 55690 4624 55692
rect 4568 55638 4570 55690
rect 4570 55638 4622 55690
rect 4622 55638 4624 55690
rect 4568 55636 4624 55638
rect 4672 55690 4728 55692
rect 4672 55638 4674 55690
rect 4674 55638 4726 55690
rect 4726 55638 4728 55690
rect 4672 55636 4728 55638
rect 1372 55244 1428 55300
rect 1036 55132 1092 55188
rect 1036 54290 1092 54292
rect 1036 54238 1038 54290
rect 1038 54238 1090 54290
rect 1090 54238 1092 54290
rect 1036 54236 1092 54238
rect 1036 53340 1092 53396
rect 1036 52444 1092 52500
rect 1036 51548 1092 51604
rect 924 50652 980 50708
rect 1036 49756 1092 49812
rect 1036 48860 1092 48916
rect 1148 48412 1204 48468
rect 812 48076 868 48132
rect 1036 48018 1092 48020
rect 1036 47966 1038 48018
rect 1038 47966 1090 48018
rect 1090 47966 1092 48018
rect 1036 47964 1092 47966
rect 1036 47068 1092 47124
rect 924 45276 980 45332
rect 812 43596 868 43652
rect 1148 44380 1204 44436
rect 924 43484 980 43540
rect 252 41020 308 41076
rect 364 39004 420 39060
rect 1148 42588 1204 42644
rect 476 37212 532 37268
rect 364 36764 420 36820
rect 588 36316 644 36372
rect 700 40236 756 40292
rect 364 35420 420 35476
rect 588 35756 644 35812
rect 140 30716 196 30772
rect 364 30716 420 30772
rect 140 27356 196 27412
rect 140 27020 196 27076
rect 588 33292 644 33348
rect 476 26348 532 26404
rect 588 33068 644 33124
rect 364 22092 420 22148
rect 364 20636 420 20692
rect 812 36764 868 36820
rect 1596 52162 1652 52164
rect 1596 52110 1598 52162
rect 1598 52110 1650 52162
rect 1650 52110 1652 52162
rect 1596 52108 1652 52110
rect 1596 51266 1652 51268
rect 1596 51214 1598 51266
rect 1598 51214 1650 51266
rect 1650 51214 1652 51266
rect 1596 51212 1652 51214
rect 1596 50482 1652 50484
rect 1596 50430 1598 50482
rect 1598 50430 1650 50482
rect 1650 50430 1652 50482
rect 1596 50428 1652 50430
rect 2380 50428 2436 50484
rect 1596 48130 1652 48132
rect 1596 48078 1598 48130
rect 1598 48078 1650 48130
rect 1650 48078 1652 48130
rect 1596 48076 1652 48078
rect 1596 46562 1652 46564
rect 1596 46510 1598 46562
rect 1598 46510 1650 46562
rect 1650 46510 1652 46562
rect 1596 46508 1652 46510
rect 1484 46284 1540 46340
rect 1596 45778 1652 45780
rect 1596 45726 1598 45778
rect 1598 45726 1650 45778
rect 1650 45726 1652 45778
rect 1596 45724 1652 45726
rect 1596 44380 1652 44436
rect 1596 43708 1652 43764
rect 1596 43426 1652 43428
rect 1596 43374 1598 43426
rect 1598 43374 1650 43426
rect 1650 43374 1652 43426
rect 1596 43372 1652 43374
rect 1932 46172 1988 46228
rect 1708 42812 1764 42868
rect 1596 42140 1652 42196
rect 1708 42588 1764 42644
rect 1372 42028 1428 42084
rect 1596 41858 1652 41860
rect 1596 41806 1598 41858
rect 1598 41806 1650 41858
rect 1650 41806 1652 41858
rect 1596 41804 1652 41806
rect 1596 41074 1652 41076
rect 1596 41022 1598 41074
rect 1598 41022 1650 41074
rect 1650 41022 1652 41074
rect 1596 41020 1652 41022
rect 1372 40572 1428 40628
rect 2380 42924 2436 42980
rect 2604 43372 2660 43428
rect 2380 42642 2436 42644
rect 2380 42590 2382 42642
rect 2382 42590 2434 42642
rect 2434 42590 2436 42642
rect 2380 42588 2436 42590
rect 2044 42140 2100 42196
rect 1932 41746 1988 41748
rect 1932 41694 1934 41746
rect 1934 41694 1986 41746
rect 1986 41694 1988 41746
rect 1932 41692 1988 41694
rect 1820 40796 1876 40852
rect 2268 41580 2324 41636
rect 1596 40290 1652 40292
rect 1596 40238 1598 40290
rect 1598 40238 1650 40290
rect 1650 40238 1652 40290
rect 1596 40236 1652 40238
rect 1596 38946 1652 38948
rect 1596 38894 1598 38946
rect 1598 38894 1650 38946
rect 1650 38894 1652 38946
rect 1596 38892 1652 38894
rect 1708 38556 1764 38612
rect 1820 37996 1876 38052
rect 2044 39900 2100 39956
rect 2156 40236 2212 40292
rect 2268 39788 2324 39844
rect 2156 38556 2212 38612
rect 1932 37884 1988 37940
rect 1708 37100 1764 37156
rect 1372 35756 1428 35812
rect 1708 36876 1764 36932
rect 1260 35644 1316 35700
rect 812 33628 868 33684
rect 1372 35084 1428 35140
rect 1148 34524 1204 34580
rect 1260 34972 1316 35028
rect 1596 34802 1652 34804
rect 1596 34750 1598 34802
rect 1598 34750 1650 34802
rect 1650 34750 1652 34802
rect 1596 34748 1652 34750
rect 1596 34412 1652 34468
rect 1484 34130 1540 34132
rect 1484 34078 1486 34130
rect 1486 34078 1538 34130
rect 1538 34078 1540 34130
rect 1484 34076 1540 34078
rect 1260 33628 1316 33684
rect 1484 33628 1540 33684
rect 1148 33516 1204 33572
rect 924 31836 980 31892
rect 1148 33292 1204 33348
rect 1148 32284 1204 32340
rect 1148 31724 1204 31780
rect 1260 32396 1316 32452
rect 1036 30940 1092 30996
rect 1932 35196 1988 35252
rect 1708 33628 1764 33684
rect 1596 33234 1652 33236
rect 1596 33182 1598 33234
rect 1598 33182 1650 33234
rect 1650 33182 1652 33234
rect 1596 33180 1652 33182
rect 2268 36652 2324 36708
rect 2156 36370 2212 36372
rect 2156 36318 2158 36370
rect 2158 36318 2210 36370
rect 2210 36318 2212 36370
rect 2156 36316 2212 36318
rect 2268 35586 2324 35588
rect 2268 35534 2270 35586
rect 2270 35534 2322 35586
rect 2322 35534 2324 35586
rect 2268 35532 2324 35534
rect 2156 35420 2212 35476
rect 2268 35196 2324 35252
rect 2268 34412 2324 34468
rect 1932 33852 1988 33908
rect 1820 32732 1876 32788
rect 2044 33628 2100 33684
rect 1708 32450 1764 32452
rect 1708 32398 1710 32450
rect 1710 32398 1762 32450
rect 1762 32398 1764 32450
rect 1708 32396 1764 32398
rect 2044 31890 2100 31892
rect 2044 31838 2046 31890
rect 2046 31838 2098 31890
rect 2098 31838 2100 31890
rect 2044 31836 2100 31838
rect 1708 31778 1764 31780
rect 1708 31726 1710 31778
rect 1710 31726 1762 31778
rect 1762 31726 1764 31778
rect 1708 31724 1764 31726
rect 1260 30268 1316 30324
rect 1036 30044 1092 30100
rect 1036 29202 1092 29204
rect 1036 29150 1038 29202
rect 1038 29150 1090 29202
rect 1090 29150 1092 29202
rect 1036 29148 1092 29150
rect 1036 28924 1092 28980
rect 1932 30044 1988 30100
rect 1484 28476 1540 28532
rect 588 13132 644 13188
rect 700 23884 756 23940
rect 812 18620 868 18676
rect 812 18396 868 18452
rect 812 9212 868 9268
rect 700 5516 756 5572
rect 364 2828 420 2884
rect 1036 27020 1092 27076
rect 1260 27074 1316 27076
rect 1260 27022 1262 27074
rect 1262 27022 1314 27074
rect 1314 27022 1316 27074
rect 1260 27020 1316 27022
rect 1708 27298 1764 27300
rect 1708 27246 1710 27298
rect 1710 27246 1762 27298
rect 1762 27246 1764 27298
rect 1708 27244 1764 27246
rect 1260 26460 1316 26516
rect 1372 24892 1428 24948
rect 1036 23772 1092 23828
rect 1148 22316 1204 22372
rect 1260 22258 1316 22260
rect 1260 22206 1262 22258
rect 1262 22206 1314 22258
rect 1314 22206 1316 22258
rect 1260 22204 1316 22206
rect 1596 24108 1652 24164
rect 1484 23212 1540 23268
rect 1596 23548 1652 23604
rect 1820 27020 1876 27076
rect 1820 25452 1876 25508
rect 2044 28530 2100 28532
rect 2044 28478 2046 28530
rect 2046 28478 2098 28530
rect 2098 28478 2100 28530
rect 2044 28476 2100 28478
rect 2268 33516 2324 33572
rect 2268 30210 2324 30212
rect 2268 30158 2270 30210
rect 2270 30158 2322 30210
rect 2322 30158 2324 30210
rect 2268 30156 2324 30158
rect 2492 40514 2548 40516
rect 2492 40462 2494 40514
rect 2494 40462 2546 40514
rect 2546 40462 2548 40514
rect 2492 40460 2548 40462
rect 2492 39842 2548 39844
rect 2492 39790 2494 39842
rect 2494 39790 2546 39842
rect 2546 39790 2548 39842
rect 2492 39788 2548 39790
rect 2492 37996 2548 38052
rect 2716 38444 2772 38500
rect 3052 41916 3108 41972
rect 2828 38108 2884 38164
rect 2828 37884 2884 37940
rect 2716 37378 2772 37380
rect 2716 37326 2718 37378
rect 2718 37326 2770 37378
rect 2770 37326 2772 37378
rect 2716 37324 2772 37326
rect 2604 36652 2660 36708
rect 2716 35810 2772 35812
rect 2716 35758 2718 35810
rect 2718 35758 2770 35810
rect 2770 35758 2772 35810
rect 2716 35756 2772 35758
rect 2604 35308 2660 35364
rect 2828 35196 2884 35252
rect 2492 34188 2548 34244
rect 2492 33964 2548 34020
rect 3052 36540 3108 36596
rect 3164 36428 3220 36484
rect 3164 35644 3220 35700
rect 2716 33516 2772 33572
rect 6188 55804 6244 55860
rect 6076 55132 6132 55188
rect 3804 54906 3860 54908
rect 3804 54854 3806 54906
rect 3806 54854 3858 54906
rect 3858 54854 3860 54906
rect 3804 54852 3860 54854
rect 3908 54906 3964 54908
rect 3908 54854 3910 54906
rect 3910 54854 3962 54906
rect 3962 54854 3964 54906
rect 3908 54852 3964 54854
rect 4012 54906 4068 54908
rect 4012 54854 4014 54906
rect 4014 54854 4066 54906
rect 4066 54854 4068 54906
rect 4012 54852 4068 54854
rect 4464 54122 4520 54124
rect 4464 54070 4466 54122
rect 4466 54070 4518 54122
rect 4518 54070 4520 54122
rect 4464 54068 4520 54070
rect 4568 54122 4624 54124
rect 4568 54070 4570 54122
rect 4570 54070 4622 54122
rect 4622 54070 4624 54122
rect 4568 54068 4624 54070
rect 4672 54122 4728 54124
rect 4672 54070 4674 54122
rect 4674 54070 4726 54122
rect 4726 54070 4728 54122
rect 4672 54068 4728 54070
rect 3804 53338 3860 53340
rect 3804 53286 3806 53338
rect 3806 53286 3858 53338
rect 3858 53286 3860 53338
rect 3804 53284 3860 53286
rect 3908 53338 3964 53340
rect 3908 53286 3910 53338
rect 3910 53286 3962 53338
rect 3962 53286 3964 53338
rect 3908 53284 3964 53286
rect 4012 53338 4068 53340
rect 4012 53286 4014 53338
rect 4014 53286 4066 53338
rect 4066 53286 4068 53338
rect 4012 53284 4068 53286
rect 4464 52554 4520 52556
rect 4464 52502 4466 52554
rect 4466 52502 4518 52554
rect 4518 52502 4520 52554
rect 4464 52500 4520 52502
rect 4568 52554 4624 52556
rect 4568 52502 4570 52554
rect 4570 52502 4622 52554
rect 4622 52502 4624 52554
rect 4568 52500 4624 52502
rect 4672 52554 4728 52556
rect 4672 52502 4674 52554
rect 4674 52502 4726 52554
rect 4726 52502 4728 52554
rect 4672 52500 4728 52502
rect 3804 51770 3860 51772
rect 3804 51718 3806 51770
rect 3806 51718 3858 51770
rect 3858 51718 3860 51770
rect 3804 51716 3860 51718
rect 3908 51770 3964 51772
rect 3908 51718 3910 51770
rect 3910 51718 3962 51770
rect 3962 51718 3964 51770
rect 3908 51716 3964 51718
rect 4012 51770 4068 51772
rect 4012 51718 4014 51770
rect 4014 51718 4066 51770
rect 4066 51718 4068 51770
rect 4012 51716 4068 51718
rect 5852 51212 5908 51268
rect 4464 50986 4520 50988
rect 4464 50934 4466 50986
rect 4466 50934 4518 50986
rect 4518 50934 4520 50986
rect 4464 50932 4520 50934
rect 4568 50986 4624 50988
rect 4568 50934 4570 50986
rect 4570 50934 4622 50986
rect 4622 50934 4624 50986
rect 4568 50932 4624 50934
rect 4672 50986 4728 50988
rect 4672 50934 4674 50986
rect 4674 50934 4726 50986
rect 4726 50934 4728 50986
rect 4672 50932 4728 50934
rect 3804 50202 3860 50204
rect 3804 50150 3806 50202
rect 3806 50150 3858 50202
rect 3858 50150 3860 50202
rect 3804 50148 3860 50150
rect 3908 50202 3964 50204
rect 3908 50150 3910 50202
rect 3910 50150 3962 50202
rect 3962 50150 3964 50202
rect 3908 50148 3964 50150
rect 4012 50202 4068 50204
rect 4012 50150 4014 50202
rect 4014 50150 4066 50202
rect 4066 50150 4068 50202
rect 4012 50148 4068 50150
rect 4464 49418 4520 49420
rect 4464 49366 4466 49418
rect 4466 49366 4518 49418
rect 4518 49366 4520 49418
rect 4464 49364 4520 49366
rect 4568 49418 4624 49420
rect 4568 49366 4570 49418
rect 4570 49366 4622 49418
rect 4622 49366 4624 49418
rect 4568 49364 4624 49366
rect 4672 49418 4728 49420
rect 4672 49366 4674 49418
rect 4674 49366 4726 49418
rect 4726 49366 4728 49418
rect 4672 49364 4728 49366
rect 3804 48634 3860 48636
rect 3804 48582 3806 48634
rect 3806 48582 3858 48634
rect 3858 48582 3860 48634
rect 3804 48580 3860 48582
rect 3908 48634 3964 48636
rect 3908 48582 3910 48634
rect 3910 48582 3962 48634
rect 3962 48582 3964 48634
rect 3908 48580 3964 48582
rect 4012 48634 4068 48636
rect 4012 48582 4014 48634
rect 4014 48582 4066 48634
rect 4066 48582 4068 48634
rect 4012 48580 4068 48582
rect 5628 48412 5684 48468
rect 4464 47850 4520 47852
rect 4464 47798 4466 47850
rect 4466 47798 4518 47850
rect 4518 47798 4520 47850
rect 4464 47796 4520 47798
rect 4568 47850 4624 47852
rect 4568 47798 4570 47850
rect 4570 47798 4622 47850
rect 4622 47798 4624 47850
rect 4568 47796 4624 47798
rect 4672 47850 4728 47852
rect 4672 47798 4674 47850
rect 4674 47798 4726 47850
rect 4726 47798 4728 47850
rect 4672 47796 4728 47798
rect 3804 47066 3860 47068
rect 3804 47014 3806 47066
rect 3806 47014 3858 47066
rect 3858 47014 3860 47066
rect 3804 47012 3860 47014
rect 3908 47066 3964 47068
rect 3908 47014 3910 47066
rect 3910 47014 3962 47066
rect 3962 47014 3964 47066
rect 3908 47012 3964 47014
rect 4012 47066 4068 47068
rect 4012 47014 4014 47066
rect 4014 47014 4066 47066
rect 4066 47014 4068 47066
rect 4012 47012 4068 47014
rect 4464 46282 4520 46284
rect 4464 46230 4466 46282
rect 4466 46230 4518 46282
rect 4518 46230 4520 46282
rect 4464 46228 4520 46230
rect 4568 46282 4624 46284
rect 4568 46230 4570 46282
rect 4570 46230 4622 46282
rect 4622 46230 4624 46282
rect 4568 46228 4624 46230
rect 4672 46282 4728 46284
rect 4672 46230 4674 46282
rect 4674 46230 4726 46282
rect 4726 46230 4728 46282
rect 4672 46228 4728 46230
rect 3804 45498 3860 45500
rect 3804 45446 3806 45498
rect 3806 45446 3858 45498
rect 3858 45446 3860 45498
rect 3804 45444 3860 45446
rect 3908 45498 3964 45500
rect 3908 45446 3910 45498
rect 3910 45446 3962 45498
rect 3962 45446 3964 45498
rect 3908 45444 3964 45446
rect 4012 45498 4068 45500
rect 4012 45446 4014 45498
rect 4014 45446 4066 45498
rect 4066 45446 4068 45498
rect 4012 45444 4068 45446
rect 4464 44714 4520 44716
rect 4464 44662 4466 44714
rect 4466 44662 4518 44714
rect 4518 44662 4520 44714
rect 4464 44660 4520 44662
rect 4568 44714 4624 44716
rect 4568 44662 4570 44714
rect 4570 44662 4622 44714
rect 4622 44662 4624 44714
rect 4568 44660 4624 44662
rect 4672 44714 4728 44716
rect 4672 44662 4674 44714
rect 4674 44662 4726 44714
rect 4726 44662 4728 44714
rect 4672 44660 4728 44662
rect 3804 43930 3860 43932
rect 3804 43878 3806 43930
rect 3806 43878 3858 43930
rect 3858 43878 3860 43930
rect 3804 43876 3860 43878
rect 3908 43930 3964 43932
rect 3908 43878 3910 43930
rect 3910 43878 3962 43930
rect 3962 43878 3964 43930
rect 3908 43876 3964 43878
rect 4012 43930 4068 43932
rect 4012 43878 4014 43930
rect 4014 43878 4066 43930
rect 4066 43878 4068 43930
rect 4012 43876 4068 43878
rect 4464 43146 4520 43148
rect 4464 43094 4466 43146
rect 4466 43094 4518 43146
rect 4518 43094 4520 43146
rect 4464 43092 4520 43094
rect 4568 43146 4624 43148
rect 4568 43094 4570 43146
rect 4570 43094 4622 43146
rect 4622 43094 4624 43146
rect 4568 43092 4624 43094
rect 4672 43146 4728 43148
rect 4672 43094 4674 43146
rect 4674 43094 4726 43146
rect 4726 43094 4728 43146
rect 4672 43092 4728 43094
rect 3804 42362 3860 42364
rect 3804 42310 3806 42362
rect 3806 42310 3858 42362
rect 3858 42310 3860 42362
rect 3804 42308 3860 42310
rect 3908 42362 3964 42364
rect 3908 42310 3910 42362
rect 3910 42310 3962 42362
rect 3962 42310 3964 42362
rect 3908 42308 3964 42310
rect 4012 42362 4068 42364
rect 4012 42310 4014 42362
rect 4014 42310 4066 42362
rect 4066 42310 4068 42362
rect 4012 42308 4068 42310
rect 5516 42028 5572 42084
rect 4464 41578 4520 41580
rect 4464 41526 4466 41578
rect 4466 41526 4518 41578
rect 4518 41526 4520 41578
rect 4464 41524 4520 41526
rect 4568 41578 4624 41580
rect 4568 41526 4570 41578
rect 4570 41526 4622 41578
rect 4622 41526 4624 41578
rect 4568 41524 4624 41526
rect 4672 41578 4728 41580
rect 4672 41526 4674 41578
rect 4674 41526 4726 41578
rect 4726 41526 4728 41578
rect 4672 41524 4728 41526
rect 3804 40794 3860 40796
rect 3804 40742 3806 40794
rect 3806 40742 3858 40794
rect 3858 40742 3860 40794
rect 3804 40740 3860 40742
rect 3908 40794 3964 40796
rect 3908 40742 3910 40794
rect 3910 40742 3962 40794
rect 3962 40742 3964 40794
rect 3908 40740 3964 40742
rect 4012 40794 4068 40796
rect 4012 40742 4014 40794
rect 4014 40742 4066 40794
rect 4066 40742 4068 40794
rect 4012 40740 4068 40742
rect 4464 40010 4520 40012
rect 4464 39958 4466 40010
rect 4466 39958 4518 40010
rect 4518 39958 4520 40010
rect 4464 39956 4520 39958
rect 4568 40010 4624 40012
rect 4568 39958 4570 40010
rect 4570 39958 4622 40010
rect 4622 39958 4624 40010
rect 4568 39956 4624 39958
rect 4672 40010 4728 40012
rect 4672 39958 4674 40010
rect 4674 39958 4726 40010
rect 4726 39958 4728 40010
rect 4672 39956 4728 39958
rect 3500 39676 3556 39732
rect 3948 39618 4004 39620
rect 3948 39566 3950 39618
rect 3950 39566 4002 39618
rect 4002 39566 4004 39618
rect 3948 39564 4004 39566
rect 3500 39340 3556 39396
rect 5180 39340 5236 39396
rect 3804 39226 3860 39228
rect 3804 39174 3806 39226
rect 3806 39174 3858 39226
rect 3858 39174 3860 39226
rect 3804 39172 3860 39174
rect 3908 39226 3964 39228
rect 3908 39174 3910 39226
rect 3910 39174 3962 39226
rect 3962 39174 3964 39226
rect 3908 39172 3964 39174
rect 4012 39226 4068 39228
rect 4012 39174 4014 39226
rect 4014 39174 4066 39226
rect 4066 39174 4068 39226
rect 4012 39172 4068 39174
rect 4172 38444 4228 38500
rect 3388 34130 3444 34132
rect 3388 34078 3390 34130
rect 3390 34078 3442 34130
rect 3442 34078 3444 34130
rect 3388 34076 3444 34078
rect 2940 33628 2996 33684
rect 2604 33404 2660 33460
rect 2380 28754 2436 28756
rect 2380 28702 2382 28754
rect 2382 28702 2434 28754
rect 2434 28702 2436 28754
rect 2380 28700 2436 28702
rect 2492 31836 2548 31892
rect 1932 26236 1988 26292
rect 1708 22988 1764 23044
rect 1932 23772 1988 23828
rect 1596 22482 1652 22484
rect 1596 22430 1598 22482
rect 1598 22430 1650 22482
rect 1650 22430 1652 22482
rect 1596 22428 1652 22430
rect 1484 22204 1540 22260
rect 1708 22204 1764 22260
rect 1596 22092 1652 22148
rect 1484 21980 1540 22036
rect 1148 19292 1204 19348
rect 1036 17500 1092 17556
rect 1260 17052 1316 17108
rect 1148 12124 1204 12180
rect 1372 16268 1428 16324
rect 1372 15260 1428 15316
rect 1372 13916 1428 13972
rect 1260 9266 1316 9268
rect 1260 9214 1262 9266
rect 1262 9214 1314 9266
rect 1314 9214 1316 9266
rect 1260 9212 1316 9214
rect 1596 18956 1652 19012
rect 1820 20914 1876 20916
rect 1820 20862 1822 20914
rect 1822 20862 1874 20914
rect 1874 20862 1876 20914
rect 1820 20860 1876 20862
rect 1596 18732 1652 18788
rect 1820 17388 1876 17444
rect 1708 17052 1764 17108
rect 1820 16828 1876 16884
rect 1596 16770 1652 16772
rect 1596 16718 1598 16770
rect 1598 16718 1650 16770
rect 1650 16718 1652 16770
rect 1596 16716 1652 16718
rect 1820 16210 1876 16212
rect 1820 16158 1822 16210
rect 1822 16158 1874 16210
rect 1874 16158 1876 16210
rect 1820 16156 1876 16158
rect 1820 15260 1876 15316
rect 1596 15148 1652 15204
rect 2716 31836 2772 31892
rect 2716 30268 2772 30324
rect 2604 30210 2660 30212
rect 2604 30158 2606 30210
rect 2606 30158 2658 30210
rect 2658 30158 2660 30210
rect 2604 30156 2660 30158
rect 2604 29426 2660 29428
rect 2604 29374 2606 29426
rect 2606 29374 2658 29426
rect 2658 29374 2660 29426
rect 2604 29372 2660 29374
rect 2604 28924 2660 28980
rect 2268 25788 2324 25844
rect 2380 24610 2436 24612
rect 2380 24558 2382 24610
rect 2382 24558 2434 24610
rect 2434 24558 2436 24610
rect 2380 24556 2436 24558
rect 2380 24332 2436 24388
rect 2380 23938 2436 23940
rect 2380 23886 2382 23938
rect 2382 23886 2434 23938
rect 2434 23886 2436 23938
rect 2380 23884 2436 23886
rect 2268 23266 2324 23268
rect 2268 23214 2270 23266
rect 2270 23214 2322 23266
rect 2322 23214 2324 23266
rect 2268 23212 2324 23214
rect 2044 22764 2100 22820
rect 2156 21644 2212 21700
rect 2268 22988 2324 23044
rect 2156 20690 2212 20692
rect 2156 20638 2158 20690
rect 2158 20638 2210 20690
rect 2210 20638 2212 20690
rect 2156 20636 2212 20638
rect 2268 19516 2324 19572
rect 2604 24780 2660 24836
rect 3804 37658 3860 37660
rect 3804 37606 3806 37658
rect 3806 37606 3858 37658
rect 3858 37606 3860 37658
rect 3804 37604 3860 37606
rect 3908 37658 3964 37660
rect 3908 37606 3910 37658
rect 3910 37606 3962 37658
rect 3962 37606 3964 37658
rect 3908 37604 3964 37606
rect 4012 37658 4068 37660
rect 4012 37606 4014 37658
rect 4014 37606 4066 37658
rect 4066 37606 4068 37658
rect 4012 37604 4068 37606
rect 4464 38442 4520 38444
rect 4464 38390 4466 38442
rect 4466 38390 4518 38442
rect 4518 38390 4520 38442
rect 4464 38388 4520 38390
rect 4568 38442 4624 38444
rect 4568 38390 4570 38442
rect 4570 38390 4622 38442
rect 4622 38390 4624 38442
rect 4568 38388 4624 38390
rect 4672 38442 4728 38444
rect 4672 38390 4674 38442
rect 4674 38390 4726 38442
rect 4726 38390 4728 38442
rect 4672 38388 4728 38390
rect 4732 37884 4788 37940
rect 4396 37772 4452 37828
rect 5068 37772 5124 37828
rect 4172 37100 4228 37156
rect 4844 37324 4900 37380
rect 3804 36090 3860 36092
rect 3804 36038 3806 36090
rect 3806 36038 3858 36090
rect 3858 36038 3860 36090
rect 3804 36036 3860 36038
rect 3908 36090 3964 36092
rect 3908 36038 3910 36090
rect 3910 36038 3962 36090
rect 3962 36038 3964 36090
rect 3908 36036 3964 36038
rect 4012 36090 4068 36092
rect 4012 36038 4014 36090
rect 4014 36038 4066 36090
rect 4066 36038 4068 36090
rect 4012 36036 4068 36038
rect 3724 35308 3780 35364
rect 3612 35084 3668 35140
rect 3948 34972 4004 35028
rect 4464 36874 4520 36876
rect 4464 36822 4466 36874
rect 4466 36822 4518 36874
rect 4518 36822 4520 36874
rect 4464 36820 4520 36822
rect 4568 36874 4624 36876
rect 4568 36822 4570 36874
rect 4570 36822 4622 36874
rect 4622 36822 4624 36874
rect 4568 36820 4624 36822
rect 4672 36874 4728 36876
rect 4672 36822 4674 36874
rect 4674 36822 4726 36874
rect 4726 36822 4728 36874
rect 4672 36820 4728 36822
rect 4396 35698 4452 35700
rect 4396 35646 4398 35698
rect 4398 35646 4450 35698
rect 4450 35646 4452 35698
rect 4396 35644 4452 35646
rect 4844 35532 4900 35588
rect 4464 35306 4520 35308
rect 4464 35254 4466 35306
rect 4466 35254 4518 35306
rect 4518 35254 4520 35306
rect 4464 35252 4520 35254
rect 4568 35306 4624 35308
rect 4568 35254 4570 35306
rect 4570 35254 4622 35306
rect 4622 35254 4624 35306
rect 4568 35252 4624 35254
rect 4672 35306 4728 35308
rect 4672 35254 4674 35306
rect 4674 35254 4726 35306
rect 4726 35254 4728 35306
rect 4672 35252 4728 35254
rect 3804 34522 3860 34524
rect 3804 34470 3806 34522
rect 3806 34470 3858 34522
rect 3858 34470 3860 34522
rect 3804 34468 3860 34470
rect 3908 34522 3964 34524
rect 3908 34470 3910 34522
rect 3910 34470 3962 34522
rect 3962 34470 3964 34522
rect 3908 34468 3964 34470
rect 4012 34522 4068 34524
rect 4012 34470 4014 34522
rect 4014 34470 4066 34522
rect 4066 34470 4068 34522
rect 4012 34468 4068 34470
rect 4284 34412 4340 34468
rect 3612 33852 3668 33908
rect 4172 34300 4228 34356
rect 3276 31778 3332 31780
rect 3276 31726 3278 31778
rect 3278 31726 3330 31778
rect 3330 31726 3332 31778
rect 3276 31724 3332 31726
rect 3164 30770 3220 30772
rect 3164 30718 3166 30770
rect 3166 30718 3218 30770
rect 3218 30718 3220 30770
rect 3164 30716 3220 30718
rect 3164 30044 3220 30100
rect 2828 27132 2884 27188
rect 3052 29820 3108 29876
rect 3804 32954 3860 32956
rect 3804 32902 3806 32954
rect 3806 32902 3858 32954
rect 3858 32902 3860 32954
rect 3804 32900 3860 32902
rect 3908 32954 3964 32956
rect 3908 32902 3910 32954
rect 3910 32902 3962 32954
rect 3962 32902 3964 32954
rect 3908 32900 3964 32902
rect 4012 32954 4068 32956
rect 4012 32902 4014 32954
rect 4014 32902 4066 32954
rect 4066 32902 4068 32954
rect 4012 32900 4068 32902
rect 4844 34076 4900 34132
rect 3612 31724 3668 31780
rect 4464 33738 4520 33740
rect 4464 33686 4466 33738
rect 4466 33686 4518 33738
rect 4518 33686 4520 33738
rect 4464 33684 4520 33686
rect 4568 33738 4624 33740
rect 4568 33686 4570 33738
rect 4570 33686 4622 33738
rect 4622 33686 4624 33738
rect 4568 33684 4624 33686
rect 4672 33738 4728 33740
rect 4672 33686 4674 33738
rect 4674 33686 4726 33738
rect 4726 33686 4728 33738
rect 4672 33684 4728 33686
rect 4464 32170 4520 32172
rect 4464 32118 4466 32170
rect 4466 32118 4518 32170
rect 4518 32118 4520 32170
rect 4464 32116 4520 32118
rect 4568 32170 4624 32172
rect 4568 32118 4570 32170
rect 4570 32118 4622 32170
rect 4622 32118 4624 32170
rect 4568 32116 4624 32118
rect 4672 32170 4728 32172
rect 4672 32118 4674 32170
rect 4674 32118 4726 32170
rect 4726 32118 4728 32170
rect 4672 32116 4728 32118
rect 3804 31386 3860 31388
rect 3804 31334 3806 31386
rect 3806 31334 3858 31386
rect 3858 31334 3860 31386
rect 3804 31332 3860 31334
rect 3908 31386 3964 31388
rect 3908 31334 3910 31386
rect 3910 31334 3962 31386
rect 3962 31334 3964 31386
rect 3908 31332 3964 31334
rect 4012 31386 4068 31388
rect 4012 31334 4014 31386
rect 4014 31334 4066 31386
rect 4066 31334 4068 31386
rect 4012 31332 4068 31334
rect 4284 31218 4340 31220
rect 4284 31166 4286 31218
rect 4286 31166 4338 31218
rect 4338 31166 4340 31218
rect 4284 31164 4340 31166
rect 4464 30602 4520 30604
rect 4464 30550 4466 30602
rect 4466 30550 4518 30602
rect 4518 30550 4520 30602
rect 4464 30548 4520 30550
rect 4568 30602 4624 30604
rect 4568 30550 4570 30602
rect 4570 30550 4622 30602
rect 4622 30550 4624 30602
rect 4568 30548 4624 30550
rect 4672 30602 4728 30604
rect 4672 30550 4674 30602
rect 4674 30550 4726 30602
rect 4726 30550 4728 30602
rect 4672 30548 4728 30550
rect 4172 30268 4228 30324
rect 3388 29932 3444 29988
rect 3500 28812 3556 28868
rect 3804 29818 3860 29820
rect 3804 29766 3806 29818
rect 3806 29766 3858 29818
rect 3858 29766 3860 29818
rect 3804 29764 3860 29766
rect 3908 29818 3964 29820
rect 3908 29766 3910 29818
rect 3910 29766 3962 29818
rect 3962 29766 3964 29818
rect 3908 29764 3964 29766
rect 4012 29818 4068 29820
rect 4012 29766 4014 29818
rect 4014 29766 4066 29818
rect 4066 29766 4068 29818
rect 4012 29764 4068 29766
rect 4396 30380 4452 30436
rect 4284 30044 4340 30100
rect 4284 29650 4340 29652
rect 4284 29598 4286 29650
rect 4286 29598 4338 29650
rect 4338 29598 4340 29650
rect 4284 29596 4340 29598
rect 3164 27244 3220 27300
rect 4508 30156 4564 30212
rect 4172 29372 4228 29428
rect 3276 27132 3332 27188
rect 3276 26962 3332 26964
rect 3276 26910 3278 26962
rect 3278 26910 3330 26962
rect 3330 26910 3332 26962
rect 3276 26908 3332 26910
rect 3052 26460 3108 26516
rect 3052 25788 3108 25844
rect 2716 23100 2772 23156
rect 2604 22764 2660 22820
rect 2940 22988 2996 23044
rect 2716 21698 2772 21700
rect 2716 21646 2718 21698
rect 2718 21646 2770 21698
rect 2770 21646 2772 21698
rect 2716 21644 2772 21646
rect 2380 18844 2436 18900
rect 2156 18620 2212 18676
rect 2268 18508 2324 18564
rect 2044 16716 2100 16772
rect 2380 16156 2436 16212
rect 2268 15148 2324 15204
rect 2156 15036 2212 15092
rect 1708 13692 1764 13748
rect 1820 13244 1876 13300
rect 1596 11618 1652 11620
rect 1596 11566 1598 11618
rect 1598 11566 1650 11618
rect 1650 11566 1652 11618
rect 1596 11564 1652 11566
rect 2044 12178 2100 12180
rect 2044 12126 2046 12178
rect 2046 12126 2098 12178
rect 2098 12126 2100 12178
rect 2044 12124 2100 12126
rect 1932 11564 1988 11620
rect 1932 10668 1988 10724
rect 2044 10444 2100 10500
rect 1596 8204 1652 8260
rect 1484 6748 1540 6804
rect 1596 5516 1652 5572
rect 1036 4956 1092 5012
rect 1484 4060 1540 4116
rect 1260 3164 1316 3220
rect 1484 2882 1540 2884
rect 1484 2830 1486 2882
rect 1486 2830 1538 2882
rect 1538 2830 1540 2882
rect 1484 2828 1540 2830
rect 1036 2268 1092 2324
rect 2268 13522 2324 13524
rect 2268 13470 2270 13522
rect 2270 13470 2322 13522
rect 2322 13470 2324 13522
rect 2268 13468 2324 13470
rect 2268 13244 2324 13300
rect 2268 12124 2324 12180
rect 2380 12908 2436 12964
rect 3164 23772 3220 23828
rect 3388 25340 3444 25396
rect 3804 28250 3860 28252
rect 3804 28198 3806 28250
rect 3806 28198 3858 28250
rect 3858 28198 3860 28250
rect 3804 28196 3860 28198
rect 3908 28250 3964 28252
rect 3908 28198 3910 28250
rect 3910 28198 3962 28250
rect 3962 28198 3964 28250
rect 3908 28196 3964 28198
rect 4012 28250 4068 28252
rect 4012 28198 4014 28250
rect 4014 28198 4066 28250
rect 4066 28198 4068 28250
rect 4012 28196 4068 28198
rect 4464 29034 4520 29036
rect 4464 28982 4466 29034
rect 4466 28982 4518 29034
rect 4518 28982 4520 29034
rect 4464 28980 4520 28982
rect 4568 29034 4624 29036
rect 4568 28982 4570 29034
rect 4570 28982 4622 29034
rect 4622 28982 4624 29034
rect 4568 28980 4624 28982
rect 4672 29034 4728 29036
rect 4672 28982 4674 29034
rect 4674 28982 4726 29034
rect 4726 28982 4728 29034
rect 4672 28980 4728 28982
rect 4060 27132 4116 27188
rect 4464 27466 4520 27468
rect 4464 27414 4466 27466
rect 4466 27414 4518 27466
rect 4518 27414 4520 27466
rect 4464 27412 4520 27414
rect 4568 27466 4624 27468
rect 4568 27414 4570 27466
rect 4570 27414 4622 27466
rect 4622 27414 4624 27466
rect 4568 27412 4624 27414
rect 4672 27466 4728 27468
rect 4672 27414 4674 27466
rect 4674 27414 4726 27466
rect 4726 27414 4728 27466
rect 4672 27412 4728 27414
rect 4284 27298 4340 27300
rect 4284 27246 4286 27298
rect 4286 27246 4338 27298
rect 4338 27246 4340 27298
rect 4284 27244 4340 27246
rect 3804 26682 3860 26684
rect 3804 26630 3806 26682
rect 3806 26630 3858 26682
rect 3858 26630 3860 26682
rect 3804 26628 3860 26630
rect 3908 26682 3964 26684
rect 3908 26630 3910 26682
rect 3910 26630 3962 26682
rect 3962 26630 3964 26682
rect 3908 26628 3964 26630
rect 4012 26682 4068 26684
rect 4012 26630 4014 26682
rect 4014 26630 4066 26682
rect 4066 26630 4068 26682
rect 4012 26628 4068 26630
rect 3612 25730 3668 25732
rect 3612 25678 3614 25730
rect 3614 25678 3666 25730
rect 3666 25678 3668 25730
rect 3612 25676 3668 25678
rect 3804 25114 3860 25116
rect 3804 25062 3806 25114
rect 3806 25062 3858 25114
rect 3858 25062 3860 25114
rect 3804 25060 3860 25062
rect 3908 25114 3964 25116
rect 3908 25062 3910 25114
rect 3910 25062 3962 25114
rect 3962 25062 3964 25114
rect 3908 25060 3964 25062
rect 4012 25114 4068 25116
rect 4012 25062 4014 25114
rect 4014 25062 4066 25114
rect 4066 25062 4068 25114
rect 4012 25060 4068 25062
rect 4172 25116 4228 25172
rect 3724 24668 3780 24724
rect 3388 23548 3444 23604
rect 3500 23996 3556 24052
rect 3276 23100 3332 23156
rect 3052 22428 3108 22484
rect 2828 18508 2884 18564
rect 2716 17724 2772 17780
rect 3052 20972 3108 21028
rect 4172 24332 4228 24388
rect 3724 23996 3780 24052
rect 3804 23546 3860 23548
rect 3804 23494 3806 23546
rect 3806 23494 3858 23546
rect 3858 23494 3860 23546
rect 3804 23492 3860 23494
rect 3908 23546 3964 23548
rect 3908 23494 3910 23546
rect 3910 23494 3962 23546
rect 3962 23494 3964 23546
rect 3908 23492 3964 23494
rect 4012 23546 4068 23548
rect 4012 23494 4014 23546
rect 4014 23494 4066 23546
rect 4066 23494 4068 23546
rect 4012 23492 4068 23494
rect 4464 25898 4520 25900
rect 4464 25846 4466 25898
rect 4466 25846 4518 25898
rect 4518 25846 4520 25898
rect 4464 25844 4520 25846
rect 4568 25898 4624 25900
rect 4568 25846 4570 25898
rect 4570 25846 4622 25898
rect 4622 25846 4624 25898
rect 4568 25844 4624 25846
rect 4672 25898 4728 25900
rect 4672 25846 4674 25898
rect 4674 25846 4726 25898
rect 4726 25846 4728 25898
rect 4672 25844 4728 25846
rect 4956 32732 5012 32788
rect 5068 33852 5124 33908
rect 5404 39228 5460 39284
rect 5404 37772 5460 37828
rect 5292 35420 5348 35476
rect 5404 36092 5460 36148
rect 4956 31836 5012 31892
rect 5068 31666 5124 31668
rect 5068 31614 5070 31666
rect 5070 31614 5122 31666
rect 5122 31614 5124 31666
rect 5068 31612 5124 31614
rect 4956 30604 5012 30660
rect 5068 30156 5124 30212
rect 4956 29596 5012 29652
rect 5068 29932 5124 29988
rect 4956 29372 5012 29428
rect 4956 27804 5012 27860
rect 4956 27244 5012 27300
rect 4956 25676 5012 25732
rect 4620 24556 4676 24612
rect 4464 24330 4520 24332
rect 4464 24278 4466 24330
rect 4466 24278 4518 24330
rect 4518 24278 4520 24330
rect 4464 24276 4520 24278
rect 4568 24330 4624 24332
rect 4568 24278 4570 24330
rect 4570 24278 4622 24330
rect 4622 24278 4624 24330
rect 4568 24276 4624 24278
rect 4672 24330 4728 24332
rect 4672 24278 4674 24330
rect 4674 24278 4726 24330
rect 4726 24278 4728 24330
rect 4672 24276 4728 24278
rect 4620 23548 4676 23604
rect 4464 22762 4520 22764
rect 4464 22710 4466 22762
rect 4466 22710 4518 22762
rect 4518 22710 4520 22762
rect 4464 22708 4520 22710
rect 4568 22762 4624 22764
rect 4568 22710 4570 22762
rect 4570 22710 4622 22762
rect 4622 22710 4624 22762
rect 4568 22708 4624 22710
rect 4672 22762 4728 22764
rect 4672 22710 4674 22762
rect 4674 22710 4726 22762
rect 4726 22710 4728 22762
rect 4672 22708 4728 22710
rect 3804 21978 3860 21980
rect 3804 21926 3806 21978
rect 3806 21926 3858 21978
rect 3858 21926 3860 21978
rect 3804 21924 3860 21926
rect 3908 21978 3964 21980
rect 3908 21926 3910 21978
rect 3910 21926 3962 21978
rect 3962 21926 3964 21978
rect 3908 21924 3964 21926
rect 4012 21978 4068 21980
rect 4012 21926 4014 21978
rect 4014 21926 4066 21978
rect 4066 21926 4068 21978
rect 4012 21924 4068 21926
rect 5292 34860 5348 34916
rect 5292 34412 5348 34468
rect 5628 34076 5684 34132
rect 5516 33906 5572 33908
rect 5516 33854 5518 33906
rect 5518 33854 5570 33906
rect 5570 33854 5572 33906
rect 5516 33852 5572 33854
rect 5516 32338 5572 32340
rect 5516 32286 5518 32338
rect 5518 32286 5570 32338
rect 5570 32286 5572 32338
rect 5516 32284 5572 32286
rect 5404 31164 5460 31220
rect 5628 31612 5684 31668
rect 5292 30604 5348 30660
rect 5292 29372 5348 29428
rect 5180 28924 5236 28980
rect 5180 28700 5236 28756
rect 5292 27074 5348 27076
rect 5292 27022 5294 27074
rect 5294 27022 5346 27074
rect 5346 27022 5348 27074
rect 5292 27020 5348 27022
rect 5516 30828 5572 30884
rect 6860 55186 6916 55188
rect 6860 55134 6862 55186
rect 6862 55134 6914 55186
rect 6914 55134 6916 55186
rect 6860 55132 6916 55134
rect 7756 51212 7812 51268
rect 5852 41356 5908 41412
rect 7644 45724 7700 45780
rect 6748 42924 6804 42980
rect 5964 40236 6020 40292
rect 6076 40124 6132 40180
rect 5852 39788 5908 39844
rect 6300 40124 6356 40180
rect 6300 38668 6356 38724
rect 5852 34914 5908 34916
rect 5852 34862 5854 34914
rect 5854 34862 5906 34914
rect 5906 34862 5908 34914
rect 5852 34860 5908 34862
rect 6412 39452 6468 39508
rect 6636 39340 6692 39396
rect 6524 37884 6580 37940
rect 6524 37378 6580 37380
rect 6524 37326 6526 37378
rect 6526 37326 6578 37378
rect 6578 37326 6580 37378
rect 6524 37324 6580 37326
rect 6412 36428 6468 36484
rect 6524 35810 6580 35812
rect 6524 35758 6526 35810
rect 6526 35758 6578 35810
rect 6578 35758 6580 35810
rect 6524 35756 6580 35758
rect 6300 34076 6356 34132
rect 6188 33852 6244 33908
rect 5964 31836 6020 31892
rect 5740 30828 5796 30884
rect 5628 29426 5684 29428
rect 5628 29374 5630 29426
rect 5630 29374 5682 29426
rect 5682 29374 5684 29426
rect 5628 29372 5684 29374
rect 5628 28364 5684 28420
rect 5852 28700 5908 28756
rect 6076 28924 6132 28980
rect 5740 28140 5796 28196
rect 5964 28252 6020 28308
rect 5516 27356 5572 27412
rect 5740 27692 5796 27748
rect 5516 26684 5572 26740
rect 5516 25564 5572 25620
rect 5404 25004 5460 25060
rect 5292 24668 5348 24724
rect 5740 25676 5796 25732
rect 5740 25506 5796 25508
rect 5740 25454 5742 25506
rect 5742 25454 5794 25506
rect 5794 25454 5796 25506
rect 5740 25452 5796 25454
rect 5852 25116 5908 25172
rect 5964 27132 6020 27188
rect 5516 23938 5572 23940
rect 5516 23886 5518 23938
rect 5518 23886 5570 23938
rect 5570 23886 5572 23938
rect 5516 23884 5572 23886
rect 5852 23996 5908 24052
rect 4956 21756 5012 21812
rect 4956 21532 5012 21588
rect 3164 20914 3220 20916
rect 3164 20862 3166 20914
rect 3166 20862 3218 20914
rect 3218 20862 3220 20914
rect 3164 20860 3220 20862
rect 3804 20410 3860 20412
rect 3804 20358 3806 20410
rect 3806 20358 3858 20410
rect 3858 20358 3860 20410
rect 3804 20356 3860 20358
rect 3908 20410 3964 20412
rect 3908 20358 3910 20410
rect 3910 20358 3962 20410
rect 3962 20358 3964 20410
rect 3908 20356 3964 20358
rect 4012 20410 4068 20412
rect 4012 20358 4014 20410
rect 4014 20358 4066 20410
rect 4066 20358 4068 20410
rect 4012 20356 4068 20358
rect 3388 19516 3444 19572
rect 3388 18732 3444 18788
rect 3804 18842 3860 18844
rect 3804 18790 3806 18842
rect 3806 18790 3858 18842
rect 3858 18790 3860 18842
rect 3804 18788 3860 18790
rect 3908 18842 3964 18844
rect 3908 18790 3910 18842
rect 3910 18790 3962 18842
rect 3962 18790 3964 18842
rect 3908 18788 3964 18790
rect 4012 18842 4068 18844
rect 4012 18790 4014 18842
rect 4014 18790 4066 18842
rect 4066 18790 4068 18842
rect 4012 18788 4068 18790
rect 3052 18508 3108 18564
rect 3836 18508 3892 18564
rect 2940 17612 2996 17668
rect 2828 16156 2884 16212
rect 2828 15708 2884 15764
rect 2604 15314 2660 15316
rect 2604 15262 2606 15314
rect 2606 15262 2658 15314
rect 2658 15262 2660 15314
rect 2604 15260 2660 15262
rect 2716 15036 2772 15092
rect 2492 12236 2548 12292
rect 2604 12684 2660 12740
rect 2380 11564 2436 11620
rect 2492 9996 2548 10052
rect 2156 8652 2212 8708
rect 2716 11452 2772 11508
rect 2716 9996 2772 10052
rect 3164 16828 3220 16884
rect 3052 15148 3108 15204
rect 3948 17500 4004 17556
rect 3804 17274 3860 17276
rect 3804 17222 3806 17274
rect 3806 17222 3858 17274
rect 3858 17222 3860 17274
rect 3804 17220 3860 17222
rect 3908 17274 3964 17276
rect 3908 17222 3910 17274
rect 3910 17222 3962 17274
rect 3962 17222 3964 17274
rect 3908 17220 3964 17222
rect 4012 17274 4068 17276
rect 4012 17222 4014 17274
rect 4014 17222 4066 17274
rect 4066 17222 4068 17274
rect 4012 17220 4068 17222
rect 3836 16994 3892 16996
rect 3836 16942 3838 16994
rect 3838 16942 3890 16994
rect 3890 16942 3892 16994
rect 3836 16940 3892 16942
rect 4464 21194 4520 21196
rect 4464 21142 4466 21194
rect 4466 21142 4518 21194
rect 4518 21142 4520 21194
rect 4464 21140 4520 21142
rect 4568 21194 4624 21196
rect 4568 21142 4570 21194
rect 4570 21142 4622 21194
rect 4622 21142 4624 21194
rect 4568 21140 4624 21142
rect 4672 21194 4728 21196
rect 4672 21142 4674 21194
rect 4674 21142 4726 21194
rect 4726 21142 4728 21194
rect 4672 21140 4728 21142
rect 4956 20860 5012 20916
rect 4396 20636 4452 20692
rect 4284 19964 4340 20020
rect 4844 20188 4900 20244
rect 4464 19626 4520 19628
rect 4464 19574 4466 19626
rect 4466 19574 4518 19626
rect 4518 19574 4520 19626
rect 4464 19572 4520 19574
rect 4568 19626 4624 19628
rect 4568 19574 4570 19626
rect 4570 19574 4622 19626
rect 4622 19574 4624 19626
rect 4568 19572 4624 19574
rect 4672 19626 4728 19628
rect 4672 19574 4674 19626
rect 4674 19574 4726 19626
rect 4726 19574 4728 19626
rect 4672 19572 4728 19574
rect 4620 19234 4676 19236
rect 4620 19182 4622 19234
rect 4622 19182 4674 19234
rect 4674 19182 4676 19234
rect 4620 19180 4676 19182
rect 4464 18058 4520 18060
rect 4464 18006 4466 18058
rect 4466 18006 4518 18058
rect 4518 18006 4520 18058
rect 4464 18004 4520 18006
rect 4568 18058 4624 18060
rect 4568 18006 4570 18058
rect 4570 18006 4622 18058
rect 4622 18006 4624 18058
rect 4568 18004 4624 18006
rect 4672 18058 4728 18060
rect 4672 18006 4674 18058
rect 4674 18006 4726 18058
rect 4726 18006 4728 18058
rect 4672 18004 4728 18006
rect 4284 17836 4340 17892
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 4732 17164 4788 17220
rect 4464 16490 4520 16492
rect 4464 16438 4466 16490
rect 4466 16438 4518 16490
rect 4518 16438 4520 16490
rect 4464 16436 4520 16438
rect 4568 16490 4624 16492
rect 4568 16438 4570 16490
rect 4570 16438 4622 16490
rect 4622 16438 4624 16490
rect 4568 16436 4624 16438
rect 4672 16490 4728 16492
rect 4672 16438 4674 16490
rect 4674 16438 4726 16490
rect 4726 16438 4728 16490
rect 4672 16436 4728 16438
rect 4172 16268 4228 16324
rect 3612 16098 3668 16100
rect 3612 16046 3614 16098
rect 3614 16046 3666 16098
rect 3666 16046 3668 16098
rect 3612 16044 3668 16046
rect 3804 15706 3860 15708
rect 3804 15654 3806 15706
rect 3806 15654 3858 15706
rect 3858 15654 3860 15706
rect 3804 15652 3860 15654
rect 3908 15706 3964 15708
rect 3908 15654 3910 15706
rect 3910 15654 3962 15706
rect 3962 15654 3964 15706
rect 3908 15652 3964 15654
rect 4012 15706 4068 15708
rect 4012 15654 4014 15706
rect 4014 15654 4066 15706
rect 4066 15654 4068 15706
rect 4012 15652 4068 15654
rect 4060 15484 4116 15540
rect 3500 15372 3556 15428
rect 3388 13634 3444 13636
rect 3388 13582 3390 13634
rect 3390 13582 3442 13634
rect 3442 13582 3444 13634
rect 3388 13580 3444 13582
rect 3164 13132 3220 13188
rect 2940 9996 2996 10052
rect 3052 13020 3108 13076
rect 2940 9436 2996 9492
rect 2268 7980 2324 8036
rect 2380 7644 2436 7700
rect 2492 7532 2548 7588
rect 3724 15202 3780 15204
rect 3724 15150 3726 15202
rect 3726 15150 3778 15202
rect 3778 15150 3780 15202
rect 3724 15148 3780 15150
rect 4464 14922 4520 14924
rect 4464 14870 4466 14922
rect 4466 14870 4518 14922
rect 4518 14870 4520 14922
rect 4464 14868 4520 14870
rect 4568 14922 4624 14924
rect 4568 14870 4570 14922
rect 4570 14870 4622 14922
rect 4622 14870 4624 14922
rect 4568 14868 4624 14870
rect 4672 14922 4728 14924
rect 4672 14870 4674 14922
rect 4674 14870 4726 14922
rect 4726 14870 4728 14922
rect 4672 14868 4728 14870
rect 4172 14700 4228 14756
rect 4284 14530 4340 14532
rect 4284 14478 4286 14530
rect 4286 14478 4338 14530
rect 4338 14478 4340 14530
rect 4284 14476 4340 14478
rect 3804 14138 3860 14140
rect 3804 14086 3806 14138
rect 3806 14086 3858 14138
rect 3858 14086 3860 14138
rect 3804 14084 3860 14086
rect 3908 14138 3964 14140
rect 3908 14086 3910 14138
rect 3910 14086 3962 14138
rect 3962 14086 3964 14138
rect 3908 14084 3964 14086
rect 4012 14138 4068 14140
rect 4012 14086 4014 14138
rect 4014 14086 4066 14138
rect 4066 14086 4068 14138
rect 4012 14084 4068 14086
rect 3724 13916 3780 13972
rect 3948 13804 4004 13860
rect 4732 14306 4788 14308
rect 4732 14254 4734 14306
rect 4734 14254 4786 14306
rect 4786 14254 4788 14306
rect 4732 14252 4788 14254
rect 4396 14140 4452 14196
rect 5628 23324 5684 23380
rect 5516 22876 5572 22932
rect 5292 21420 5348 21476
rect 5404 21084 5460 21140
rect 5740 22930 5796 22932
rect 5740 22878 5742 22930
rect 5742 22878 5794 22930
rect 5794 22878 5796 22930
rect 5740 22876 5796 22878
rect 5628 22258 5684 22260
rect 5628 22206 5630 22258
rect 5630 22206 5682 22258
rect 5682 22206 5684 22258
rect 5628 22204 5684 22206
rect 5628 21644 5684 21700
rect 5068 18844 5124 18900
rect 5068 18562 5124 18564
rect 5068 18510 5070 18562
rect 5070 18510 5122 18562
rect 5122 18510 5124 18562
rect 5068 18508 5124 18510
rect 5068 18284 5124 18340
rect 5068 17778 5124 17780
rect 5068 17726 5070 17778
rect 5070 17726 5122 17778
rect 5122 17726 5124 17778
rect 5068 17724 5124 17726
rect 5404 19234 5460 19236
rect 5404 19182 5406 19234
rect 5406 19182 5458 19234
rect 5458 19182 5460 19234
rect 5404 19180 5460 19182
rect 5852 20972 5908 21028
rect 5852 20578 5908 20580
rect 5852 20526 5854 20578
rect 5854 20526 5906 20578
rect 5906 20526 5908 20578
rect 5852 20524 5908 20526
rect 6412 33628 6468 33684
rect 6300 30380 6356 30436
rect 6524 30210 6580 30212
rect 6524 30158 6526 30210
rect 6526 30158 6578 30210
rect 6578 30158 6580 30210
rect 6524 30156 6580 30158
rect 6412 29596 6468 29652
rect 6188 25228 6244 25284
rect 6524 28364 6580 28420
rect 6412 26572 6468 26628
rect 6412 26402 6468 26404
rect 6412 26350 6414 26402
rect 6414 26350 6466 26402
rect 6466 26350 6468 26402
rect 6412 26348 6468 26350
rect 7308 39730 7364 39732
rect 7308 39678 7310 39730
rect 7310 39678 7362 39730
rect 7362 39678 7364 39730
rect 7308 39676 7364 39678
rect 6860 38780 6916 38836
rect 9100 52108 9156 52164
rect 8876 46508 8932 46564
rect 8092 42812 8148 42868
rect 8540 44940 8596 44996
rect 8316 42140 8372 42196
rect 8540 42028 8596 42084
rect 8652 42476 8708 42532
rect 7868 41020 7924 41076
rect 6860 38556 6916 38612
rect 7084 34412 7140 34468
rect 6972 33852 7028 33908
rect 6860 33404 6916 33460
rect 7196 33292 7252 33348
rect 7532 34524 7588 34580
rect 7868 39004 7924 39060
rect 7756 33906 7812 33908
rect 7756 33854 7758 33906
rect 7758 33854 7810 33906
rect 7810 33854 7812 33906
rect 7756 33852 7812 33854
rect 7420 31612 7476 31668
rect 7308 31388 7364 31444
rect 7308 30882 7364 30884
rect 7308 30830 7310 30882
rect 7310 30830 7362 30882
rect 7362 30830 7364 30882
rect 7308 30828 7364 30830
rect 6972 29708 7028 29764
rect 7196 29650 7252 29652
rect 7196 29598 7198 29650
rect 7198 29598 7250 29650
rect 7250 29598 7252 29650
rect 7196 29596 7252 29598
rect 7308 29484 7364 29540
rect 7308 28364 7364 28420
rect 7420 28252 7476 28308
rect 7420 28082 7476 28084
rect 7420 28030 7422 28082
rect 7422 28030 7474 28082
rect 7474 28030 7476 28082
rect 7420 28028 7476 28030
rect 6300 23996 6356 24052
rect 6748 26012 6804 26068
rect 6076 23100 6132 23156
rect 6300 23154 6356 23156
rect 6300 23102 6302 23154
rect 6302 23102 6354 23154
rect 6354 23102 6356 23154
rect 6300 23100 6356 23102
rect 6188 20748 6244 20804
rect 5740 18956 5796 19012
rect 6076 18732 6132 18788
rect 5404 18284 5460 18340
rect 5180 17276 5236 17332
rect 5516 17276 5572 17332
rect 4956 16492 5012 16548
rect 4844 13916 4900 13972
rect 4956 16268 5012 16324
rect 4956 13804 5012 13860
rect 4956 13634 5012 13636
rect 4956 13582 4958 13634
rect 4958 13582 5010 13634
rect 5010 13582 5012 13634
rect 4956 13580 5012 13582
rect 4844 13468 4900 13524
rect 4464 13354 4520 13356
rect 4464 13302 4466 13354
rect 4466 13302 4518 13354
rect 4518 13302 4520 13354
rect 4464 13300 4520 13302
rect 4568 13354 4624 13356
rect 4568 13302 4570 13354
rect 4570 13302 4622 13354
rect 4622 13302 4624 13354
rect 4568 13300 4624 13302
rect 4672 13354 4728 13356
rect 4672 13302 4674 13354
rect 4674 13302 4726 13354
rect 4726 13302 4728 13354
rect 4672 13300 4728 13302
rect 3164 12124 3220 12180
rect 3276 11228 3332 11284
rect 3164 8652 3220 8708
rect 3804 12570 3860 12572
rect 3804 12518 3806 12570
rect 3806 12518 3858 12570
rect 3858 12518 3860 12570
rect 3804 12516 3860 12518
rect 3908 12570 3964 12572
rect 3908 12518 3910 12570
rect 3910 12518 3962 12570
rect 3962 12518 3964 12570
rect 3908 12516 3964 12518
rect 4012 12570 4068 12572
rect 4012 12518 4014 12570
rect 4014 12518 4066 12570
rect 4066 12518 4068 12570
rect 4012 12516 4068 12518
rect 4172 12460 4228 12516
rect 3612 12402 3668 12404
rect 3612 12350 3614 12402
rect 3614 12350 3666 12402
rect 3666 12350 3668 12402
rect 3612 12348 3668 12350
rect 3612 11900 3668 11956
rect 4172 12012 4228 12068
rect 3804 11002 3860 11004
rect 3804 10950 3806 11002
rect 3806 10950 3858 11002
rect 3858 10950 3860 11002
rect 3804 10948 3860 10950
rect 3908 11002 3964 11004
rect 3908 10950 3910 11002
rect 3910 10950 3962 11002
rect 3962 10950 3964 11002
rect 3908 10948 3964 10950
rect 4012 11002 4068 11004
rect 4012 10950 4014 11002
rect 4014 10950 4066 11002
rect 4066 10950 4068 11002
rect 4012 10948 4068 10950
rect 3836 9826 3892 9828
rect 3836 9774 3838 9826
rect 3838 9774 3890 9826
rect 3890 9774 3892 9826
rect 3836 9772 3892 9774
rect 3804 9434 3860 9436
rect 3804 9382 3806 9434
rect 3806 9382 3858 9434
rect 3858 9382 3860 9434
rect 3804 9380 3860 9382
rect 3908 9434 3964 9436
rect 3908 9382 3910 9434
rect 3910 9382 3962 9434
rect 3962 9382 3964 9434
rect 3908 9380 3964 9382
rect 4012 9434 4068 9436
rect 4012 9382 4014 9434
rect 4014 9382 4066 9434
rect 4066 9382 4068 9434
rect 4012 9380 4068 9382
rect 4464 11786 4520 11788
rect 4464 11734 4466 11786
rect 4466 11734 4518 11786
rect 4518 11734 4520 11786
rect 4464 11732 4520 11734
rect 4568 11786 4624 11788
rect 4568 11734 4570 11786
rect 4570 11734 4622 11786
rect 4622 11734 4624 11786
rect 4568 11732 4624 11734
rect 4672 11786 4728 11788
rect 4672 11734 4674 11786
rect 4674 11734 4726 11786
rect 4726 11734 4728 11786
rect 4672 11732 4728 11734
rect 4284 11116 4340 11172
rect 5292 16604 5348 16660
rect 5180 15484 5236 15540
rect 5068 12348 5124 12404
rect 5404 15260 5460 15316
rect 5740 16828 5796 16884
rect 5628 15932 5684 15988
rect 5964 18284 6020 18340
rect 6076 17778 6132 17780
rect 6076 17726 6078 17778
rect 6078 17726 6130 17778
rect 6130 17726 6132 17778
rect 6076 17724 6132 17726
rect 5964 17500 6020 17556
rect 5852 16268 5908 16324
rect 5852 15260 5908 15316
rect 5516 13970 5572 13972
rect 5516 13918 5518 13970
rect 5518 13918 5570 13970
rect 5570 13918 5572 13970
rect 5516 13916 5572 13918
rect 5740 13244 5796 13300
rect 6300 15932 6356 15988
rect 6748 24108 6804 24164
rect 6860 25676 6916 25732
rect 6524 24050 6580 24052
rect 6524 23998 6526 24050
rect 6526 23998 6578 24050
rect 6578 23998 6580 24050
rect 6524 23996 6580 23998
rect 7420 26012 7476 26068
rect 7084 25228 7140 25284
rect 6972 24780 7028 24836
rect 6972 24332 7028 24388
rect 6524 21586 6580 21588
rect 6524 21534 6526 21586
rect 6526 21534 6578 21586
rect 6578 21534 6580 21586
rect 6524 21532 6580 21534
rect 6524 20524 6580 20580
rect 7196 23884 7252 23940
rect 6860 22764 6916 22820
rect 6860 21532 6916 21588
rect 7644 33458 7700 33460
rect 7644 33406 7646 33458
rect 7646 33406 7698 33458
rect 7698 33406 7700 33458
rect 7644 33404 7700 33406
rect 7644 32450 7700 32452
rect 7644 32398 7646 32450
rect 7646 32398 7698 32450
rect 7698 32398 7700 32450
rect 7644 32396 7700 32398
rect 8204 39004 8260 39060
rect 7980 38722 8036 38724
rect 7980 38670 7982 38722
rect 7982 38670 8034 38722
rect 8034 38670 8036 38722
rect 7980 38668 8036 38670
rect 8204 38274 8260 38276
rect 8204 38222 8206 38274
rect 8206 38222 8258 38274
rect 8258 38222 8260 38274
rect 8204 38220 8260 38222
rect 7980 35756 8036 35812
rect 8316 35868 8372 35924
rect 8204 34690 8260 34692
rect 8204 34638 8206 34690
rect 8206 34638 8258 34690
rect 8258 34638 8260 34690
rect 8204 34636 8260 34638
rect 8092 34076 8148 34132
rect 8204 34412 8260 34468
rect 7980 31612 8036 31668
rect 7756 29708 7812 29764
rect 7644 28140 7700 28196
rect 7084 23212 7140 23268
rect 6972 20914 7028 20916
rect 6972 20862 6974 20914
rect 6974 20862 7026 20914
rect 7026 20862 7028 20914
rect 6972 20860 7028 20862
rect 6860 20636 6916 20692
rect 6972 20188 7028 20244
rect 7196 20860 7252 20916
rect 7532 22876 7588 22932
rect 8204 31612 8260 31668
rect 8092 30268 8148 30324
rect 8092 29708 8148 29764
rect 7980 28252 8036 28308
rect 8092 28476 8148 28532
rect 8764 39116 8820 39172
rect 8764 38834 8820 38836
rect 8764 38782 8766 38834
rect 8766 38782 8818 38834
rect 8818 38782 8820 38834
rect 8764 38780 8820 38782
rect 8652 37266 8708 37268
rect 8652 37214 8654 37266
rect 8654 37214 8706 37266
rect 8706 37214 8708 37266
rect 8652 37212 8708 37214
rect 8764 36540 8820 36596
rect 8652 35420 8708 35476
rect 9100 45276 9156 45332
rect 9772 42700 9828 42756
rect 9548 39900 9604 39956
rect 9212 38668 9268 38724
rect 9884 42588 9940 42644
rect 10220 55244 10276 55300
rect 10108 41298 10164 41300
rect 10108 41246 10110 41298
rect 10110 41246 10162 41298
rect 10162 41246 10164 41298
rect 10108 41244 10164 41246
rect 9996 39676 10052 39732
rect 9884 38668 9940 38724
rect 9324 35420 9380 35476
rect 9212 35084 9268 35140
rect 9324 34972 9380 35028
rect 8876 34412 8932 34468
rect 9100 34636 9156 34692
rect 8652 33964 8708 34020
rect 8540 32732 8596 32788
rect 8652 33628 8708 33684
rect 8540 30044 8596 30100
rect 8540 29538 8596 29540
rect 8540 29486 8542 29538
rect 8542 29486 8594 29538
rect 8594 29486 8596 29538
rect 8540 29484 8596 29486
rect 8876 33628 8932 33684
rect 9324 33628 9380 33684
rect 8876 33458 8932 33460
rect 8876 33406 8878 33458
rect 8878 33406 8930 33458
rect 8930 33406 8932 33458
rect 8876 33404 8932 33406
rect 9548 38108 9604 38164
rect 8764 32844 8820 32900
rect 8652 27746 8708 27748
rect 8652 27694 8654 27746
rect 8654 27694 8706 27746
rect 8706 27694 8708 27746
rect 8652 27692 8708 27694
rect 8764 32620 8820 32676
rect 7756 26348 7812 26404
rect 7980 26066 8036 26068
rect 7980 26014 7982 26066
rect 7982 26014 8034 26066
rect 8034 26014 8036 26066
rect 7980 26012 8036 26014
rect 7756 25116 7812 25172
rect 8204 24668 8260 24724
rect 8428 24722 8484 24724
rect 8428 24670 8430 24722
rect 8430 24670 8482 24722
rect 8482 24670 8484 24722
rect 8428 24668 8484 24670
rect 8316 24444 8372 24500
rect 7756 23212 7812 23268
rect 7756 21868 7812 21924
rect 6524 18226 6580 18228
rect 6524 18174 6526 18226
rect 6526 18174 6578 18226
rect 6578 18174 6580 18226
rect 6524 18172 6580 18174
rect 6524 17836 6580 17892
rect 6636 15986 6692 15988
rect 6636 15934 6638 15986
rect 6638 15934 6690 15986
rect 6690 15934 6692 15986
rect 6636 15932 6692 15934
rect 6748 15708 6804 15764
rect 6972 16210 7028 16212
rect 6972 16158 6974 16210
rect 6974 16158 7026 16210
rect 7026 16158 7028 16210
rect 6972 16156 7028 16158
rect 7084 15708 7140 15764
rect 6188 14812 6244 14868
rect 6972 15148 7028 15204
rect 5404 11900 5460 11956
rect 5628 12236 5684 12292
rect 5404 11506 5460 11508
rect 5404 11454 5406 11506
rect 5406 11454 5458 11506
rect 5458 11454 5460 11506
rect 5404 11452 5460 11454
rect 4956 10780 5012 10836
rect 4464 10218 4520 10220
rect 4464 10166 4466 10218
rect 4466 10166 4518 10218
rect 4518 10166 4520 10218
rect 4464 10164 4520 10166
rect 4568 10218 4624 10220
rect 4568 10166 4570 10218
rect 4570 10166 4622 10218
rect 4622 10166 4624 10218
rect 4568 10164 4624 10166
rect 4672 10218 4728 10220
rect 4672 10166 4674 10218
rect 4674 10166 4726 10218
rect 4726 10166 4728 10218
rect 4672 10164 4728 10166
rect 5180 10780 5236 10836
rect 5852 11452 5908 11508
rect 5180 10332 5236 10388
rect 4464 8650 4520 8652
rect 4464 8598 4466 8650
rect 4466 8598 4518 8650
rect 4518 8598 4520 8650
rect 4464 8596 4520 8598
rect 4568 8650 4624 8652
rect 4568 8598 4570 8650
rect 4570 8598 4622 8650
rect 4622 8598 4624 8650
rect 4568 8596 4624 8598
rect 4672 8650 4728 8652
rect 4672 8598 4674 8650
rect 4674 8598 4726 8650
rect 4726 8598 4728 8650
rect 4672 8596 4728 8598
rect 5068 8034 5124 8036
rect 5068 7982 5070 8034
rect 5070 7982 5122 8034
rect 5122 7982 5124 8034
rect 5068 7980 5124 7982
rect 3804 7866 3860 7868
rect 3804 7814 3806 7866
rect 3806 7814 3858 7866
rect 3858 7814 3860 7866
rect 3804 7812 3860 7814
rect 3908 7866 3964 7868
rect 3908 7814 3910 7866
rect 3910 7814 3962 7866
rect 3962 7814 3964 7866
rect 3908 7812 3964 7814
rect 4012 7866 4068 7868
rect 4012 7814 4014 7866
rect 4014 7814 4066 7866
rect 4066 7814 4068 7866
rect 4012 7812 4068 7814
rect 3836 7474 3892 7476
rect 3836 7422 3838 7474
rect 3838 7422 3890 7474
rect 3890 7422 3892 7474
rect 3836 7420 3892 7422
rect 5292 9938 5348 9940
rect 5292 9886 5294 9938
rect 5294 9886 5346 9938
rect 5346 9886 5348 9938
rect 5292 9884 5348 9886
rect 5516 9154 5572 9156
rect 5516 9102 5518 9154
rect 5518 9102 5570 9154
rect 5570 9102 5572 9154
rect 5516 9100 5572 9102
rect 5516 8428 5572 8484
rect 4464 7082 4520 7084
rect 4464 7030 4466 7082
rect 4466 7030 4518 7082
rect 4518 7030 4520 7082
rect 4464 7028 4520 7030
rect 4568 7082 4624 7084
rect 4568 7030 4570 7082
rect 4570 7030 4622 7082
rect 4622 7030 4624 7082
rect 4568 7028 4624 7030
rect 4672 7082 4728 7084
rect 4672 7030 4674 7082
rect 4674 7030 4726 7082
rect 4726 7030 4728 7082
rect 4672 7028 4728 7030
rect 2828 5852 2884 5908
rect 3836 6524 3892 6580
rect 3500 6412 3556 6468
rect 3164 5794 3220 5796
rect 3164 5742 3166 5794
rect 3166 5742 3218 5794
rect 3218 5742 3220 5794
rect 3164 5740 3220 5742
rect 3804 6298 3860 6300
rect 3804 6246 3806 6298
rect 3806 6246 3858 6298
rect 3858 6246 3860 6298
rect 3804 6244 3860 6246
rect 3908 6298 3964 6300
rect 3908 6246 3910 6298
rect 3910 6246 3962 6298
rect 3962 6246 3964 6298
rect 3908 6244 3964 6246
rect 4012 6298 4068 6300
rect 4012 6246 4014 6298
rect 4014 6246 4066 6298
rect 4066 6246 4068 6298
rect 4012 6244 4068 6246
rect 6188 10220 6244 10276
rect 6188 8370 6244 8372
rect 6188 8318 6190 8370
rect 6190 8318 6242 8370
rect 6242 8318 6244 8370
rect 6188 8316 6244 8318
rect 6076 6076 6132 6132
rect 4464 5514 4520 5516
rect 4464 5462 4466 5514
rect 4466 5462 4518 5514
rect 4518 5462 4520 5514
rect 4464 5460 4520 5462
rect 4568 5514 4624 5516
rect 4568 5462 4570 5514
rect 4570 5462 4622 5514
rect 4622 5462 4624 5514
rect 4568 5460 4624 5462
rect 4672 5514 4728 5516
rect 4672 5462 4674 5514
rect 4674 5462 4726 5514
rect 4726 5462 4728 5514
rect 4672 5460 4728 5462
rect 4060 5122 4116 5124
rect 4060 5070 4062 5122
rect 4062 5070 4114 5122
rect 4114 5070 4116 5122
rect 4060 5068 4116 5070
rect 3804 4730 3860 4732
rect 3804 4678 3806 4730
rect 3806 4678 3858 4730
rect 3858 4678 3860 4730
rect 3804 4676 3860 4678
rect 3908 4730 3964 4732
rect 3908 4678 3910 4730
rect 3910 4678 3962 4730
rect 3962 4678 3964 4730
rect 3908 4676 3964 4678
rect 4012 4730 4068 4732
rect 4012 4678 4014 4730
rect 4014 4678 4066 4730
rect 4066 4678 4068 4730
rect 4012 4676 4068 4678
rect 2044 4284 2100 4340
rect 924 1596 980 1652
rect 700 588 756 644
rect 2268 4226 2324 4228
rect 2268 4174 2270 4226
rect 2270 4174 2322 4226
rect 2322 4174 2324 4226
rect 2268 4172 2324 4174
rect 4464 3946 4520 3948
rect 4464 3894 4466 3946
rect 4466 3894 4518 3946
rect 4518 3894 4520 3946
rect 4464 3892 4520 3894
rect 4568 3946 4624 3948
rect 4568 3894 4570 3946
rect 4570 3894 4622 3946
rect 4622 3894 4624 3946
rect 4568 3892 4624 3894
rect 4672 3946 4728 3948
rect 4672 3894 4674 3946
rect 4674 3894 4726 3946
rect 4726 3894 4728 3946
rect 4672 3892 4728 3894
rect 2268 3554 2324 3556
rect 2268 3502 2270 3554
rect 2270 3502 2322 3554
rect 2322 3502 2324 3554
rect 2268 3500 2324 3502
rect 6412 14588 6468 14644
rect 6412 12124 6468 12180
rect 6860 14642 6916 14644
rect 6860 14590 6862 14642
rect 6862 14590 6914 14642
rect 6914 14590 6916 14642
rect 6860 14588 6916 14590
rect 6972 12348 7028 12404
rect 7084 15036 7140 15092
rect 7308 20018 7364 20020
rect 7308 19966 7310 20018
rect 7310 19966 7362 20018
rect 7362 19966 7364 20018
rect 7308 19964 7364 19966
rect 7532 20076 7588 20132
rect 7420 19628 7476 19684
rect 7308 17164 7364 17220
rect 7420 16268 7476 16324
rect 7980 20748 8036 20804
rect 7756 20188 7812 20244
rect 7868 20076 7924 20132
rect 7532 16044 7588 16100
rect 7756 17388 7812 17444
rect 7756 16940 7812 16996
rect 7420 15148 7476 15204
rect 7532 15314 7588 15316
rect 7532 15262 7534 15314
rect 7534 15262 7586 15314
rect 7586 15262 7588 15314
rect 7532 15260 7588 15262
rect 7308 14476 7364 14532
rect 7420 14924 7476 14980
rect 7308 14306 7364 14308
rect 7308 14254 7310 14306
rect 7310 14254 7362 14306
rect 7362 14254 7364 14306
rect 7308 14252 7364 14254
rect 8204 18956 8260 19012
rect 8540 22428 8596 22484
rect 8652 25452 8708 25508
rect 8540 21474 8596 21476
rect 8540 21422 8542 21474
rect 8542 21422 8594 21474
rect 8594 21422 8596 21474
rect 8540 21420 8596 21422
rect 8428 20860 8484 20916
rect 8316 18732 8372 18788
rect 8092 18284 8148 18340
rect 8204 17666 8260 17668
rect 8204 17614 8206 17666
rect 8206 17614 8258 17666
rect 8258 17614 8260 17666
rect 8204 17612 8260 17614
rect 8204 16828 8260 16884
rect 8092 15932 8148 15988
rect 7868 15372 7924 15428
rect 7980 15820 8036 15876
rect 7644 15202 7700 15204
rect 7644 15150 7646 15202
rect 7646 15150 7698 15202
rect 7698 15150 7700 15202
rect 7644 15148 7700 15150
rect 8316 15484 8372 15540
rect 7756 15036 7812 15092
rect 7756 14588 7812 14644
rect 7420 13634 7476 13636
rect 7420 13582 7422 13634
rect 7422 13582 7474 13634
rect 7474 13582 7476 13634
rect 7420 13580 7476 13582
rect 7196 13468 7252 13524
rect 7196 13132 7252 13188
rect 6748 12012 6804 12068
rect 6524 11676 6580 11732
rect 6636 11506 6692 11508
rect 6636 11454 6638 11506
rect 6638 11454 6690 11506
rect 6690 11454 6692 11506
rect 6636 11452 6692 11454
rect 6524 10444 6580 10500
rect 6524 10050 6580 10052
rect 6524 9998 6526 10050
rect 6526 9998 6578 10050
rect 6578 9998 6580 10050
rect 6524 9996 6580 9998
rect 6412 9154 6468 9156
rect 6412 9102 6414 9154
rect 6414 9102 6466 9154
rect 6466 9102 6468 9154
rect 6412 9100 6468 9102
rect 6748 10498 6804 10500
rect 6748 10446 6750 10498
rect 6750 10446 6802 10498
rect 6802 10446 6804 10498
rect 6748 10444 6804 10446
rect 6972 11452 7028 11508
rect 7420 12572 7476 12628
rect 7308 11900 7364 11956
rect 7644 13132 7700 13188
rect 7196 10892 7252 10948
rect 7084 10108 7140 10164
rect 6860 9324 6916 9380
rect 6972 9996 7028 10052
rect 8204 14530 8260 14532
rect 8204 14478 8206 14530
rect 8206 14478 8258 14530
rect 8258 14478 8260 14530
rect 8204 14476 8260 14478
rect 8876 32338 8932 32340
rect 8876 32286 8878 32338
rect 8878 32286 8930 32338
rect 8930 32286 8932 32338
rect 8876 32284 8932 32286
rect 9100 31724 9156 31780
rect 9100 30156 9156 30212
rect 9100 28700 9156 28756
rect 8876 28364 8932 28420
rect 9660 37212 9716 37268
rect 9660 33964 9716 34020
rect 9660 33628 9716 33684
rect 10108 39004 10164 39060
rect 10108 38834 10164 38836
rect 10108 38782 10110 38834
rect 10110 38782 10162 38834
rect 10162 38782 10164 38834
rect 10108 38780 10164 38782
rect 15484 56252 15540 56308
rect 16492 56306 16548 56308
rect 16492 56254 16494 56306
rect 16494 56254 16546 56306
rect 16546 56254 16548 56306
rect 16492 56252 16548 56254
rect 11452 55132 11508 55188
rect 14028 55970 14084 55972
rect 14028 55918 14030 55970
rect 14030 55918 14082 55970
rect 14082 55918 14084 55970
rect 14028 55916 14084 55918
rect 14700 55804 14756 55860
rect 11900 55186 11956 55188
rect 11900 55134 11902 55186
rect 11902 55134 11954 55186
rect 11954 55134 11956 55186
rect 11900 55132 11956 55134
rect 11564 54460 11620 54516
rect 11900 54236 11956 54292
rect 11116 53116 11172 53172
rect 10892 52332 10948 52388
rect 10780 43596 10836 43652
rect 10444 39340 10500 39396
rect 10444 38556 10500 38612
rect 10668 37324 10724 37380
rect 10444 34748 10500 34804
rect 10220 34130 10276 34132
rect 10220 34078 10222 34130
rect 10222 34078 10274 34130
rect 10274 34078 10276 34130
rect 10220 34076 10276 34078
rect 9660 30156 9716 30212
rect 9436 29932 9492 29988
rect 9548 28028 9604 28084
rect 9548 27692 9604 27748
rect 8988 25340 9044 25396
rect 8876 25228 8932 25284
rect 8988 25004 9044 25060
rect 9324 24892 9380 24948
rect 9884 31612 9940 31668
rect 10668 35084 10724 35140
rect 10892 41916 10948 41972
rect 10892 41244 10948 41300
rect 11004 38668 11060 38724
rect 10892 38556 10948 38612
rect 11788 41186 11844 41188
rect 11788 41134 11790 41186
rect 11790 41134 11842 41186
rect 11842 41134 11844 41186
rect 11788 41132 11844 41134
rect 11788 39452 11844 39508
rect 11788 37212 11844 37268
rect 11116 35308 11172 35364
rect 10892 34914 10948 34916
rect 10892 34862 10894 34914
rect 10894 34862 10946 34914
rect 10946 34862 10948 34914
rect 10892 34860 10948 34862
rect 10892 33292 10948 33348
rect 10892 32172 10948 32228
rect 10668 31666 10724 31668
rect 10668 31614 10670 31666
rect 10670 31614 10722 31666
rect 10722 31614 10724 31666
rect 10668 31612 10724 31614
rect 10220 31164 10276 31220
rect 9996 30994 10052 30996
rect 9996 30942 9998 30994
rect 9998 30942 10050 30994
rect 10050 30942 10052 30994
rect 9996 30940 10052 30942
rect 10556 30994 10612 30996
rect 10556 30942 10558 30994
rect 10558 30942 10610 30994
rect 10610 30942 10612 30994
rect 10556 30940 10612 30942
rect 9884 29932 9940 29988
rect 10108 30828 10164 30884
rect 10332 30604 10388 30660
rect 9884 28754 9940 28756
rect 9884 28702 9886 28754
rect 9886 28702 9938 28754
rect 9938 28702 9940 28754
rect 9884 28700 9940 28702
rect 10108 27298 10164 27300
rect 10108 27246 10110 27298
rect 10110 27246 10162 27298
rect 10162 27246 10164 27298
rect 10108 27244 10164 27246
rect 9212 24556 9268 24612
rect 9212 24220 9268 24276
rect 9660 23212 9716 23268
rect 9324 22764 9380 22820
rect 9436 22876 9492 22932
rect 8876 21196 8932 21252
rect 8876 20802 8932 20804
rect 8876 20750 8878 20802
rect 8878 20750 8930 20802
rect 8930 20750 8932 20802
rect 8876 20748 8932 20750
rect 8764 18338 8820 18340
rect 8764 18286 8766 18338
rect 8766 18286 8818 18338
rect 8818 18286 8820 18338
rect 8764 18284 8820 18286
rect 8540 16380 8596 16436
rect 8652 17612 8708 17668
rect 8428 14364 8484 14420
rect 8092 13692 8148 13748
rect 8204 14252 8260 14308
rect 8092 13132 8148 13188
rect 8876 17778 8932 17780
rect 8876 17726 8878 17778
rect 8878 17726 8930 17778
rect 8930 17726 8932 17778
rect 8876 17724 8932 17726
rect 8988 16940 9044 16996
rect 9100 21420 9156 21476
rect 8876 15260 8932 15316
rect 8764 14924 8820 14980
rect 8876 14642 8932 14644
rect 8876 14590 8878 14642
rect 8878 14590 8930 14642
rect 8930 14590 8932 14642
rect 8876 14588 8932 14590
rect 8764 14530 8820 14532
rect 8764 14478 8766 14530
rect 8766 14478 8818 14530
rect 8818 14478 8820 14530
rect 8764 14476 8820 14478
rect 8540 13858 8596 13860
rect 8540 13806 8542 13858
rect 8542 13806 8594 13858
rect 8594 13806 8596 13858
rect 8540 13804 8596 13806
rect 9212 17612 9268 17668
rect 9548 22764 9604 22820
rect 9548 21308 9604 21364
rect 9436 19516 9492 19572
rect 9436 18284 9492 18340
rect 9212 16940 9268 16996
rect 9324 16882 9380 16884
rect 9324 16830 9326 16882
rect 9326 16830 9378 16882
rect 9378 16830 9380 16882
rect 9324 16828 9380 16830
rect 9324 16156 9380 16212
rect 9212 15874 9268 15876
rect 9212 15822 9214 15874
rect 9214 15822 9266 15874
rect 9266 15822 9268 15874
rect 9212 15820 9268 15822
rect 9100 15148 9156 15204
rect 9548 15148 9604 15204
rect 9212 14700 9268 14756
rect 9324 14812 9380 14868
rect 9324 13804 9380 13860
rect 8764 13356 8820 13412
rect 8316 13132 8372 13188
rect 8204 12738 8260 12740
rect 8204 12686 8206 12738
rect 8206 12686 8258 12738
rect 8258 12686 8260 12738
rect 8204 12684 8260 12686
rect 8316 12012 8372 12068
rect 8428 13020 8484 13076
rect 8316 11788 8372 11844
rect 8204 11506 8260 11508
rect 8204 11454 8206 11506
rect 8206 11454 8258 11506
rect 8258 11454 8260 11506
rect 8204 11452 8260 11454
rect 8316 11228 8372 11284
rect 8092 10892 8148 10948
rect 7980 10722 8036 10724
rect 7980 10670 7982 10722
rect 7982 10670 8034 10722
rect 8034 10670 8036 10722
rect 7980 10668 8036 10670
rect 7868 10610 7924 10612
rect 7868 10558 7870 10610
rect 7870 10558 7922 10610
rect 7922 10558 7924 10610
rect 7868 10556 7924 10558
rect 7756 10444 7812 10500
rect 8092 10386 8148 10388
rect 8092 10334 8094 10386
rect 8094 10334 8146 10386
rect 8146 10334 8148 10386
rect 8092 10332 8148 10334
rect 8204 10220 8260 10276
rect 7644 10108 7700 10164
rect 7532 9996 7588 10052
rect 6860 8316 6916 8372
rect 7308 9324 7364 9380
rect 7420 9154 7476 9156
rect 7420 9102 7422 9154
rect 7422 9102 7474 9154
rect 7474 9102 7476 9154
rect 7420 9100 7476 9102
rect 7868 9884 7924 9940
rect 7196 8652 7252 8708
rect 8092 8540 8148 8596
rect 8316 10108 8372 10164
rect 7084 8204 7140 8260
rect 7756 8146 7812 8148
rect 7756 8094 7758 8146
rect 7758 8094 7810 8146
rect 7810 8094 7812 8146
rect 7756 8092 7812 8094
rect 8540 12066 8596 12068
rect 8540 12014 8542 12066
rect 8542 12014 8594 12066
rect 8594 12014 8596 12066
rect 8540 12012 8596 12014
rect 8652 11788 8708 11844
rect 8764 11900 8820 11956
rect 8764 10892 8820 10948
rect 8764 10668 8820 10724
rect 9100 12124 9156 12180
rect 8988 12012 9044 12068
rect 9212 11452 9268 11508
rect 9324 12684 9380 12740
rect 9436 12460 9492 12516
rect 9436 12290 9492 12292
rect 9436 12238 9438 12290
rect 9438 12238 9490 12290
rect 9490 12238 9492 12290
rect 9436 12236 9492 12238
rect 9324 11788 9380 11844
rect 8988 9996 9044 10052
rect 9100 11004 9156 11060
rect 8876 9884 8932 9940
rect 9212 10892 9268 10948
rect 8540 8652 8596 8708
rect 8428 8428 8484 8484
rect 7308 7644 7364 7700
rect 7756 6130 7812 6132
rect 7756 6078 7758 6130
rect 7758 6078 7810 6130
rect 7810 6078 7812 6130
rect 7756 6076 7812 6078
rect 9884 26290 9940 26292
rect 9884 26238 9886 26290
rect 9886 26238 9938 26290
rect 9938 26238 9940 26290
rect 9884 26236 9940 26238
rect 10220 26124 10276 26180
rect 9884 26012 9940 26068
rect 9996 25452 10052 25508
rect 10108 24668 10164 24724
rect 10220 23996 10276 24052
rect 10556 29708 10612 29764
rect 10556 28476 10612 28532
rect 10444 28028 10500 28084
rect 10220 23772 10276 23828
rect 10108 23436 10164 23492
rect 9996 22482 10052 22484
rect 9996 22430 9998 22482
rect 9998 22430 10050 22482
rect 10050 22430 10052 22482
rect 9996 22428 10052 22430
rect 10332 23154 10388 23156
rect 10332 23102 10334 23154
rect 10334 23102 10386 23154
rect 10386 23102 10388 23154
rect 10332 23100 10388 23102
rect 10556 25340 10612 25396
rect 10668 25452 10724 25508
rect 10556 24722 10612 24724
rect 10556 24670 10558 24722
rect 10558 24670 10610 24722
rect 10610 24670 10612 24722
rect 10556 24668 10612 24670
rect 10444 22204 10500 22260
rect 10444 21586 10500 21588
rect 10444 21534 10446 21586
rect 10446 21534 10498 21586
rect 10498 21534 10500 21586
rect 10444 21532 10500 21534
rect 10444 21308 10500 21364
rect 10220 20860 10276 20916
rect 10332 20972 10388 21028
rect 9996 19852 10052 19908
rect 9884 19516 9940 19572
rect 9884 19346 9940 19348
rect 9884 19294 9886 19346
rect 9886 19294 9938 19346
rect 9938 19294 9940 19346
rect 9884 19292 9940 19294
rect 9884 17948 9940 18004
rect 9772 17276 9828 17332
rect 9996 17388 10052 17444
rect 9996 17052 10052 17108
rect 9884 16882 9940 16884
rect 9884 16830 9886 16882
rect 9886 16830 9938 16882
rect 9938 16830 9940 16882
rect 9884 16828 9940 16830
rect 9884 15932 9940 15988
rect 10220 19740 10276 19796
rect 10892 30716 10948 30772
rect 10892 29372 10948 29428
rect 11228 32732 11284 32788
rect 11116 31890 11172 31892
rect 11116 31838 11118 31890
rect 11118 31838 11170 31890
rect 11170 31838 11172 31890
rect 11116 31836 11172 31838
rect 11788 34130 11844 34132
rect 11788 34078 11790 34130
rect 11790 34078 11842 34130
rect 11842 34078 11844 34130
rect 11788 34076 11844 34078
rect 11340 31612 11396 31668
rect 11228 31164 11284 31220
rect 11452 30940 11508 30996
rect 11340 30380 11396 30436
rect 11004 29148 11060 29204
rect 11116 28642 11172 28644
rect 11116 28590 11118 28642
rect 11118 28590 11170 28642
rect 11170 28590 11172 28642
rect 11116 28588 11172 28590
rect 11004 27746 11060 27748
rect 11004 27694 11006 27746
rect 11006 27694 11058 27746
rect 11058 27694 11060 27746
rect 11004 27692 11060 27694
rect 10892 26236 10948 26292
rect 11116 26572 11172 26628
rect 11340 29932 11396 29988
rect 11340 28700 11396 28756
rect 12572 52780 12628 52836
rect 12460 46956 12516 47012
rect 12124 41074 12180 41076
rect 12124 41022 12126 41074
rect 12126 41022 12178 41074
rect 12178 41022 12180 41074
rect 12124 41020 12180 41022
rect 12236 40236 12292 40292
rect 12124 40178 12180 40180
rect 12124 40126 12126 40178
rect 12126 40126 12178 40178
rect 12178 40126 12180 40178
rect 12124 40124 12180 40126
rect 12012 37378 12068 37380
rect 12012 37326 12014 37378
rect 12014 37326 12066 37378
rect 12066 37326 12068 37378
rect 12012 37324 12068 37326
rect 11676 30156 11732 30212
rect 12012 32844 12068 32900
rect 11564 29596 11620 29652
rect 11564 28812 11620 28868
rect 11676 27916 11732 27972
rect 11564 26962 11620 26964
rect 11564 26910 11566 26962
rect 11566 26910 11618 26962
rect 11618 26910 11620 26962
rect 11564 26908 11620 26910
rect 12124 32060 12180 32116
rect 12236 31612 12292 31668
rect 14364 53788 14420 53844
rect 13692 45276 13748 45332
rect 12572 39788 12628 39844
rect 12572 38892 12628 38948
rect 12572 36540 12628 36596
rect 12908 40012 12964 40068
rect 13244 41356 13300 41412
rect 12684 35084 12740 35140
rect 12796 37212 12852 37268
rect 12684 33628 12740 33684
rect 12684 32956 12740 33012
rect 12572 32620 12628 32676
rect 13132 38220 13188 38276
rect 12908 32844 12964 32900
rect 13020 37324 13076 37380
rect 12796 31948 12852 32004
rect 12908 32060 12964 32116
rect 12460 31890 12516 31892
rect 12460 31838 12462 31890
rect 12462 31838 12514 31890
rect 12514 31838 12516 31890
rect 12460 31836 12516 31838
rect 13132 33628 13188 33684
rect 13468 40572 13524 40628
rect 13356 38668 13412 38724
rect 13356 34076 13412 34132
rect 12236 31164 12292 31220
rect 11900 29596 11956 29652
rect 11900 28642 11956 28644
rect 11900 28590 11902 28642
rect 11902 28590 11954 28642
rect 11954 28590 11956 28642
rect 11900 28588 11956 28590
rect 12236 30268 12292 30324
rect 12124 30210 12180 30212
rect 12124 30158 12126 30210
rect 12126 30158 12178 30210
rect 12178 30158 12180 30210
rect 12124 30156 12180 30158
rect 12796 30380 12852 30436
rect 12124 28364 12180 28420
rect 12012 27298 12068 27300
rect 12012 27246 12014 27298
rect 12014 27246 12066 27298
rect 12066 27246 12068 27298
rect 12012 27244 12068 27246
rect 11452 25564 11508 25620
rect 11676 26124 11732 26180
rect 11452 25116 11508 25172
rect 11228 23826 11284 23828
rect 11228 23774 11230 23826
rect 11230 23774 11282 23826
rect 11282 23774 11284 23826
rect 11228 23772 11284 23774
rect 11228 22540 11284 22596
rect 10780 22428 10836 22484
rect 10892 21420 10948 21476
rect 11004 21362 11060 21364
rect 11004 21310 11006 21362
rect 11006 21310 11058 21362
rect 11058 21310 11060 21362
rect 11004 21308 11060 21310
rect 11116 21196 11172 21252
rect 11676 22652 11732 22708
rect 11788 23548 11844 23604
rect 11788 22258 11844 22260
rect 11788 22206 11790 22258
rect 11790 22206 11842 22258
rect 11842 22206 11844 22258
rect 11788 22204 11844 22206
rect 11564 21868 11620 21924
rect 11228 20412 11284 20468
rect 11116 20242 11172 20244
rect 11116 20190 11118 20242
rect 11118 20190 11170 20242
rect 11170 20190 11172 20242
rect 11116 20188 11172 20190
rect 10892 19852 10948 19908
rect 11004 19628 11060 19684
rect 10444 18620 10500 18676
rect 10780 18620 10836 18676
rect 10332 17388 10388 17444
rect 10444 18284 10500 18340
rect 10444 16210 10500 16212
rect 10444 16158 10446 16210
rect 10446 16158 10498 16210
rect 10498 16158 10500 16210
rect 10444 16156 10500 16158
rect 10556 15932 10612 15988
rect 10556 15484 10612 15540
rect 10220 13580 10276 13636
rect 9996 12850 10052 12852
rect 9996 12798 9998 12850
rect 9998 12798 10050 12850
rect 10050 12798 10052 12850
rect 9996 12796 10052 12798
rect 9660 12460 9716 12516
rect 9772 11788 9828 11844
rect 9884 11506 9940 11508
rect 9884 11454 9886 11506
rect 9886 11454 9938 11506
rect 9938 11454 9940 11506
rect 9884 11452 9940 11454
rect 9436 10556 9492 10612
rect 9660 10498 9716 10500
rect 9660 10446 9662 10498
rect 9662 10446 9714 10498
rect 9714 10446 9716 10498
rect 9660 10444 9716 10446
rect 9548 10386 9604 10388
rect 9548 10334 9550 10386
rect 9550 10334 9602 10386
rect 9602 10334 9604 10386
rect 9548 10332 9604 10334
rect 9324 8988 9380 9044
rect 9660 8540 9716 8596
rect 9324 8428 9380 8484
rect 10108 10108 10164 10164
rect 9884 9100 9940 9156
rect 9996 9548 10052 9604
rect 9996 8428 10052 8484
rect 9772 8316 9828 8372
rect 9772 7362 9828 7364
rect 9772 7310 9774 7362
rect 9774 7310 9826 7362
rect 9826 7310 9828 7362
rect 9772 7308 9828 7310
rect 10444 13468 10500 13524
rect 10332 12460 10388 12516
rect 10332 9548 10388 9604
rect 10220 8316 10276 8372
rect 8316 5404 8372 5460
rect 7756 5346 7812 5348
rect 7756 5294 7758 5346
rect 7758 5294 7810 5346
rect 7810 5294 7812 5346
rect 7756 5292 7812 5294
rect 8876 5292 8932 5348
rect 6524 4956 6580 5012
rect 6636 5068 6692 5124
rect 8764 5068 8820 5124
rect 6636 4396 6692 4452
rect 7980 4956 8036 5012
rect 3804 3162 3860 3164
rect 3804 3110 3806 3162
rect 3806 3110 3858 3162
rect 3858 3110 3860 3162
rect 3804 3108 3860 3110
rect 3908 3162 3964 3164
rect 3908 3110 3910 3162
rect 3910 3110 3962 3162
rect 3962 3110 3964 3162
rect 3908 3108 3964 3110
rect 4012 3162 4068 3164
rect 4012 3110 4014 3162
rect 4014 3110 4066 3162
rect 4066 3110 4068 3162
rect 4012 3108 4068 3110
rect 4464 2378 4520 2380
rect 4464 2326 4466 2378
rect 4466 2326 4518 2378
rect 4518 2326 4520 2378
rect 4464 2324 4520 2326
rect 4568 2378 4624 2380
rect 4568 2326 4570 2378
rect 4570 2326 4622 2378
rect 4622 2326 4624 2378
rect 4568 2324 4624 2326
rect 4672 2378 4728 2380
rect 4672 2326 4674 2378
rect 4674 2326 4726 2378
rect 4726 2326 4728 2378
rect 4672 2324 4728 2326
rect 3388 1596 3444 1652
rect 3804 1594 3860 1596
rect 3804 1542 3806 1594
rect 3806 1542 3858 1594
rect 3858 1542 3860 1594
rect 3804 1540 3860 1542
rect 3908 1594 3964 1596
rect 3908 1542 3910 1594
rect 3910 1542 3962 1594
rect 3962 1542 3964 1594
rect 3908 1540 3964 1542
rect 4012 1594 4068 1596
rect 4012 1542 4014 1594
rect 4014 1542 4066 1594
rect 4066 1542 4068 1594
rect 4012 1540 4068 1542
rect 4464 810 4520 812
rect 4464 758 4466 810
rect 4466 758 4518 810
rect 4518 758 4520 810
rect 4464 756 4520 758
rect 4568 810 4624 812
rect 4568 758 4570 810
rect 4570 758 4622 810
rect 4622 758 4624 810
rect 4568 756 4624 758
rect 4672 810 4728 812
rect 4672 758 4674 810
rect 4674 758 4726 810
rect 4726 758 4728 810
rect 4672 756 4728 758
rect 4732 364 4788 420
rect 10444 9042 10500 9044
rect 10444 8990 10446 9042
rect 10446 8990 10498 9042
rect 10498 8990 10500 9042
rect 10444 8988 10500 8990
rect 10892 15202 10948 15204
rect 10892 15150 10894 15202
rect 10894 15150 10946 15202
rect 10946 15150 10948 15202
rect 10892 15148 10948 15150
rect 11116 17948 11172 18004
rect 11116 17388 11172 17444
rect 11116 17052 11172 17108
rect 11452 17948 11508 18004
rect 11676 18172 11732 18228
rect 10780 12460 10836 12516
rect 11116 11676 11172 11732
rect 10668 10668 10724 10724
rect 10892 10892 10948 10948
rect 10892 10332 10948 10388
rect 11116 11004 11172 11060
rect 11116 10668 11172 10724
rect 11340 13580 11396 13636
rect 11564 17442 11620 17444
rect 11564 17390 11566 17442
rect 11566 17390 11618 17442
rect 11618 17390 11620 17442
rect 11564 17388 11620 17390
rect 11676 13356 11732 13412
rect 11676 13020 11732 13076
rect 11340 11004 11396 11060
rect 11452 11676 11508 11732
rect 11228 10386 11284 10388
rect 11228 10334 11230 10386
rect 11230 10334 11282 10386
rect 11282 10334 11284 10386
rect 11228 10332 11284 10334
rect 11676 11394 11732 11396
rect 11676 11342 11678 11394
rect 11678 11342 11730 11394
rect 11730 11342 11732 11394
rect 11676 11340 11732 11342
rect 11564 10892 11620 10948
rect 11676 11116 11732 11172
rect 11788 11004 11844 11060
rect 12012 26796 12068 26852
rect 12012 25004 12068 25060
rect 12684 28252 12740 28308
rect 12908 30044 12964 30100
rect 13020 28364 13076 28420
rect 13244 32508 13300 32564
rect 13580 38834 13636 38836
rect 13580 38782 13582 38834
rect 13582 38782 13634 38834
rect 13634 38782 13636 38834
rect 13580 38780 13636 38782
rect 13580 38444 13636 38500
rect 13580 37154 13636 37156
rect 13580 37102 13582 37154
rect 13582 37102 13634 37154
rect 13634 37102 13636 37154
rect 13580 37100 13636 37102
rect 13468 32060 13524 32116
rect 13356 31948 13412 32004
rect 13580 31612 13636 31668
rect 13468 31276 13524 31332
rect 13580 30828 13636 30884
rect 13356 30268 13412 30324
rect 12908 27244 12964 27300
rect 12460 26348 12516 26404
rect 12684 25676 12740 25732
rect 12236 24162 12292 24164
rect 12236 24110 12238 24162
rect 12238 24110 12290 24162
rect 12290 24110 12292 24162
rect 12236 24108 12292 24110
rect 12572 23884 12628 23940
rect 12236 22594 12292 22596
rect 12236 22542 12238 22594
rect 12238 22542 12290 22594
rect 12290 22542 12292 22594
rect 12236 22540 12292 22542
rect 12124 21868 12180 21924
rect 12124 21586 12180 21588
rect 12124 21534 12126 21586
rect 12126 21534 12178 21586
rect 12178 21534 12180 21586
rect 12124 21532 12180 21534
rect 12348 21084 12404 21140
rect 12460 20412 12516 20468
rect 12908 25452 12964 25508
rect 12796 24108 12852 24164
rect 13132 27298 13188 27300
rect 13132 27246 13134 27298
rect 13134 27246 13186 27298
rect 13186 27246 13188 27298
rect 13132 27244 13188 27246
rect 13580 28642 13636 28644
rect 13580 28590 13582 28642
rect 13582 28590 13634 28642
rect 13634 28590 13636 28642
rect 13580 28588 13636 28590
rect 13580 28252 13636 28308
rect 13580 27692 13636 27748
rect 13356 26460 13412 26516
rect 13132 25676 13188 25732
rect 13244 25788 13300 25844
rect 13132 25452 13188 25508
rect 12684 19628 12740 19684
rect 12796 19964 12852 20020
rect 12572 19516 12628 19572
rect 12796 19404 12852 19460
rect 12012 19068 12068 19124
rect 12460 19122 12516 19124
rect 12460 19070 12462 19122
rect 12462 19070 12514 19122
rect 12514 19070 12516 19122
rect 12460 19068 12516 19070
rect 13244 25340 13300 25396
rect 13916 41074 13972 41076
rect 13916 41022 13918 41074
rect 13918 41022 13970 41074
rect 13970 41022 13972 41074
rect 13916 41020 13972 41022
rect 13916 38780 13972 38836
rect 13804 38722 13860 38724
rect 13804 38670 13806 38722
rect 13806 38670 13858 38722
rect 13858 38670 13860 38722
rect 13804 38668 13860 38670
rect 13804 36988 13860 37044
rect 13804 32508 13860 32564
rect 14700 41916 14756 41972
rect 14364 41468 14420 41524
rect 19516 57260 19572 57316
rect 19852 57260 19908 57316
rect 20860 56252 20916 56308
rect 22204 56306 22260 56308
rect 22204 56254 22206 56306
rect 22206 56254 22258 56306
rect 22258 56254 22260 56306
rect 22204 56252 22260 56254
rect 22540 56140 22596 56196
rect 16828 53676 16884 53732
rect 16044 50428 16100 50484
rect 15596 41692 15652 41748
rect 15708 45836 15764 45892
rect 15036 41356 15092 41412
rect 14364 41020 14420 41076
rect 14140 39228 14196 39284
rect 14252 40124 14308 40180
rect 14476 39452 14532 39508
rect 14588 40348 14644 40404
rect 14140 32060 14196 32116
rect 13916 31164 13972 31220
rect 13916 30604 13972 30660
rect 14028 30210 14084 30212
rect 14028 30158 14030 30210
rect 14030 30158 14082 30210
rect 14082 30158 14084 30210
rect 14028 30156 14084 30158
rect 14476 31778 14532 31780
rect 14476 31726 14478 31778
rect 14478 31726 14530 31778
rect 14530 31726 14532 31778
rect 14476 31724 14532 31726
rect 14364 30828 14420 30884
rect 14252 30156 14308 30212
rect 13916 28924 13972 28980
rect 13804 28700 13860 28756
rect 13916 28588 13972 28644
rect 14812 38834 14868 38836
rect 14812 38782 14814 38834
rect 14814 38782 14866 38834
rect 14866 38782 14868 38834
rect 14812 38780 14868 38782
rect 14924 38444 14980 38500
rect 14588 30716 14644 30772
rect 14364 29820 14420 29876
rect 14924 32172 14980 32228
rect 13916 27244 13972 27300
rect 14140 27186 14196 27188
rect 14140 27134 14142 27186
rect 14142 27134 14194 27186
rect 14194 27134 14196 27186
rect 14140 27132 14196 27134
rect 13916 27020 13972 27076
rect 13692 25116 13748 25172
rect 13804 25900 13860 25956
rect 13692 24892 13748 24948
rect 13468 23938 13524 23940
rect 13468 23886 13470 23938
rect 13470 23886 13522 23938
rect 13522 23886 13524 23938
rect 13468 23884 13524 23886
rect 13580 24668 13636 24724
rect 13356 22764 13412 22820
rect 13468 23324 13524 23380
rect 13356 22594 13412 22596
rect 13356 22542 13358 22594
rect 13358 22542 13410 22594
rect 13410 22542 13412 22594
rect 13356 22540 13412 22542
rect 13468 22316 13524 22372
rect 13356 21980 13412 22036
rect 13132 20300 13188 20356
rect 13132 20018 13188 20020
rect 13132 19966 13134 20018
rect 13134 19966 13186 20018
rect 13186 19966 13188 20018
rect 13132 19964 13188 19966
rect 13804 23660 13860 23716
rect 13692 23324 13748 23380
rect 14252 26908 14308 26964
rect 13244 19234 13300 19236
rect 13244 19182 13246 19234
rect 13246 19182 13298 19234
rect 13298 19182 13300 19234
rect 13244 19180 13300 19182
rect 14028 26684 14084 26740
rect 13692 19852 13748 19908
rect 14252 25900 14308 25956
rect 14700 26908 14756 26964
rect 15260 38780 15316 38836
rect 15148 38556 15204 38612
rect 15036 32060 15092 32116
rect 15148 31948 15204 32004
rect 15036 30882 15092 30884
rect 15036 30830 15038 30882
rect 15038 30830 15090 30882
rect 15090 30830 15092 30882
rect 15036 30828 15092 30830
rect 15148 29426 15204 29428
rect 15148 29374 15150 29426
rect 15150 29374 15202 29426
rect 15202 29374 15204 29426
rect 15148 29372 15204 29374
rect 15596 39116 15652 39172
rect 15820 38834 15876 38836
rect 15820 38782 15822 38834
rect 15822 38782 15874 38834
rect 15874 38782 15876 38834
rect 15820 38780 15876 38782
rect 16828 46956 16884 47012
rect 17276 53564 17332 53620
rect 16940 46060 16996 46116
rect 16044 40460 16100 40516
rect 16716 41804 16772 41860
rect 15932 37266 15988 37268
rect 15932 37214 15934 37266
rect 15934 37214 15986 37266
rect 15986 37214 15988 37266
rect 15932 37212 15988 37214
rect 15596 34748 15652 34804
rect 15596 32674 15652 32676
rect 15596 32622 15598 32674
rect 15598 32622 15650 32674
rect 15650 32622 15652 32674
rect 15596 32620 15652 32622
rect 15820 32284 15876 32340
rect 15708 30940 15764 30996
rect 15932 31948 15988 32004
rect 15484 29596 15540 29652
rect 15484 29372 15540 29428
rect 14588 26236 14644 26292
rect 14140 24668 14196 24724
rect 14588 26012 14644 26068
rect 14476 25394 14532 25396
rect 14476 25342 14478 25394
rect 14478 25342 14530 25394
rect 14530 25342 14532 25394
rect 14476 25340 14532 25342
rect 14924 25730 14980 25732
rect 14924 25678 14926 25730
rect 14926 25678 14978 25730
rect 14978 25678 14980 25730
rect 14924 25676 14980 25678
rect 14364 24444 14420 24500
rect 14476 21420 14532 21476
rect 14364 20802 14420 20804
rect 14364 20750 14366 20802
rect 14366 20750 14418 20802
rect 14418 20750 14420 20802
rect 14364 20748 14420 20750
rect 14700 23154 14756 23156
rect 14700 23102 14702 23154
rect 14702 23102 14754 23154
rect 14754 23102 14756 23154
rect 14700 23100 14756 23102
rect 14812 22482 14868 22484
rect 14812 22430 14814 22482
rect 14814 22430 14866 22482
rect 14866 22430 14868 22482
rect 14812 22428 14868 22430
rect 14812 21586 14868 21588
rect 14812 21534 14814 21586
rect 14814 21534 14866 21586
rect 14866 21534 14868 21586
rect 14812 21532 14868 21534
rect 15708 29372 15764 29428
rect 15708 28812 15764 28868
rect 15260 26290 15316 26292
rect 15260 26238 15262 26290
rect 15262 26238 15314 26290
rect 15314 26238 15316 26290
rect 15260 26236 15316 26238
rect 15372 24722 15428 24724
rect 15372 24670 15374 24722
rect 15374 24670 15426 24722
rect 15426 24670 15428 24722
rect 15372 24668 15428 24670
rect 15148 23660 15204 23716
rect 15596 26908 15652 26964
rect 15596 25116 15652 25172
rect 15820 26178 15876 26180
rect 15820 26126 15822 26178
rect 15822 26126 15874 26178
rect 15874 26126 15876 26178
rect 15820 26124 15876 26126
rect 15820 25004 15876 25060
rect 15260 24332 15316 24388
rect 15148 23324 15204 23380
rect 15596 24108 15652 24164
rect 15372 23660 15428 23716
rect 15372 22204 15428 22260
rect 15372 21980 15428 22036
rect 14700 20188 14756 20244
rect 14924 20748 14980 20804
rect 14140 19964 14196 20020
rect 13580 19180 13636 19236
rect 14028 19852 14084 19908
rect 14028 19628 14084 19684
rect 12124 18732 12180 18788
rect 13356 18620 13412 18676
rect 12124 17052 12180 17108
rect 12572 16604 12628 16660
rect 12124 16492 12180 16548
rect 12572 15484 12628 15540
rect 12460 15260 12516 15316
rect 12012 14476 12068 14532
rect 12460 14476 12516 14532
rect 12012 14140 12068 14196
rect 12012 12460 12068 12516
rect 12908 18284 12964 18340
rect 12796 16828 12852 16884
rect 13356 18338 13412 18340
rect 13356 18286 13358 18338
rect 13358 18286 13410 18338
rect 13410 18286 13412 18338
rect 13356 18284 13412 18286
rect 13580 16716 13636 16772
rect 13468 15820 13524 15876
rect 13132 14418 13188 14420
rect 13132 14366 13134 14418
rect 13134 14366 13186 14418
rect 13186 14366 13188 14418
rect 13132 14364 13188 14366
rect 12796 13468 12852 13524
rect 12684 13356 12740 13412
rect 12908 13356 12964 13412
rect 12684 13074 12740 13076
rect 12684 13022 12686 13074
rect 12686 13022 12738 13074
rect 12738 13022 12740 13074
rect 12684 13020 12740 13022
rect 12572 12796 12628 12852
rect 12236 12236 12292 12292
rect 11452 10220 11508 10276
rect 11340 9100 11396 9156
rect 10892 8764 10948 8820
rect 11116 8370 11172 8372
rect 11116 8318 11118 8370
rect 11118 8318 11170 8370
rect 11170 8318 11172 8370
rect 11116 8316 11172 8318
rect 10668 7308 10724 7364
rect 11004 7308 11060 7364
rect 11004 6748 11060 6804
rect 11676 10108 11732 10164
rect 11564 8652 11620 8708
rect 11228 7196 11284 7252
rect 11564 6690 11620 6692
rect 11564 6638 11566 6690
rect 11566 6638 11618 6690
rect 11618 6638 11620 6690
rect 11564 6636 11620 6638
rect 11116 5292 11172 5348
rect 11564 5292 11620 5348
rect 11564 4508 11620 4564
rect 12124 10780 12180 10836
rect 12236 10556 12292 10612
rect 11900 9884 11956 9940
rect 12012 10444 12068 10500
rect 12348 10220 12404 10276
rect 12124 9884 12180 9940
rect 12236 9436 12292 9492
rect 12348 9548 12404 9604
rect 12124 8930 12180 8932
rect 12124 8878 12126 8930
rect 12126 8878 12178 8930
rect 12178 8878 12180 8930
rect 12124 8876 12180 8878
rect 12348 8876 12404 8932
rect 12460 9212 12516 9268
rect 12796 12460 12852 12516
rect 12796 10780 12852 10836
rect 12796 9042 12852 9044
rect 12796 8990 12798 9042
rect 12798 8990 12850 9042
rect 12850 8990 12852 9042
rect 12796 8988 12852 8990
rect 13244 13356 13300 13412
rect 13020 12796 13076 12852
rect 13020 11116 13076 11172
rect 13356 11676 13412 11732
rect 13244 11116 13300 11172
rect 14476 18956 14532 19012
rect 15148 20300 15204 20356
rect 14924 19964 14980 20020
rect 15036 19852 15092 19908
rect 14924 19628 14980 19684
rect 14140 16604 14196 16660
rect 14700 16940 14756 16996
rect 14476 16380 14532 16436
rect 13804 16044 13860 16100
rect 14364 15932 14420 15988
rect 14476 15484 14532 15540
rect 14700 15202 14756 15204
rect 14700 15150 14702 15202
rect 14702 15150 14754 15202
rect 14754 15150 14756 15202
rect 14700 15148 14756 15150
rect 15372 20972 15428 21028
rect 15036 16882 15092 16884
rect 15036 16830 15038 16882
rect 15038 16830 15090 16882
rect 15090 16830 15092 16882
rect 15036 16828 15092 16830
rect 15036 15874 15092 15876
rect 15036 15822 15038 15874
rect 15038 15822 15090 15874
rect 15090 15822 15092 15874
rect 15036 15820 15092 15822
rect 15148 15314 15204 15316
rect 15148 15262 15150 15314
rect 15150 15262 15202 15314
rect 15202 15262 15204 15314
rect 15148 15260 15204 15262
rect 13804 13580 13860 13636
rect 14364 14364 14420 14420
rect 13916 12684 13972 12740
rect 14028 13468 14084 13524
rect 13692 12460 13748 12516
rect 13244 10722 13300 10724
rect 13244 10670 13246 10722
rect 13246 10670 13298 10722
rect 13298 10670 13300 10722
rect 13244 10668 13300 10670
rect 13020 10610 13076 10612
rect 13020 10558 13022 10610
rect 13022 10558 13074 10610
rect 13074 10558 13076 10610
rect 13020 10556 13076 10558
rect 13132 9938 13188 9940
rect 13132 9886 13134 9938
rect 13134 9886 13186 9938
rect 13186 9886 13188 9938
rect 13132 9884 13188 9886
rect 13244 9212 13300 9268
rect 12908 8316 12964 8372
rect 14364 13468 14420 13524
rect 14700 14642 14756 14644
rect 14700 14590 14702 14642
rect 14702 14590 14754 14642
rect 14754 14590 14756 14642
rect 14700 14588 14756 14590
rect 13356 8540 13412 8596
rect 13468 8316 13524 8372
rect 13692 10386 13748 10388
rect 13692 10334 13694 10386
rect 13694 10334 13746 10386
rect 13746 10334 13748 10386
rect 13692 10332 13748 10334
rect 14028 10556 14084 10612
rect 13804 9884 13860 9940
rect 14028 9602 14084 9604
rect 14028 9550 14030 9602
rect 14030 9550 14082 9602
rect 14082 9550 14084 9602
rect 14028 9548 14084 9550
rect 13580 7420 13636 7476
rect 13916 8428 13972 8484
rect 13020 6972 13076 7028
rect 12684 6802 12740 6804
rect 12684 6750 12686 6802
rect 12686 6750 12738 6802
rect 12738 6750 12740 6802
rect 12684 6748 12740 6750
rect 12236 5852 12292 5908
rect 13244 7084 13300 7140
rect 13356 6972 13412 7028
rect 14700 13916 14756 13972
rect 14812 13468 14868 13524
rect 14924 12348 14980 12404
rect 14812 10556 14868 10612
rect 14588 9996 14644 10052
rect 14252 8204 14308 8260
rect 13804 5346 13860 5348
rect 13804 5294 13806 5346
rect 13806 5294 13858 5346
rect 13858 5294 13860 5346
rect 13804 5292 13860 5294
rect 14588 7474 14644 7476
rect 14588 7422 14590 7474
rect 14590 7422 14642 7474
rect 14642 7422 14644 7474
rect 14588 7420 14644 7422
rect 15148 13916 15204 13972
rect 15260 13692 15316 13748
rect 15596 20748 15652 20804
rect 15484 19234 15540 19236
rect 15484 19182 15486 19234
rect 15486 19182 15538 19234
rect 15538 19182 15540 19234
rect 15484 19180 15540 19182
rect 16156 36652 16212 36708
rect 16268 34860 16324 34916
rect 16380 32172 16436 32228
rect 16492 37100 16548 37156
rect 17164 37324 17220 37380
rect 16716 36706 16772 36708
rect 16716 36654 16718 36706
rect 16718 36654 16770 36706
rect 16770 36654 16772 36706
rect 16716 36652 16772 36654
rect 16604 35196 16660 35252
rect 17388 39004 17444 39060
rect 16044 28642 16100 28644
rect 16044 28590 16046 28642
rect 16046 28590 16098 28642
rect 16098 28590 16100 28642
rect 16044 28588 16100 28590
rect 17052 34636 17108 34692
rect 16828 31724 16884 31780
rect 16268 26796 16324 26852
rect 16044 24444 16100 24500
rect 16380 29426 16436 29428
rect 16380 29374 16382 29426
rect 16382 29374 16434 29426
rect 16434 29374 16436 29426
rect 16380 29372 16436 29374
rect 16268 23378 16324 23380
rect 16268 23326 16270 23378
rect 16270 23326 16322 23378
rect 16322 23326 16324 23378
rect 16268 23324 16324 23326
rect 16044 21868 16100 21924
rect 16156 22092 16212 22148
rect 15932 20972 15988 21028
rect 16044 21196 16100 21252
rect 16268 20748 16324 20804
rect 16492 28812 16548 28868
rect 16716 29596 16772 29652
rect 16604 27858 16660 27860
rect 16604 27806 16606 27858
rect 16606 27806 16658 27858
rect 16658 27806 16660 27858
rect 16604 27804 16660 27806
rect 16604 27468 16660 27524
rect 16716 27132 16772 27188
rect 16940 30882 16996 30884
rect 16940 30830 16942 30882
rect 16942 30830 16994 30882
rect 16994 30830 16996 30882
rect 16940 30828 16996 30830
rect 17276 35756 17332 35812
rect 18284 55298 18340 55300
rect 18284 55246 18286 55298
rect 18286 55246 18338 55298
rect 18338 55246 18340 55298
rect 18284 55244 18340 55246
rect 17500 37324 17556 37380
rect 17948 46508 18004 46564
rect 17500 36540 17556 36596
rect 17500 35308 17556 35364
rect 19628 55916 19684 55972
rect 21308 55970 21364 55972
rect 21308 55918 21310 55970
rect 21310 55918 21362 55970
rect 21362 55918 21364 55970
rect 21308 55916 21364 55918
rect 21644 55804 21700 55860
rect 20524 55298 20580 55300
rect 20524 55246 20526 55298
rect 20526 55246 20578 55298
rect 20578 55246 20580 55298
rect 20524 55244 20580 55246
rect 20636 54290 20692 54292
rect 20636 54238 20638 54290
rect 20638 54238 20690 54290
rect 20690 54238 20692 54290
rect 20636 54236 20692 54238
rect 21196 54514 21252 54516
rect 21196 54462 21198 54514
rect 21198 54462 21250 54514
rect 21250 54462 21252 54514
rect 21196 54460 21252 54462
rect 20860 53788 20916 53844
rect 21420 52162 21476 52164
rect 21420 52110 21422 52162
rect 21422 52110 21474 52162
rect 21474 52110 21476 52162
rect 21420 52108 21476 52110
rect 19964 48076 20020 48132
rect 19740 47292 19796 47348
rect 18396 40124 18452 40180
rect 18060 35308 18116 35364
rect 17836 34188 17892 34244
rect 17052 30210 17108 30212
rect 17052 30158 17054 30210
rect 17054 30158 17106 30210
rect 17106 30158 17108 30210
rect 17052 30156 17108 30158
rect 16940 29484 16996 29540
rect 17052 29820 17108 29876
rect 17724 33740 17780 33796
rect 17500 33628 17556 33684
rect 17500 30492 17556 30548
rect 17836 33628 17892 33684
rect 17724 30268 17780 30324
rect 18060 31948 18116 32004
rect 17388 29932 17444 29988
rect 17724 29932 17780 29988
rect 17388 28530 17444 28532
rect 17388 28478 17390 28530
rect 17390 28478 17442 28530
rect 17442 28478 17444 28530
rect 17388 28476 17444 28478
rect 17164 27580 17220 27636
rect 17388 27186 17444 27188
rect 17388 27134 17390 27186
rect 17390 27134 17442 27186
rect 17442 27134 17444 27186
rect 17388 27132 17444 27134
rect 17052 26348 17108 26404
rect 17500 26684 17556 26740
rect 16828 26012 16884 26068
rect 17276 25676 17332 25732
rect 17388 26012 17444 26068
rect 18060 31778 18116 31780
rect 18060 31726 18062 31778
rect 18062 31726 18114 31778
rect 18114 31726 18116 31778
rect 18060 31724 18116 31726
rect 17948 28812 18004 28868
rect 18060 29260 18116 29316
rect 17836 27804 17892 27860
rect 17500 25564 17556 25620
rect 18284 36594 18340 36596
rect 18284 36542 18286 36594
rect 18286 36542 18338 36594
rect 18338 36542 18340 36594
rect 18284 36540 18340 36542
rect 18284 34802 18340 34804
rect 18284 34750 18286 34802
rect 18286 34750 18338 34802
rect 18338 34750 18340 34802
rect 18284 34748 18340 34750
rect 18284 33740 18340 33796
rect 18172 27804 18228 27860
rect 18060 27580 18116 27636
rect 19068 34914 19124 34916
rect 19068 34862 19070 34914
rect 19070 34862 19122 34914
rect 19122 34862 19124 34914
rect 19068 34860 19124 34862
rect 19404 36258 19460 36260
rect 19404 36206 19406 36258
rect 19406 36206 19458 36258
rect 19458 36206 19460 36258
rect 19404 36204 19460 36206
rect 18732 33516 18788 33572
rect 19292 33516 19348 33572
rect 18508 31948 18564 32004
rect 18396 31724 18452 31780
rect 18508 30994 18564 30996
rect 18508 30942 18510 30994
rect 18510 30942 18562 30994
rect 18562 30942 18564 30994
rect 18508 30940 18564 30942
rect 18508 30492 18564 30548
rect 18620 29986 18676 29988
rect 18620 29934 18622 29986
rect 18622 29934 18674 29986
rect 18674 29934 18676 29986
rect 18620 29932 18676 29934
rect 18508 28812 18564 28868
rect 18956 33180 19012 33236
rect 20188 44268 20244 44324
rect 19852 41916 19908 41972
rect 20076 41244 20132 41300
rect 19964 38668 20020 38724
rect 19852 36204 19908 36260
rect 19964 34412 20020 34468
rect 21084 40012 21140 40068
rect 20748 37996 20804 38052
rect 20188 35644 20244 35700
rect 19740 30940 19796 30996
rect 19964 31052 20020 31108
rect 19292 30210 19348 30212
rect 19292 30158 19294 30210
rect 19294 30158 19346 30210
rect 19346 30158 19348 30210
rect 19292 30156 19348 30158
rect 18956 29932 19012 29988
rect 19068 30044 19124 30100
rect 18844 29148 18900 29204
rect 18732 28364 18788 28420
rect 18284 26012 18340 26068
rect 18396 26402 18452 26404
rect 18396 26350 18398 26402
rect 18398 26350 18450 26402
rect 18450 26350 18452 26402
rect 18396 26348 18452 26350
rect 18732 25676 18788 25732
rect 18956 25676 19012 25732
rect 16828 24108 16884 24164
rect 17388 24332 17444 24388
rect 17164 23996 17220 24052
rect 16716 23826 16772 23828
rect 16716 23774 16718 23826
rect 16718 23774 16770 23826
rect 16770 23774 16772 23826
rect 16716 23772 16772 23774
rect 17052 23324 17108 23380
rect 16828 22146 16884 22148
rect 16828 22094 16830 22146
rect 16830 22094 16882 22146
rect 16882 22094 16884 22146
rect 16828 22092 16884 22094
rect 15820 19516 15876 19572
rect 16268 20524 16324 20580
rect 15820 19180 15876 19236
rect 15932 19292 15988 19348
rect 15820 17276 15876 17332
rect 15820 17052 15876 17108
rect 15148 13634 15204 13636
rect 15148 13582 15150 13634
rect 15150 13582 15202 13634
rect 15202 13582 15204 13634
rect 15148 13580 15204 13582
rect 15596 11618 15652 11620
rect 15596 11566 15598 11618
rect 15598 11566 15650 11618
rect 15650 11566 15652 11618
rect 15596 11564 15652 11566
rect 15036 9996 15092 10052
rect 15148 10108 15204 10164
rect 15148 9660 15204 9716
rect 14924 8428 14980 8484
rect 14812 8204 14868 8260
rect 14812 7868 14868 7924
rect 15372 9660 15428 9716
rect 16044 19068 16100 19124
rect 16156 19010 16212 19012
rect 16156 18958 16158 19010
rect 16158 18958 16210 19010
rect 16210 18958 16212 19010
rect 16156 18956 16212 18958
rect 16044 18844 16100 18900
rect 16156 17388 16212 17444
rect 16268 17052 16324 17108
rect 16156 15820 16212 15876
rect 16044 12908 16100 12964
rect 16156 12236 16212 12292
rect 17500 24220 17556 24276
rect 17500 23660 17556 23716
rect 17388 22092 17444 22148
rect 17500 21756 17556 21812
rect 17052 21308 17108 21364
rect 17388 21532 17444 21588
rect 16492 20018 16548 20020
rect 16492 19966 16494 20018
rect 16494 19966 16546 20018
rect 16546 19966 16548 20018
rect 16492 19964 16548 19966
rect 17276 21196 17332 21252
rect 18396 25340 18452 25396
rect 19740 30044 19796 30100
rect 20188 30828 20244 30884
rect 20524 31500 20580 31556
rect 20636 30882 20692 30884
rect 20636 30830 20638 30882
rect 20638 30830 20690 30882
rect 20690 30830 20692 30882
rect 20636 30828 20692 30830
rect 20412 30156 20468 30212
rect 20076 30044 20132 30100
rect 19292 29932 19348 29988
rect 19180 28476 19236 28532
rect 19068 23996 19124 24052
rect 18284 23660 18340 23716
rect 18060 22540 18116 22596
rect 18396 23100 18452 23156
rect 17948 22482 18004 22484
rect 17948 22430 17950 22482
rect 17950 22430 18002 22482
rect 18002 22430 18004 22482
rect 17948 22428 18004 22430
rect 18396 22092 18452 22148
rect 18284 21756 18340 21812
rect 17388 19234 17444 19236
rect 17388 19182 17390 19234
rect 17390 19182 17442 19234
rect 17442 19182 17444 19234
rect 17388 19180 17444 19182
rect 17164 18956 17220 19012
rect 16828 17890 16884 17892
rect 16828 17838 16830 17890
rect 16830 17838 16882 17890
rect 16882 17838 16884 17890
rect 16828 17836 16884 17838
rect 16716 17666 16772 17668
rect 16716 17614 16718 17666
rect 16718 17614 16770 17666
rect 16770 17614 16772 17666
rect 16716 17612 16772 17614
rect 16940 17276 16996 17332
rect 16492 15148 16548 15204
rect 16940 16098 16996 16100
rect 16940 16046 16942 16098
rect 16942 16046 16994 16098
rect 16994 16046 16996 16098
rect 16940 16044 16996 16046
rect 17500 18844 17556 18900
rect 17612 19852 17668 19908
rect 17388 18338 17444 18340
rect 17388 18286 17390 18338
rect 17390 18286 17442 18338
rect 17442 18286 17444 18338
rect 17388 18284 17444 18286
rect 17948 21026 18004 21028
rect 17948 20974 17950 21026
rect 17950 20974 18002 21026
rect 18002 20974 18004 21026
rect 17948 20972 18004 20974
rect 17836 19852 17892 19908
rect 17500 17778 17556 17780
rect 17500 17726 17502 17778
rect 17502 17726 17554 17778
rect 17554 17726 17556 17778
rect 17500 17724 17556 17726
rect 17276 17612 17332 17668
rect 17388 17052 17444 17108
rect 17276 16828 17332 16884
rect 17388 16380 17444 16436
rect 17276 16156 17332 16212
rect 17164 15820 17220 15876
rect 16828 15260 16884 15316
rect 17052 14924 17108 14980
rect 17052 14588 17108 14644
rect 16716 14530 16772 14532
rect 16716 14478 16718 14530
rect 16718 14478 16770 14530
rect 16770 14478 16772 14530
rect 16716 14476 16772 14478
rect 16604 13916 16660 13972
rect 16828 14364 16884 14420
rect 16492 12178 16548 12180
rect 16492 12126 16494 12178
rect 16494 12126 16546 12178
rect 16546 12126 16548 12178
rect 16492 12124 16548 12126
rect 17500 15036 17556 15092
rect 17164 14028 17220 14084
rect 17276 14924 17332 14980
rect 17164 12738 17220 12740
rect 17164 12686 17166 12738
rect 17166 12686 17218 12738
rect 17218 12686 17220 12738
rect 17164 12684 17220 12686
rect 16380 11564 16436 11620
rect 17052 11900 17108 11956
rect 15596 9660 15652 9716
rect 15484 9602 15540 9604
rect 15484 9550 15486 9602
rect 15486 9550 15538 9602
rect 15538 9550 15540 9602
rect 15484 9548 15540 9550
rect 15708 9548 15764 9604
rect 15372 8818 15428 8820
rect 15372 8766 15374 8818
rect 15374 8766 15426 8818
rect 15426 8766 15428 8818
rect 15372 8764 15428 8766
rect 15596 8370 15652 8372
rect 15596 8318 15598 8370
rect 15598 8318 15650 8370
rect 15650 8318 15652 8370
rect 15596 8316 15652 8318
rect 15260 8204 15316 8260
rect 15036 8034 15092 8036
rect 15036 7982 15038 8034
rect 15038 7982 15090 8034
rect 15090 7982 15092 8034
rect 15036 7980 15092 7982
rect 15372 7980 15428 8036
rect 15484 7420 15540 7476
rect 14924 7308 14980 7364
rect 15596 7362 15652 7364
rect 15596 7310 15598 7362
rect 15598 7310 15650 7362
rect 15650 7310 15652 7362
rect 15596 7308 15652 7310
rect 15708 7250 15764 7252
rect 15708 7198 15710 7250
rect 15710 7198 15762 7250
rect 15762 7198 15764 7250
rect 15708 7196 15764 7198
rect 16044 10108 16100 10164
rect 16268 10108 16324 10164
rect 16492 9996 16548 10052
rect 16044 9660 16100 9716
rect 14812 5682 14868 5684
rect 14812 5630 14814 5682
rect 14814 5630 14866 5682
rect 14866 5630 14868 5682
rect 14812 5628 14868 5630
rect 14476 5292 14532 5348
rect 15372 5628 15428 5684
rect 16156 9436 16212 9492
rect 16604 9548 16660 9604
rect 17164 11452 17220 11508
rect 16828 11228 16884 11284
rect 17388 13970 17444 13972
rect 17388 13918 17390 13970
rect 17390 13918 17442 13970
rect 17442 13918 17444 13970
rect 17388 13916 17444 13918
rect 17276 10780 17332 10836
rect 17388 12908 17444 12964
rect 18172 18620 18228 18676
rect 18060 17388 18116 17444
rect 18284 18284 18340 18340
rect 18284 17388 18340 17444
rect 18284 17106 18340 17108
rect 18284 17054 18286 17106
rect 18286 17054 18338 17106
rect 18338 17054 18340 17106
rect 18284 17052 18340 17054
rect 17948 16380 18004 16436
rect 17724 15596 17780 15652
rect 17836 15148 17892 15204
rect 18284 16098 18340 16100
rect 18284 16046 18286 16098
rect 18286 16046 18338 16098
rect 18338 16046 18340 16098
rect 18284 16044 18340 16046
rect 18508 21196 18564 21252
rect 18956 23938 19012 23940
rect 18956 23886 18958 23938
rect 18958 23886 19010 23938
rect 19010 23886 19012 23938
rect 18956 23884 19012 23886
rect 19404 23884 19460 23940
rect 20188 26796 20244 26852
rect 19068 22316 19124 22372
rect 19068 21868 19124 21924
rect 18844 20972 18900 21028
rect 19068 21196 19124 21252
rect 18732 19964 18788 20020
rect 18620 19906 18676 19908
rect 18620 19854 18622 19906
rect 18622 19854 18674 19906
rect 18674 19854 18676 19906
rect 18620 19852 18676 19854
rect 18508 18956 18564 19012
rect 18620 19516 18676 19572
rect 18508 17612 18564 17668
rect 18508 17106 18564 17108
rect 18508 17054 18510 17106
rect 18510 17054 18562 17106
rect 18562 17054 18564 17106
rect 18508 17052 18564 17054
rect 18844 19628 18900 19684
rect 19292 22092 19348 22148
rect 19292 21586 19348 21588
rect 19292 21534 19294 21586
rect 19294 21534 19346 21586
rect 19346 21534 19348 21586
rect 19292 21532 19348 21534
rect 19292 21084 19348 21140
rect 19740 25394 19796 25396
rect 19740 25342 19742 25394
rect 19742 25342 19794 25394
rect 19794 25342 19796 25394
rect 19740 25340 19796 25342
rect 20972 31778 21028 31780
rect 20972 31726 20974 31778
rect 20974 31726 21026 31778
rect 21026 31726 21028 31778
rect 20972 31724 21028 31726
rect 20972 31052 21028 31108
rect 21308 34076 21364 34132
rect 22428 55298 22484 55300
rect 22428 55246 22430 55298
rect 22430 55246 22482 55298
rect 22482 55246 22484 55298
rect 22428 55244 22484 55246
rect 24332 56588 24388 56644
rect 23804 56474 23860 56476
rect 23804 56422 23806 56474
rect 23806 56422 23858 56474
rect 23858 56422 23860 56474
rect 23804 56420 23860 56422
rect 23908 56474 23964 56476
rect 23908 56422 23910 56474
rect 23910 56422 23962 56474
rect 23962 56422 23964 56474
rect 23908 56420 23964 56422
rect 24012 56474 24068 56476
rect 24012 56422 24014 56474
rect 24014 56422 24066 56474
rect 24066 56422 24068 56474
rect 24012 56420 24068 56422
rect 23548 56252 23604 56308
rect 23548 55356 23604 55412
rect 21980 54012 22036 54068
rect 22764 53730 22820 53732
rect 22764 53678 22766 53730
rect 22766 53678 22818 53730
rect 22818 53678 22820 53730
rect 22764 53676 22820 53678
rect 24220 55916 24276 55972
rect 23804 54906 23860 54908
rect 23804 54854 23806 54906
rect 23806 54854 23858 54906
rect 23858 54854 23860 54906
rect 23804 54852 23860 54854
rect 23908 54906 23964 54908
rect 23908 54854 23910 54906
rect 23910 54854 23962 54906
rect 23962 54854 23964 54906
rect 23908 54852 23964 54854
rect 24012 54906 24068 54908
rect 24012 54854 24014 54906
rect 24014 54854 24066 54906
rect 24066 54854 24068 54906
rect 24012 54852 24068 54854
rect 23772 54738 23828 54740
rect 23772 54686 23774 54738
rect 23774 54686 23826 54738
rect 23826 54686 23828 54738
rect 23772 54684 23828 54686
rect 24108 54514 24164 54516
rect 24108 54462 24110 54514
rect 24110 54462 24162 54514
rect 24162 54462 24164 54514
rect 24108 54460 24164 54462
rect 23660 54012 23716 54068
rect 23804 53338 23860 53340
rect 23804 53286 23806 53338
rect 23806 53286 23858 53338
rect 23858 53286 23860 53338
rect 23804 53284 23860 53286
rect 23908 53338 23964 53340
rect 23908 53286 23910 53338
rect 23910 53286 23962 53338
rect 23962 53286 23964 53338
rect 23908 53284 23964 53286
rect 24012 53338 24068 53340
rect 24012 53286 24014 53338
rect 24014 53286 24066 53338
rect 24066 53286 24068 53338
rect 24012 53284 24068 53286
rect 22764 52162 22820 52164
rect 22764 52110 22766 52162
rect 22766 52110 22818 52162
rect 22818 52110 22820 52162
rect 22764 52108 22820 52110
rect 22428 50764 22484 50820
rect 24444 56306 24500 56308
rect 24444 56254 24446 56306
rect 24446 56254 24498 56306
rect 24498 56254 24500 56306
rect 24444 56252 24500 56254
rect 24892 56252 24948 56308
rect 25004 57148 25060 57204
rect 24464 55690 24520 55692
rect 24464 55638 24466 55690
rect 24466 55638 24518 55690
rect 24518 55638 24520 55690
rect 24464 55636 24520 55638
rect 24568 55690 24624 55692
rect 24568 55638 24570 55690
rect 24570 55638 24622 55690
rect 24622 55638 24624 55690
rect 24568 55636 24624 55638
rect 24672 55690 24728 55692
rect 24672 55638 24674 55690
rect 24674 55638 24726 55690
rect 24726 55638 24728 55690
rect 24672 55636 24728 55638
rect 24892 55298 24948 55300
rect 24892 55246 24894 55298
rect 24894 55246 24946 55298
rect 24946 55246 24948 55298
rect 24892 55244 24948 55246
rect 24464 54122 24520 54124
rect 24464 54070 24466 54122
rect 24466 54070 24518 54122
rect 24518 54070 24520 54122
rect 24464 54068 24520 54070
rect 24568 54122 24624 54124
rect 24568 54070 24570 54122
rect 24570 54070 24622 54122
rect 24622 54070 24624 54122
rect 24568 54068 24624 54070
rect 24672 54122 24728 54124
rect 24672 54070 24674 54122
rect 24674 54070 24726 54122
rect 24726 54070 24728 54122
rect 24672 54068 24728 54070
rect 24892 53900 24948 53956
rect 24668 53564 24724 53620
rect 23660 52722 23716 52724
rect 23660 52670 23662 52722
rect 23662 52670 23714 52722
rect 23714 52670 23716 52722
rect 23660 52668 23716 52670
rect 24668 52834 24724 52836
rect 24668 52782 24670 52834
rect 24670 52782 24722 52834
rect 24722 52782 24724 52834
rect 24668 52780 24724 52782
rect 25452 55970 25508 55972
rect 25452 55918 25454 55970
rect 25454 55918 25506 55970
rect 25506 55918 25508 55970
rect 25452 55916 25508 55918
rect 25004 52668 25060 52724
rect 25340 55244 25396 55300
rect 24464 52554 24520 52556
rect 24464 52502 24466 52554
rect 24466 52502 24518 52554
rect 24518 52502 24520 52554
rect 24464 52500 24520 52502
rect 24568 52554 24624 52556
rect 24568 52502 24570 52554
rect 24570 52502 24622 52554
rect 24622 52502 24624 52554
rect 24568 52500 24624 52502
rect 24672 52554 24728 52556
rect 24672 52502 24674 52554
rect 24674 52502 24726 52554
rect 24726 52502 24728 52554
rect 24672 52500 24728 52502
rect 24892 52162 24948 52164
rect 24892 52110 24894 52162
rect 24894 52110 24946 52162
rect 24946 52110 24948 52162
rect 24892 52108 24948 52110
rect 23804 51770 23860 51772
rect 23804 51718 23806 51770
rect 23806 51718 23858 51770
rect 23858 51718 23860 51770
rect 23804 51716 23860 51718
rect 23908 51770 23964 51772
rect 23908 51718 23910 51770
rect 23910 51718 23962 51770
rect 23962 51718 23964 51770
rect 23908 51716 23964 51718
rect 24012 51770 24068 51772
rect 24012 51718 24014 51770
rect 24014 51718 24066 51770
rect 24066 51718 24068 51770
rect 24012 51716 24068 51718
rect 24668 51266 24724 51268
rect 24668 51214 24670 51266
rect 24670 51214 24722 51266
rect 24722 51214 24724 51266
rect 24668 51212 24724 51214
rect 24464 50986 24520 50988
rect 24464 50934 24466 50986
rect 24466 50934 24518 50986
rect 24518 50934 24520 50986
rect 24464 50932 24520 50934
rect 24568 50986 24624 50988
rect 24568 50934 24570 50986
rect 24570 50934 24622 50986
rect 24622 50934 24624 50986
rect 24568 50932 24624 50934
rect 24672 50986 24728 50988
rect 24672 50934 24674 50986
rect 24674 50934 24726 50986
rect 24726 50934 24728 50986
rect 24672 50932 24728 50934
rect 23884 50594 23940 50596
rect 23884 50542 23886 50594
rect 23886 50542 23938 50594
rect 23938 50542 23940 50594
rect 23884 50540 23940 50542
rect 24668 50428 24724 50484
rect 23804 50202 23860 50204
rect 23804 50150 23806 50202
rect 23806 50150 23858 50202
rect 23858 50150 23860 50202
rect 23804 50148 23860 50150
rect 23908 50202 23964 50204
rect 23908 50150 23910 50202
rect 23910 50150 23962 50202
rect 23962 50150 23964 50202
rect 23908 50148 23964 50150
rect 24012 50202 24068 50204
rect 24012 50150 24014 50202
rect 24014 50150 24066 50202
rect 24066 50150 24068 50202
rect 24012 50148 24068 50150
rect 24668 49698 24724 49700
rect 24668 49646 24670 49698
rect 24670 49646 24722 49698
rect 24722 49646 24724 49698
rect 24668 49644 24724 49646
rect 24464 49418 24520 49420
rect 24464 49366 24466 49418
rect 24466 49366 24518 49418
rect 24518 49366 24520 49418
rect 24464 49364 24520 49366
rect 24568 49418 24624 49420
rect 24568 49366 24570 49418
rect 24570 49366 24622 49418
rect 24622 49366 24624 49418
rect 24568 49364 24624 49366
rect 24672 49418 24728 49420
rect 24672 49366 24674 49418
rect 24674 49366 24726 49418
rect 24726 49366 24728 49418
rect 24672 49364 24728 49366
rect 24668 49026 24724 49028
rect 24668 48974 24670 49026
rect 24670 48974 24722 49026
rect 24722 48974 24724 49026
rect 24668 48972 24724 48974
rect 23804 48634 23860 48636
rect 23804 48582 23806 48634
rect 23806 48582 23858 48634
rect 23858 48582 23860 48634
rect 23804 48580 23860 48582
rect 23908 48634 23964 48636
rect 23908 48582 23910 48634
rect 23910 48582 23962 48634
rect 23962 48582 23964 48634
rect 23908 48580 23964 48582
rect 24012 48634 24068 48636
rect 24012 48582 24014 48634
rect 24014 48582 24066 48634
rect 24066 48582 24068 48634
rect 24012 48580 24068 48582
rect 24464 47850 24520 47852
rect 24464 47798 24466 47850
rect 24466 47798 24518 47850
rect 24518 47798 24520 47850
rect 24464 47796 24520 47798
rect 24568 47850 24624 47852
rect 24568 47798 24570 47850
rect 24570 47798 24622 47850
rect 24622 47798 24624 47850
rect 24568 47796 24624 47798
rect 24672 47850 24728 47852
rect 24672 47798 24674 47850
rect 24674 47798 24726 47850
rect 24726 47798 24728 47850
rect 24672 47796 24728 47798
rect 24668 47458 24724 47460
rect 24668 47406 24670 47458
rect 24670 47406 24722 47458
rect 24722 47406 24724 47458
rect 24668 47404 24724 47406
rect 23804 47066 23860 47068
rect 23804 47014 23806 47066
rect 23806 47014 23858 47066
rect 23858 47014 23860 47066
rect 23804 47012 23860 47014
rect 23908 47066 23964 47068
rect 23908 47014 23910 47066
rect 23910 47014 23962 47066
rect 23962 47014 23964 47066
rect 23908 47012 23964 47014
rect 24012 47066 24068 47068
rect 24012 47014 24014 47066
rect 24014 47014 24066 47066
rect 24066 47014 24068 47066
rect 24012 47012 24068 47014
rect 24668 46562 24724 46564
rect 24668 46510 24670 46562
rect 24670 46510 24722 46562
rect 24722 46510 24724 46562
rect 24668 46508 24724 46510
rect 24464 46282 24520 46284
rect 24464 46230 24466 46282
rect 24466 46230 24518 46282
rect 24518 46230 24520 46282
rect 24464 46228 24520 46230
rect 24568 46282 24624 46284
rect 24568 46230 24570 46282
rect 24570 46230 24622 46282
rect 24622 46230 24624 46282
rect 24568 46228 24624 46230
rect 24672 46282 24728 46284
rect 24672 46230 24674 46282
rect 24674 46230 24726 46282
rect 24726 46230 24728 46282
rect 24672 46228 24728 46230
rect 24668 45890 24724 45892
rect 24668 45838 24670 45890
rect 24670 45838 24722 45890
rect 24722 45838 24724 45890
rect 24668 45836 24724 45838
rect 23804 45498 23860 45500
rect 23804 45446 23806 45498
rect 23806 45446 23858 45498
rect 23858 45446 23860 45498
rect 23804 45444 23860 45446
rect 23908 45498 23964 45500
rect 23908 45446 23910 45498
rect 23910 45446 23962 45498
rect 23962 45446 23964 45498
rect 23908 45444 23964 45446
rect 24012 45498 24068 45500
rect 24012 45446 24014 45498
rect 24014 45446 24066 45498
rect 24066 45446 24068 45498
rect 24012 45444 24068 45446
rect 24464 44714 24520 44716
rect 24464 44662 24466 44714
rect 24466 44662 24518 44714
rect 24518 44662 24520 44714
rect 24464 44660 24520 44662
rect 24568 44714 24624 44716
rect 24568 44662 24570 44714
rect 24570 44662 24622 44714
rect 24622 44662 24624 44714
rect 24568 44660 24624 44662
rect 24672 44714 24728 44716
rect 24672 44662 24674 44714
rect 24674 44662 24726 44714
rect 24726 44662 24728 44714
rect 24672 44660 24728 44662
rect 24668 44322 24724 44324
rect 24668 44270 24670 44322
rect 24670 44270 24722 44322
rect 24722 44270 24724 44322
rect 24668 44268 24724 44270
rect 23804 43930 23860 43932
rect 23804 43878 23806 43930
rect 23806 43878 23858 43930
rect 23858 43878 23860 43930
rect 23804 43876 23860 43878
rect 23908 43930 23964 43932
rect 23908 43878 23910 43930
rect 23910 43878 23962 43930
rect 23962 43878 23964 43930
rect 23908 43876 23964 43878
rect 24012 43930 24068 43932
rect 24012 43878 24014 43930
rect 24014 43878 24066 43930
rect 24066 43878 24068 43930
rect 24012 43876 24068 43878
rect 23324 42812 23380 42868
rect 22316 39564 22372 39620
rect 21532 33068 21588 33124
rect 21868 34524 21924 34580
rect 21420 31948 21476 32004
rect 21532 31724 21588 31780
rect 20524 25900 20580 25956
rect 20188 25228 20244 25284
rect 20524 25340 20580 25396
rect 19628 22370 19684 22372
rect 19628 22318 19630 22370
rect 19630 22318 19682 22370
rect 19682 22318 19684 22370
rect 19628 22316 19684 22318
rect 20748 25340 20804 25396
rect 20188 23436 20244 23492
rect 21308 31500 21364 31556
rect 21420 30210 21476 30212
rect 21420 30158 21422 30210
rect 21422 30158 21474 30210
rect 21474 30158 21476 30210
rect 21420 30156 21476 30158
rect 21308 27132 21364 27188
rect 21084 25900 21140 25956
rect 21308 26066 21364 26068
rect 21308 26014 21310 26066
rect 21310 26014 21362 26066
rect 21362 26014 21364 26066
rect 21308 26012 21364 26014
rect 21644 30268 21700 30324
rect 21756 30156 21812 30212
rect 22092 32674 22148 32676
rect 22092 32622 22094 32674
rect 22094 32622 22146 32674
rect 22146 32622 22148 32674
rect 22092 32620 22148 32622
rect 22092 30994 22148 30996
rect 22092 30942 22094 30994
rect 22094 30942 22146 30994
rect 22146 30942 22148 30994
rect 22092 30940 22148 30942
rect 21532 27468 21588 27524
rect 21532 27132 21588 27188
rect 21308 25340 21364 25396
rect 21420 25228 21476 25284
rect 21084 24108 21140 24164
rect 20972 24050 21028 24052
rect 20972 23998 20974 24050
rect 20974 23998 21026 24050
rect 21026 23998 21028 24050
rect 20972 23996 21028 23998
rect 20076 23100 20132 23156
rect 19740 21980 19796 22036
rect 19852 22092 19908 22148
rect 19516 21532 19572 21588
rect 20076 22204 20132 22260
rect 20188 22316 20244 22372
rect 19628 21362 19684 21364
rect 19628 21310 19630 21362
rect 19630 21310 19682 21362
rect 19682 21310 19684 21362
rect 19628 21308 19684 21310
rect 19404 20972 19460 21028
rect 19516 21084 19572 21140
rect 19964 21084 20020 21140
rect 20076 20972 20132 21028
rect 19404 20188 19460 20244
rect 19740 20188 19796 20244
rect 19964 20188 20020 20244
rect 20636 21308 20692 21364
rect 20748 21196 20804 21252
rect 20188 20076 20244 20132
rect 19740 19852 19796 19908
rect 19852 19964 19908 20020
rect 19516 19628 19572 19684
rect 19180 18956 19236 19012
rect 18844 18844 18900 18900
rect 19292 18844 19348 18900
rect 18844 18172 18900 18228
rect 19068 18060 19124 18116
rect 19292 18172 19348 18228
rect 18844 17778 18900 17780
rect 18844 17726 18846 17778
rect 18846 17726 18898 17778
rect 18898 17726 18900 17778
rect 18844 17724 18900 17726
rect 19292 17666 19348 17668
rect 19292 17614 19294 17666
rect 19294 17614 19346 17666
rect 19346 17614 19348 17666
rect 19292 17612 19348 17614
rect 20412 19516 20468 19572
rect 19852 19180 19908 19236
rect 21084 21586 21140 21588
rect 21084 21534 21086 21586
rect 21086 21534 21138 21586
rect 21138 21534 21140 21586
rect 21084 21532 21140 21534
rect 20972 20412 21028 20468
rect 20860 20188 20916 20244
rect 20972 20130 21028 20132
rect 20972 20078 20974 20130
rect 20974 20078 21026 20130
rect 21026 20078 21028 20130
rect 20972 20076 21028 20078
rect 20860 19906 20916 19908
rect 20860 19854 20862 19906
rect 20862 19854 20914 19906
rect 20914 19854 20916 19906
rect 20860 19852 20916 19854
rect 21196 21308 21252 21364
rect 23212 31388 23268 31444
rect 22428 30716 22484 30772
rect 22092 26908 22148 26964
rect 21868 26012 21924 26068
rect 21756 25228 21812 25284
rect 21084 19852 21140 19908
rect 21196 20412 21252 20468
rect 20076 18844 20132 18900
rect 19516 17836 19572 17892
rect 19404 17164 19460 17220
rect 18732 17052 18788 17108
rect 18172 15820 18228 15876
rect 18620 16604 18676 16660
rect 18732 16492 18788 16548
rect 18956 16380 19012 16436
rect 18732 16044 18788 16100
rect 18508 15708 18564 15764
rect 18396 15314 18452 15316
rect 18396 15262 18398 15314
rect 18398 15262 18450 15314
rect 18450 15262 18452 15314
rect 18396 15260 18452 15262
rect 17948 14252 18004 14308
rect 18060 14530 18116 14532
rect 18060 14478 18062 14530
rect 18062 14478 18114 14530
rect 18114 14478 18116 14530
rect 18060 14476 18116 14478
rect 17836 13074 17892 13076
rect 17836 13022 17838 13074
rect 17838 13022 17890 13074
rect 17890 13022 17892 13074
rect 17836 13020 17892 13022
rect 18060 12796 18116 12852
rect 17724 12684 17780 12740
rect 17612 12236 17668 12292
rect 17836 11788 17892 11844
rect 18060 11788 18116 11844
rect 16828 10220 16884 10276
rect 16940 9884 16996 9940
rect 17276 9996 17332 10052
rect 17052 9826 17108 9828
rect 17052 9774 17054 9826
rect 17054 9774 17106 9826
rect 17106 9774 17108 9826
rect 17052 9772 17108 9774
rect 17276 9826 17332 9828
rect 17276 9774 17278 9826
rect 17278 9774 17330 9826
rect 17330 9774 17332 9826
rect 17276 9772 17332 9774
rect 16940 8258 16996 8260
rect 16940 8206 16942 8258
rect 16942 8206 16994 8258
rect 16994 8206 16996 8258
rect 16940 8204 16996 8206
rect 16156 8034 16212 8036
rect 16156 7982 16158 8034
rect 16158 7982 16210 8034
rect 16210 7982 16212 8034
rect 16156 7980 16212 7982
rect 16156 7474 16212 7476
rect 16156 7422 16158 7474
rect 16158 7422 16210 7474
rect 16210 7422 16212 7474
rect 16156 7420 16212 7422
rect 16380 7308 16436 7364
rect 17724 10722 17780 10724
rect 17724 10670 17726 10722
rect 17726 10670 17778 10722
rect 17778 10670 17780 10722
rect 17724 10668 17780 10670
rect 17612 9884 17668 9940
rect 17724 10220 17780 10276
rect 17836 9996 17892 10052
rect 18060 10108 18116 10164
rect 17724 9772 17780 9828
rect 17612 9324 17668 9380
rect 17836 9436 17892 9492
rect 17836 8428 17892 8484
rect 16716 8034 16772 8036
rect 16716 7982 16718 8034
rect 16718 7982 16770 8034
rect 16770 7982 16772 8034
rect 16716 7980 16772 7982
rect 16604 7756 16660 7812
rect 17052 7756 17108 7812
rect 16716 7698 16772 7700
rect 16716 7646 16718 7698
rect 16718 7646 16770 7698
rect 16770 7646 16772 7698
rect 16716 7644 16772 7646
rect 17388 7644 17444 7700
rect 16492 6524 16548 6580
rect 16940 7420 16996 7476
rect 17388 7474 17444 7476
rect 17388 7422 17390 7474
rect 17390 7422 17442 7474
rect 17442 7422 17444 7474
rect 17388 7420 17444 7422
rect 15932 5292 15988 5348
rect 15708 5068 15764 5124
rect 15484 4844 15540 4900
rect 10108 924 10164 980
rect 13244 2098 13300 2100
rect 13244 2046 13246 2098
rect 13246 2046 13298 2098
rect 13298 2046 13300 2098
rect 13244 2044 13300 2046
rect 11900 924 11956 980
rect 13804 1986 13860 1988
rect 13804 1934 13806 1986
rect 13806 1934 13858 1986
rect 13858 1934 13860 1986
rect 13804 1932 13860 1934
rect 12012 588 12068 644
rect 12796 1260 12852 1316
rect 14140 924 14196 980
rect 18396 15090 18452 15092
rect 18396 15038 18398 15090
rect 18398 15038 18450 15090
rect 18450 15038 18452 15090
rect 18396 15036 18452 15038
rect 18844 15820 18900 15876
rect 18620 14588 18676 14644
rect 18396 14252 18452 14308
rect 18284 13020 18340 13076
rect 19404 16380 19460 16436
rect 19740 16828 19796 16884
rect 19964 17836 20020 17892
rect 20860 18620 20916 18676
rect 20524 18172 20580 18228
rect 19628 16044 19684 16100
rect 19740 16380 19796 16436
rect 19180 15932 19236 15988
rect 19740 15314 19796 15316
rect 19740 15262 19742 15314
rect 19742 15262 19794 15314
rect 19794 15262 19796 15314
rect 19740 15260 19796 15262
rect 19180 14476 19236 14532
rect 19292 14588 19348 14644
rect 19740 14588 19796 14644
rect 19068 14028 19124 14084
rect 19292 13970 19348 13972
rect 19292 13918 19294 13970
rect 19294 13918 19346 13970
rect 19346 13918 19348 13970
rect 19292 13916 19348 13918
rect 19740 13858 19796 13860
rect 19740 13806 19742 13858
rect 19742 13806 19794 13858
rect 19794 13806 19796 13858
rect 19740 13804 19796 13806
rect 19740 13522 19796 13524
rect 19740 13470 19742 13522
rect 19742 13470 19794 13522
rect 19794 13470 19796 13522
rect 19740 13468 19796 13470
rect 19516 13244 19572 13300
rect 19180 13074 19236 13076
rect 19180 13022 19182 13074
rect 19182 13022 19234 13074
rect 19234 13022 19236 13074
rect 19180 13020 19236 13022
rect 18396 12962 18452 12964
rect 18396 12910 18398 12962
rect 18398 12910 18450 12962
rect 18450 12910 18452 12962
rect 18396 12908 18452 12910
rect 19628 12796 19684 12852
rect 19628 12236 19684 12292
rect 18508 12178 18564 12180
rect 18508 12126 18510 12178
rect 18510 12126 18562 12178
rect 18562 12126 18564 12178
rect 18508 12124 18564 12126
rect 18396 11452 18452 11508
rect 18284 10834 18340 10836
rect 18284 10782 18286 10834
rect 18286 10782 18338 10834
rect 18338 10782 18340 10834
rect 18284 10780 18340 10782
rect 18508 11394 18564 11396
rect 18508 11342 18510 11394
rect 18510 11342 18562 11394
rect 18562 11342 18564 11394
rect 18508 11340 18564 11342
rect 18508 11004 18564 11060
rect 17948 5180 18004 5236
rect 17500 4172 17556 4228
rect 18844 11954 18900 11956
rect 18844 11902 18846 11954
rect 18846 11902 18898 11954
rect 18898 11902 18900 11954
rect 18844 11900 18900 11902
rect 19516 11900 19572 11956
rect 19292 11788 19348 11844
rect 19180 11506 19236 11508
rect 19180 11454 19182 11506
rect 19182 11454 19234 11506
rect 19234 11454 19236 11506
rect 19180 11452 19236 11454
rect 18620 10668 18676 10724
rect 18956 10050 19012 10052
rect 18956 9998 18958 10050
rect 18958 9998 19010 10050
rect 19010 9998 19012 10050
rect 18956 9996 19012 9998
rect 19404 11116 19460 11172
rect 19292 9884 19348 9940
rect 19404 10108 19460 10164
rect 18172 8988 18228 9044
rect 18844 8316 18900 8372
rect 20076 15372 20132 15428
rect 20300 18060 20356 18116
rect 20076 15202 20132 15204
rect 20076 15150 20078 15202
rect 20078 15150 20130 15202
rect 20130 15150 20132 15202
rect 20076 15148 20132 15150
rect 19964 13916 20020 13972
rect 20076 14252 20132 14308
rect 19964 13634 20020 13636
rect 19964 13582 19966 13634
rect 19966 13582 20018 13634
rect 20018 13582 20020 13634
rect 19964 13580 20020 13582
rect 19740 11900 19796 11956
rect 19852 12908 19908 12964
rect 20076 12796 20132 12852
rect 19964 12178 20020 12180
rect 19964 12126 19966 12178
rect 19966 12126 20018 12178
rect 20018 12126 20020 12178
rect 19964 12124 20020 12126
rect 20188 11788 20244 11844
rect 20076 11340 20132 11396
rect 19964 10780 20020 10836
rect 19852 10610 19908 10612
rect 19852 10558 19854 10610
rect 19854 10558 19906 10610
rect 19906 10558 19908 10610
rect 19852 10556 19908 10558
rect 19516 8428 19572 8484
rect 20076 8204 20132 8260
rect 19068 7980 19124 8036
rect 18060 2716 18116 2772
rect 18508 6524 18564 6580
rect 20412 16156 20468 16212
rect 20636 17612 20692 17668
rect 20972 18172 21028 18228
rect 20972 17276 21028 17332
rect 20972 16882 21028 16884
rect 20972 16830 20974 16882
rect 20974 16830 21026 16882
rect 21026 16830 21028 16882
rect 20972 16828 21028 16830
rect 20636 16492 20692 16548
rect 20636 15596 20692 15652
rect 20860 16658 20916 16660
rect 20860 16606 20862 16658
rect 20862 16606 20914 16658
rect 20914 16606 20916 16658
rect 20860 16604 20916 16606
rect 20636 15426 20692 15428
rect 20636 15374 20638 15426
rect 20638 15374 20690 15426
rect 20690 15374 20692 15426
rect 20636 15372 20692 15374
rect 20524 15260 20580 15316
rect 20524 14924 20580 14980
rect 20748 14530 20804 14532
rect 20748 14478 20750 14530
rect 20750 14478 20802 14530
rect 20802 14478 20804 14530
rect 20748 14476 20804 14478
rect 21308 20300 21364 20356
rect 21420 22204 21476 22260
rect 21308 19964 21364 20020
rect 22092 24162 22148 24164
rect 22092 24110 22094 24162
rect 22094 24110 22146 24162
rect 22146 24110 22148 24162
rect 22092 24108 22148 24110
rect 21868 22428 21924 22484
rect 22316 26908 22372 26964
rect 23100 30210 23156 30212
rect 23100 30158 23102 30210
rect 23102 30158 23154 30210
rect 23154 30158 23156 30210
rect 23100 30156 23156 30158
rect 22988 28924 23044 28980
rect 22540 24050 22596 24052
rect 22540 23998 22542 24050
rect 22542 23998 22594 24050
rect 22594 23998 22596 24050
rect 22540 23996 22596 23998
rect 21980 21756 22036 21812
rect 21756 20802 21812 20804
rect 21756 20750 21758 20802
rect 21758 20750 21810 20802
rect 21810 20750 21812 20802
rect 21756 20748 21812 20750
rect 21644 20300 21700 20356
rect 21644 18396 21700 18452
rect 21420 18060 21476 18116
rect 21532 18172 21588 18228
rect 21644 17948 21700 18004
rect 21308 16492 21364 16548
rect 21532 17612 21588 17668
rect 21084 15036 21140 15092
rect 21196 15260 21252 15316
rect 21196 14924 21252 14980
rect 21084 14476 21140 14532
rect 20972 14252 21028 14308
rect 21420 15932 21476 15988
rect 21420 15708 21476 15764
rect 21420 14306 21476 14308
rect 21420 14254 21422 14306
rect 21422 14254 21474 14306
rect 21474 14254 21476 14306
rect 21420 14252 21476 14254
rect 20860 13692 20916 13748
rect 20524 13356 20580 13412
rect 20300 8316 20356 8372
rect 20412 12796 20468 12852
rect 20524 12460 20580 12516
rect 21420 13746 21476 13748
rect 21420 13694 21422 13746
rect 21422 13694 21474 13746
rect 21474 13694 21476 13746
rect 21420 13692 21476 13694
rect 20972 13580 21028 13636
rect 20748 13522 20804 13524
rect 20748 13470 20750 13522
rect 20750 13470 20802 13522
rect 20802 13470 20804 13522
rect 20748 13468 20804 13470
rect 20860 13356 20916 13412
rect 21644 15148 21700 15204
rect 21084 13244 21140 13300
rect 21644 13692 21700 13748
rect 20860 12460 20916 12516
rect 21084 11954 21140 11956
rect 21084 11902 21086 11954
rect 21086 11902 21138 11954
rect 21138 11902 21140 11954
rect 21084 11900 21140 11902
rect 20636 11788 20692 11844
rect 20860 11452 20916 11508
rect 20860 10220 20916 10276
rect 21084 9826 21140 9828
rect 21084 9774 21086 9826
rect 21086 9774 21138 9826
rect 21138 9774 21140 9826
rect 21084 9772 21140 9774
rect 20860 8988 20916 9044
rect 21420 13244 21476 13300
rect 21420 12962 21476 12964
rect 21420 12910 21422 12962
rect 21422 12910 21474 12962
rect 21474 12910 21476 12962
rect 21420 12908 21476 12910
rect 21532 12460 21588 12516
rect 21308 8204 21364 8260
rect 21420 11900 21476 11956
rect 20300 7644 20356 7700
rect 20076 7196 20132 7252
rect 19068 5404 19124 5460
rect 18508 2044 18564 2100
rect 16828 1596 16884 1652
rect 20860 1596 20916 1652
rect 18172 1260 18228 1316
rect 19516 140 19572 196
rect 21644 8258 21700 8260
rect 21644 8206 21646 8258
rect 21646 8206 21698 8258
rect 21698 8206 21700 8258
rect 21644 8204 21700 8206
rect 21644 6748 21700 6804
rect 21980 21196 22036 21252
rect 22092 20748 22148 20804
rect 22204 20076 22260 20132
rect 21980 18284 22036 18340
rect 21980 17500 22036 17556
rect 22092 17388 22148 17444
rect 22092 15314 22148 15316
rect 22092 15262 22094 15314
rect 22094 15262 22146 15314
rect 22146 15262 22148 15314
rect 22092 15260 22148 15262
rect 21868 14252 21924 14308
rect 21868 11676 21924 11732
rect 21868 9996 21924 10052
rect 21868 8092 21924 8148
rect 22204 14140 22260 14196
rect 22204 11452 22260 11508
rect 21980 3500 22036 3556
rect 21644 1820 21700 1876
rect 22204 1932 22260 1988
rect 21420 924 21476 980
rect 22652 21196 22708 21252
rect 22764 19964 22820 20020
rect 22876 22428 22932 22484
rect 22540 18396 22596 18452
rect 22652 18284 22708 18340
rect 22876 18396 22932 18452
rect 22652 17612 22708 17668
rect 22540 16268 22596 16324
rect 22540 13132 22596 13188
rect 22764 14588 22820 14644
rect 22764 13804 22820 13860
rect 22652 11788 22708 11844
rect 23100 24556 23156 24612
rect 24464 43146 24520 43148
rect 24464 43094 24466 43146
rect 24466 43094 24518 43146
rect 24518 43094 24520 43146
rect 24464 43092 24520 43094
rect 24568 43146 24624 43148
rect 24568 43094 24570 43146
rect 24570 43094 24622 43146
rect 24622 43094 24624 43146
rect 24568 43092 24624 43094
rect 24672 43146 24728 43148
rect 24672 43094 24674 43146
rect 24674 43094 24726 43146
rect 24726 43094 24728 43146
rect 24672 43092 24728 43094
rect 24668 42588 24724 42644
rect 23804 42362 23860 42364
rect 23804 42310 23806 42362
rect 23806 42310 23858 42362
rect 23858 42310 23860 42362
rect 23804 42308 23860 42310
rect 23908 42362 23964 42364
rect 23908 42310 23910 42362
rect 23910 42310 23962 42362
rect 23962 42310 23964 42362
rect 23908 42308 23964 42310
rect 24012 42362 24068 42364
rect 24012 42310 24014 42362
rect 24014 42310 24066 42362
rect 24066 42310 24068 42362
rect 24012 42308 24068 42310
rect 24464 41578 24520 41580
rect 24464 41526 24466 41578
rect 24466 41526 24518 41578
rect 24518 41526 24520 41578
rect 24464 41524 24520 41526
rect 24568 41578 24624 41580
rect 24568 41526 24570 41578
rect 24570 41526 24622 41578
rect 24622 41526 24624 41578
rect 24568 41524 24624 41526
rect 24672 41578 24728 41580
rect 24672 41526 24674 41578
rect 24674 41526 24726 41578
rect 24726 41526 24728 41578
rect 24672 41524 24728 41526
rect 23804 40794 23860 40796
rect 23804 40742 23806 40794
rect 23806 40742 23858 40794
rect 23858 40742 23860 40794
rect 23804 40740 23860 40742
rect 23908 40794 23964 40796
rect 23908 40742 23910 40794
rect 23910 40742 23962 40794
rect 23962 40742 23964 40794
rect 23908 40740 23964 40742
rect 24012 40794 24068 40796
rect 24012 40742 24014 40794
rect 24014 40742 24066 40794
rect 24066 40742 24068 40794
rect 24012 40740 24068 40742
rect 23804 39226 23860 39228
rect 23804 39174 23806 39226
rect 23806 39174 23858 39226
rect 23858 39174 23860 39226
rect 23804 39172 23860 39174
rect 23908 39226 23964 39228
rect 23908 39174 23910 39226
rect 23910 39174 23962 39226
rect 23962 39174 23964 39226
rect 23908 39172 23964 39174
rect 24012 39226 24068 39228
rect 24012 39174 24014 39226
rect 24014 39174 24066 39226
rect 24066 39174 24068 39226
rect 24012 39172 24068 39174
rect 23660 37884 23716 37940
rect 23804 37658 23860 37660
rect 23804 37606 23806 37658
rect 23806 37606 23858 37658
rect 23858 37606 23860 37658
rect 23804 37604 23860 37606
rect 23908 37658 23964 37660
rect 23908 37606 23910 37658
rect 23910 37606 23962 37658
rect 23962 37606 23964 37658
rect 23908 37604 23964 37606
rect 24012 37658 24068 37660
rect 24012 37606 24014 37658
rect 24014 37606 24066 37658
rect 24066 37606 24068 37658
rect 24012 37604 24068 37606
rect 23804 36090 23860 36092
rect 23804 36038 23806 36090
rect 23806 36038 23858 36090
rect 23858 36038 23860 36090
rect 23804 36036 23860 36038
rect 23908 36090 23964 36092
rect 23908 36038 23910 36090
rect 23910 36038 23962 36090
rect 23962 36038 23964 36090
rect 23908 36036 23964 36038
rect 24012 36090 24068 36092
rect 24012 36038 24014 36090
rect 24014 36038 24066 36090
rect 24066 36038 24068 36090
rect 24012 36036 24068 36038
rect 23804 34522 23860 34524
rect 23804 34470 23806 34522
rect 23806 34470 23858 34522
rect 23858 34470 23860 34522
rect 23804 34468 23860 34470
rect 23908 34522 23964 34524
rect 23908 34470 23910 34522
rect 23910 34470 23962 34522
rect 23962 34470 23964 34522
rect 23908 34468 23964 34470
rect 24012 34522 24068 34524
rect 24012 34470 24014 34522
rect 24014 34470 24066 34522
rect 24066 34470 24068 34522
rect 24012 34468 24068 34470
rect 23804 32954 23860 32956
rect 23804 32902 23806 32954
rect 23806 32902 23858 32954
rect 23858 32902 23860 32954
rect 23804 32900 23860 32902
rect 23908 32954 23964 32956
rect 23908 32902 23910 32954
rect 23910 32902 23962 32954
rect 23962 32902 23964 32954
rect 23908 32900 23964 32902
rect 24012 32954 24068 32956
rect 24012 32902 24014 32954
rect 24014 32902 24066 32954
rect 24066 32902 24068 32954
rect 24012 32900 24068 32902
rect 24780 40124 24836 40180
rect 24464 40010 24520 40012
rect 24332 39900 24388 39956
rect 24464 39958 24466 40010
rect 24466 39958 24518 40010
rect 24518 39958 24520 40010
rect 24464 39956 24520 39958
rect 24568 40010 24624 40012
rect 24568 39958 24570 40010
rect 24570 39958 24622 40010
rect 24622 39958 24624 40010
rect 24568 39956 24624 39958
rect 24672 40010 24728 40012
rect 24672 39958 24674 40010
rect 24674 39958 24726 40010
rect 24726 39958 24728 40010
rect 24672 39956 24728 39958
rect 24668 39618 24724 39620
rect 24668 39566 24670 39618
rect 24670 39566 24722 39618
rect 24722 39566 24724 39618
rect 24668 39564 24724 39566
rect 24464 38442 24520 38444
rect 24464 38390 24466 38442
rect 24466 38390 24518 38442
rect 24518 38390 24520 38442
rect 24464 38388 24520 38390
rect 24568 38442 24624 38444
rect 24568 38390 24570 38442
rect 24570 38390 24622 38442
rect 24622 38390 24624 38442
rect 24568 38388 24624 38390
rect 24672 38442 24728 38444
rect 24672 38390 24674 38442
rect 24674 38390 24726 38442
rect 24726 38390 24728 38442
rect 24672 38388 24728 38390
rect 24892 38220 24948 38276
rect 24668 37154 24724 37156
rect 24668 37102 24670 37154
rect 24670 37102 24722 37154
rect 24722 37102 24724 37154
rect 24668 37100 24724 37102
rect 24464 36874 24520 36876
rect 24464 36822 24466 36874
rect 24466 36822 24518 36874
rect 24518 36822 24520 36874
rect 24464 36820 24520 36822
rect 24568 36874 24624 36876
rect 24568 36822 24570 36874
rect 24570 36822 24622 36874
rect 24622 36822 24624 36874
rect 24568 36820 24624 36822
rect 24672 36874 24728 36876
rect 24672 36822 24674 36874
rect 24674 36822 24726 36874
rect 24726 36822 24728 36874
rect 24672 36820 24728 36822
rect 24892 36204 24948 36260
rect 24464 35306 24520 35308
rect 24464 35254 24466 35306
rect 24466 35254 24518 35306
rect 24518 35254 24520 35306
rect 24464 35252 24520 35254
rect 24568 35306 24624 35308
rect 24568 35254 24570 35306
rect 24570 35254 24622 35306
rect 24622 35254 24624 35306
rect 24568 35252 24624 35254
rect 24672 35306 24728 35308
rect 24672 35254 24674 35306
rect 24674 35254 24726 35306
rect 24726 35254 24728 35306
rect 24672 35252 24728 35254
rect 24668 33852 24724 33908
rect 24464 33738 24520 33740
rect 24464 33686 24466 33738
rect 24466 33686 24518 33738
rect 24518 33686 24520 33738
rect 24464 33684 24520 33686
rect 24568 33738 24624 33740
rect 24568 33686 24570 33738
rect 24570 33686 24622 33738
rect 24622 33686 24624 33738
rect 24568 33684 24624 33686
rect 24672 33738 24728 33740
rect 24672 33686 24674 33738
rect 24674 33686 24726 33738
rect 24726 33686 24728 33738
rect 24672 33684 24728 33686
rect 24464 32170 24520 32172
rect 24464 32118 24466 32170
rect 24466 32118 24518 32170
rect 24518 32118 24520 32170
rect 24464 32116 24520 32118
rect 24568 32170 24624 32172
rect 24568 32118 24570 32170
rect 24570 32118 24622 32170
rect 24622 32118 24624 32170
rect 24568 32116 24624 32118
rect 24672 32170 24728 32172
rect 24672 32118 24674 32170
rect 24674 32118 24726 32170
rect 24726 32118 24728 32170
rect 24672 32116 24728 32118
rect 24220 31948 24276 32004
rect 24780 31836 24836 31892
rect 23660 31388 23716 31444
rect 23804 31386 23860 31388
rect 23804 31334 23806 31386
rect 23806 31334 23858 31386
rect 23858 31334 23860 31386
rect 23804 31332 23860 31334
rect 23908 31386 23964 31388
rect 23908 31334 23910 31386
rect 23910 31334 23962 31386
rect 23962 31334 23964 31386
rect 23908 31332 23964 31334
rect 24012 31386 24068 31388
rect 24012 31334 24014 31386
rect 24014 31334 24066 31386
rect 24066 31334 24068 31386
rect 24012 31332 24068 31334
rect 23660 30994 23716 30996
rect 23660 30942 23662 30994
rect 23662 30942 23714 30994
rect 23714 30942 23716 30994
rect 23660 30940 23716 30942
rect 24892 31164 24948 31220
rect 24464 30602 24520 30604
rect 24464 30550 24466 30602
rect 24466 30550 24518 30602
rect 24518 30550 24520 30602
rect 24464 30548 24520 30550
rect 24568 30602 24624 30604
rect 24568 30550 24570 30602
rect 24570 30550 24622 30602
rect 24622 30550 24624 30602
rect 24568 30548 24624 30550
rect 24672 30602 24728 30604
rect 24672 30550 24674 30602
rect 24674 30550 24726 30602
rect 24726 30550 24728 30602
rect 24672 30548 24728 30550
rect 23804 29818 23860 29820
rect 23804 29766 23806 29818
rect 23806 29766 23858 29818
rect 23858 29766 23860 29818
rect 23804 29764 23860 29766
rect 23908 29818 23964 29820
rect 23908 29766 23910 29818
rect 23910 29766 23962 29818
rect 23962 29766 23964 29818
rect 23908 29764 23964 29766
rect 24012 29818 24068 29820
rect 24012 29766 24014 29818
rect 24014 29766 24066 29818
rect 24066 29766 24068 29818
rect 24012 29764 24068 29766
rect 24464 29034 24520 29036
rect 24464 28982 24466 29034
rect 24466 28982 24518 29034
rect 24518 28982 24520 29034
rect 24464 28980 24520 28982
rect 24568 29034 24624 29036
rect 24568 28982 24570 29034
rect 24570 28982 24622 29034
rect 24622 28982 24624 29034
rect 24568 28980 24624 28982
rect 24672 29034 24728 29036
rect 24672 28982 24674 29034
rect 24674 28982 24726 29034
rect 24726 28982 24728 29034
rect 24672 28980 24728 28982
rect 23804 28250 23860 28252
rect 23804 28198 23806 28250
rect 23806 28198 23858 28250
rect 23858 28198 23860 28250
rect 23804 28196 23860 28198
rect 23908 28250 23964 28252
rect 23908 28198 23910 28250
rect 23910 28198 23962 28250
rect 23962 28198 23964 28250
rect 23908 28196 23964 28198
rect 24012 28250 24068 28252
rect 24012 28198 24014 28250
rect 24014 28198 24066 28250
rect 24066 28198 24068 28250
rect 24012 28196 24068 28198
rect 25004 28028 25060 28084
rect 24464 27466 24520 27468
rect 24464 27414 24466 27466
rect 24466 27414 24518 27466
rect 24518 27414 24520 27466
rect 24464 27412 24520 27414
rect 24568 27466 24624 27468
rect 24568 27414 24570 27466
rect 24570 27414 24622 27466
rect 24622 27414 24624 27466
rect 24568 27412 24624 27414
rect 24672 27466 24728 27468
rect 24672 27414 24674 27466
rect 24674 27414 24726 27466
rect 24726 27414 24728 27466
rect 24672 27412 24728 27414
rect 24892 27244 24948 27300
rect 23804 26682 23860 26684
rect 23804 26630 23806 26682
rect 23806 26630 23858 26682
rect 23858 26630 23860 26682
rect 23804 26628 23860 26630
rect 23908 26682 23964 26684
rect 23908 26630 23910 26682
rect 23910 26630 23962 26682
rect 23962 26630 23964 26682
rect 23908 26628 23964 26630
rect 24012 26682 24068 26684
rect 24012 26630 24014 26682
rect 24014 26630 24066 26682
rect 24066 26630 24068 26682
rect 24012 26628 24068 26630
rect 23804 25114 23860 25116
rect 23804 25062 23806 25114
rect 23806 25062 23858 25114
rect 23858 25062 23860 25114
rect 23804 25060 23860 25062
rect 23908 25114 23964 25116
rect 23908 25062 23910 25114
rect 23910 25062 23962 25114
rect 23962 25062 23964 25114
rect 23908 25060 23964 25062
rect 24012 25114 24068 25116
rect 24012 25062 24014 25114
rect 24014 25062 24066 25114
rect 24066 25062 24068 25114
rect 24012 25060 24068 25062
rect 23436 22876 23492 22932
rect 23548 23436 23604 23492
rect 23436 22482 23492 22484
rect 23436 22430 23438 22482
rect 23438 22430 23490 22482
rect 23490 22430 23492 22482
rect 23436 22428 23492 22430
rect 23548 22092 23604 22148
rect 23804 23546 23860 23548
rect 23804 23494 23806 23546
rect 23806 23494 23858 23546
rect 23858 23494 23860 23546
rect 23804 23492 23860 23494
rect 23908 23546 23964 23548
rect 23908 23494 23910 23546
rect 23910 23494 23962 23546
rect 23962 23494 23964 23546
rect 23908 23492 23964 23494
rect 24012 23546 24068 23548
rect 24012 23494 24014 23546
rect 24014 23494 24066 23546
rect 24066 23494 24068 23546
rect 24012 23492 24068 23494
rect 23804 21978 23860 21980
rect 23804 21926 23806 21978
rect 23806 21926 23858 21978
rect 23858 21926 23860 21978
rect 23804 21924 23860 21926
rect 23908 21978 23964 21980
rect 23908 21926 23910 21978
rect 23910 21926 23962 21978
rect 23962 21926 23964 21978
rect 23908 21924 23964 21926
rect 24012 21978 24068 21980
rect 24012 21926 24014 21978
rect 24014 21926 24066 21978
rect 24066 21926 24068 21978
rect 24012 21924 24068 21926
rect 23996 21698 24052 21700
rect 23996 21646 23998 21698
rect 23998 21646 24050 21698
rect 24050 21646 24052 21698
rect 23996 21644 24052 21646
rect 23804 20410 23860 20412
rect 23804 20358 23806 20410
rect 23806 20358 23858 20410
rect 23858 20358 23860 20410
rect 23804 20356 23860 20358
rect 23908 20410 23964 20412
rect 23908 20358 23910 20410
rect 23910 20358 23962 20410
rect 23962 20358 23964 20410
rect 23908 20356 23964 20358
rect 24012 20410 24068 20412
rect 24012 20358 24014 20410
rect 24014 20358 24066 20410
rect 24066 20358 24068 20410
rect 24012 20356 24068 20358
rect 24332 26124 24388 26180
rect 24464 25898 24520 25900
rect 24464 25846 24466 25898
rect 24466 25846 24518 25898
rect 24518 25846 24520 25898
rect 24464 25844 24520 25846
rect 24568 25898 24624 25900
rect 24568 25846 24570 25898
rect 24570 25846 24622 25898
rect 24622 25846 24624 25898
rect 24568 25844 24624 25846
rect 24672 25898 24728 25900
rect 24672 25846 24674 25898
rect 24674 25846 24726 25898
rect 24726 25846 24728 25898
rect 24672 25844 24728 25846
rect 24668 24444 24724 24500
rect 24464 24330 24520 24332
rect 24464 24278 24466 24330
rect 24466 24278 24518 24330
rect 24518 24278 24520 24330
rect 24464 24276 24520 24278
rect 24568 24330 24624 24332
rect 24568 24278 24570 24330
rect 24570 24278 24622 24330
rect 24622 24278 24624 24330
rect 24568 24276 24624 24278
rect 24672 24330 24728 24332
rect 24672 24278 24674 24330
rect 24674 24278 24726 24330
rect 24726 24278 24728 24330
rect 24672 24276 24728 24278
rect 24892 23212 24948 23268
rect 24464 22762 24520 22764
rect 24464 22710 24466 22762
rect 24466 22710 24518 22762
rect 24518 22710 24520 22762
rect 24464 22708 24520 22710
rect 24568 22762 24624 22764
rect 24568 22710 24570 22762
rect 24570 22710 24622 22762
rect 24622 22710 24624 22762
rect 24568 22708 24624 22710
rect 24672 22762 24728 22764
rect 24672 22710 24674 22762
rect 24674 22710 24726 22762
rect 24726 22710 24728 22762
rect 24672 22708 24728 22710
rect 25900 57260 25956 57316
rect 26236 57260 26292 57316
rect 25788 56700 25844 56756
rect 25676 54460 25732 54516
rect 25676 53618 25732 53620
rect 25676 53566 25678 53618
rect 25678 53566 25730 53618
rect 25730 53566 25732 53618
rect 25676 53564 25732 53566
rect 25452 52668 25508 52724
rect 25676 51772 25732 51828
rect 27580 56588 27636 56644
rect 26012 56306 26068 56308
rect 26012 56254 26014 56306
rect 26014 56254 26066 56306
rect 26066 56254 26068 56306
rect 26012 56252 26068 56254
rect 26236 55298 26292 55300
rect 26236 55246 26238 55298
rect 26238 55246 26290 55298
rect 26290 55246 26292 55298
rect 26236 55244 26292 55246
rect 26236 53116 26292 53172
rect 26236 52332 26292 52388
rect 26236 51100 26292 51156
rect 26236 50706 26292 50708
rect 26236 50654 26238 50706
rect 26238 50654 26290 50706
rect 26290 50654 26292 50706
rect 26236 50652 26292 50654
rect 25676 50482 25732 50484
rect 25676 50430 25678 50482
rect 25678 50430 25730 50482
rect 25730 50430 25732 50482
rect 25676 50428 25732 50430
rect 25676 49532 25732 49588
rect 26236 49196 26292 49252
rect 26236 48860 26292 48916
rect 25676 48636 25732 48692
rect 26236 47458 26292 47460
rect 26236 47406 26238 47458
rect 26238 47406 26290 47458
rect 26290 47406 26292 47458
rect 26236 47404 26292 47406
rect 25676 47346 25732 47348
rect 25676 47294 25678 47346
rect 25678 47294 25730 47346
rect 25730 47294 25732 47346
rect 25676 47292 25732 47294
rect 25676 46396 25732 46452
rect 26236 46060 26292 46116
rect 25676 45500 25732 45556
rect 25564 44268 25620 44324
rect 25452 36988 25508 37044
rect 25676 44210 25732 44212
rect 25676 44158 25678 44210
rect 25678 44158 25730 44210
rect 25730 44158 25732 44210
rect 25676 44156 25732 44158
rect 25676 43260 25732 43316
rect 25676 42364 25732 42420
rect 25676 41074 25732 41076
rect 25676 41022 25678 41074
rect 25678 41022 25730 41074
rect 25730 41022 25732 41074
rect 25676 41020 25732 41022
rect 26236 44994 26292 44996
rect 26236 44942 26238 44994
rect 26238 44942 26290 44994
rect 26290 44942 26292 44994
rect 26236 44940 26292 44942
rect 26236 44322 26292 44324
rect 26236 44270 26238 44322
rect 26238 44270 26290 44322
rect 26290 44270 26292 44322
rect 26236 44268 26292 44270
rect 27244 54012 27300 54068
rect 27020 53116 27076 53172
rect 26460 48412 26516 48468
rect 26572 52108 26628 52164
rect 25788 40236 25844 40292
rect 25676 40124 25732 40180
rect 25676 39228 25732 39284
rect 25676 37938 25732 37940
rect 25676 37886 25678 37938
rect 25678 37886 25730 37938
rect 25730 37886 25732 37938
rect 25676 37884 25732 37886
rect 25676 36092 25732 36148
rect 25564 35756 25620 35812
rect 25788 35084 25844 35140
rect 25676 34802 25732 34804
rect 25676 34750 25678 34802
rect 25678 34750 25730 34802
rect 25730 34750 25732 34802
rect 25676 34748 25732 34750
rect 25676 33852 25732 33908
rect 25676 32956 25732 33012
rect 25676 31666 25732 31668
rect 25676 31614 25678 31666
rect 25678 31614 25730 31666
rect 25730 31614 25732 31666
rect 25676 31612 25732 31614
rect 25452 30716 25508 30772
rect 25788 29372 25844 29428
rect 25788 29148 25844 29204
rect 25676 27132 25732 27188
rect 25116 26460 25172 26516
rect 25228 26236 25284 26292
rect 24220 19404 24276 19460
rect 24332 22092 24388 22148
rect 23804 18842 23860 18844
rect 23804 18790 23806 18842
rect 23806 18790 23858 18842
rect 23858 18790 23860 18842
rect 23804 18788 23860 18790
rect 23908 18842 23964 18844
rect 23908 18790 23910 18842
rect 23910 18790 23962 18842
rect 23962 18790 23964 18842
rect 23908 18788 23964 18790
rect 24012 18842 24068 18844
rect 24012 18790 24014 18842
rect 24014 18790 24066 18842
rect 24066 18790 24068 18842
rect 24012 18788 24068 18790
rect 23324 17724 23380 17780
rect 22988 15260 23044 15316
rect 23660 18450 23716 18452
rect 23660 18398 23662 18450
rect 23662 18398 23714 18450
rect 23714 18398 23716 18450
rect 23660 18396 23716 18398
rect 23804 17274 23860 17276
rect 23804 17222 23806 17274
rect 23806 17222 23858 17274
rect 23858 17222 23860 17274
rect 23804 17220 23860 17222
rect 23908 17274 23964 17276
rect 23908 17222 23910 17274
rect 23910 17222 23962 17274
rect 23962 17222 23964 17274
rect 23908 17220 23964 17222
rect 24012 17274 24068 17276
rect 24012 17222 24014 17274
rect 24014 17222 24066 17274
rect 24066 17222 24068 17274
rect 24012 17220 24068 17222
rect 23548 17052 23604 17108
rect 23804 15706 23860 15708
rect 23804 15654 23806 15706
rect 23806 15654 23858 15706
rect 23858 15654 23860 15706
rect 23804 15652 23860 15654
rect 23908 15706 23964 15708
rect 23908 15654 23910 15706
rect 23910 15654 23962 15706
rect 23962 15654 23964 15706
rect 23908 15652 23964 15654
rect 24012 15706 24068 15708
rect 24012 15654 24014 15706
rect 24014 15654 24066 15706
rect 24066 15654 24068 15706
rect 24012 15652 24068 15654
rect 23660 15036 23716 15092
rect 23804 14138 23860 14140
rect 23804 14086 23806 14138
rect 23806 14086 23858 14138
rect 23858 14086 23860 14138
rect 23804 14084 23860 14086
rect 23908 14138 23964 14140
rect 23908 14086 23910 14138
rect 23910 14086 23962 14138
rect 23962 14086 23964 14138
rect 23908 14084 23964 14086
rect 24012 14138 24068 14140
rect 24012 14086 24014 14138
rect 24014 14086 24066 14138
rect 24066 14086 24068 14138
rect 24012 14084 24068 14086
rect 23324 13132 23380 13188
rect 23772 13468 23828 13524
rect 25004 21756 25060 21812
rect 24464 21194 24520 21196
rect 24464 21142 24466 21194
rect 24466 21142 24518 21194
rect 24518 21142 24520 21194
rect 24464 21140 24520 21142
rect 24568 21194 24624 21196
rect 24568 21142 24570 21194
rect 24570 21142 24622 21194
rect 24622 21142 24624 21194
rect 24568 21140 24624 21142
rect 24672 21194 24728 21196
rect 24672 21142 24674 21194
rect 24674 21142 24726 21194
rect 24726 21142 24728 21194
rect 24672 21140 24728 21142
rect 24464 19626 24520 19628
rect 24464 19574 24466 19626
rect 24466 19574 24518 19626
rect 24518 19574 24520 19626
rect 24464 19572 24520 19574
rect 24568 19626 24624 19628
rect 24568 19574 24570 19626
rect 24570 19574 24622 19626
rect 24622 19574 24624 19626
rect 24568 19572 24624 19574
rect 24672 19626 24728 19628
rect 24672 19574 24674 19626
rect 24674 19574 24726 19626
rect 24726 19574 24728 19626
rect 24672 19572 24728 19574
rect 24464 18058 24520 18060
rect 24464 18006 24466 18058
rect 24466 18006 24518 18058
rect 24518 18006 24520 18058
rect 24464 18004 24520 18006
rect 24568 18058 24624 18060
rect 24568 18006 24570 18058
rect 24570 18006 24622 18058
rect 24622 18006 24624 18058
rect 24568 18004 24624 18006
rect 24672 18058 24728 18060
rect 24672 18006 24674 18058
rect 24674 18006 24726 18058
rect 24726 18006 24728 18058
rect 24672 18004 24728 18006
rect 24556 17778 24612 17780
rect 24556 17726 24558 17778
rect 24558 17726 24610 17778
rect 24610 17726 24612 17778
rect 24556 17724 24612 17726
rect 25340 20524 25396 20580
rect 25228 17724 25284 17780
rect 25340 19068 25396 19124
rect 24464 16490 24520 16492
rect 24464 16438 24466 16490
rect 24466 16438 24518 16490
rect 24518 16438 24520 16490
rect 24464 16436 24520 16438
rect 24568 16490 24624 16492
rect 24568 16438 24570 16490
rect 24570 16438 24622 16490
rect 24622 16438 24624 16490
rect 24568 16436 24624 16438
rect 24672 16490 24728 16492
rect 24672 16438 24674 16490
rect 24674 16438 24726 16490
rect 24726 16438 24728 16490
rect 24672 16436 24728 16438
rect 24464 14922 24520 14924
rect 24464 14870 24466 14922
rect 24466 14870 24518 14922
rect 24518 14870 24520 14922
rect 24464 14868 24520 14870
rect 24568 14922 24624 14924
rect 24568 14870 24570 14922
rect 24570 14870 24622 14922
rect 24622 14870 24624 14922
rect 24568 14868 24624 14870
rect 24672 14922 24728 14924
rect 24672 14870 24674 14922
rect 24674 14870 24726 14922
rect 24726 14870 24728 14922
rect 24672 14868 24728 14870
rect 24220 13692 24276 13748
rect 23660 12572 23716 12628
rect 24332 13580 24388 13636
rect 24892 13692 24948 13748
rect 24464 13354 24520 13356
rect 24464 13302 24466 13354
rect 24466 13302 24518 13354
rect 24518 13302 24520 13354
rect 24464 13300 24520 13302
rect 24568 13354 24624 13356
rect 24568 13302 24570 13354
rect 24570 13302 24622 13354
rect 24622 13302 24624 13354
rect 24568 13300 24624 13302
rect 24672 13354 24728 13356
rect 24672 13302 24674 13354
rect 24674 13302 24726 13354
rect 24726 13302 24728 13354
rect 24672 13300 24728 13302
rect 25228 13746 25284 13748
rect 25228 13694 25230 13746
rect 25230 13694 25282 13746
rect 25282 13694 25284 13746
rect 25228 13692 25284 13694
rect 25228 13468 25284 13524
rect 24220 12684 24276 12740
rect 23804 12570 23860 12572
rect 23804 12518 23806 12570
rect 23806 12518 23858 12570
rect 23858 12518 23860 12570
rect 23804 12516 23860 12518
rect 23908 12570 23964 12572
rect 23908 12518 23910 12570
rect 23910 12518 23962 12570
rect 23962 12518 23964 12570
rect 23908 12516 23964 12518
rect 24012 12570 24068 12572
rect 24012 12518 24014 12570
rect 24014 12518 24066 12570
rect 24066 12518 24068 12570
rect 24012 12516 24068 12518
rect 23212 11788 23268 11844
rect 23660 11788 23716 11844
rect 24464 11786 24520 11788
rect 24464 11734 24466 11786
rect 24466 11734 24518 11786
rect 24518 11734 24520 11786
rect 24464 11732 24520 11734
rect 24568 11786 24624 11788
rect 24568 11734 24570 11786
rect 24570 11734 24622 11786
rect 24622 11734 24624 11786
rect 24568 11732 24624 11734
rect 24672 11786 24728 11788
rect 24672 11734 24674 11786
rect 24674 11734 24726 11786
rect 24726 11734 24728 11786
rect 24672 11732 24728 11734
rect 23772 11506 23828 11508
rect 23772 11454 23774 11506
rect 23774 11454 23826 11506
rect 23826 11454 23828 11506
rect 23772 11452 23828 11454
rect 25004 11116 25060 11172
rect 23804 11002 23860 11004
rect 23804 10950 23806 11002
rect 23806 10950 23858 11002
rect 23858 10950 23860 11002
rect 23804 10948 23860 10950
rect 23908 11002 23964 11004
rect 23908 10950 23910 11002
rect 23910 10950 23962 11002
rect 23962 10950 23964 11002
rect 23908 10948 23964 10950
rect 24012 11002 24068 11004
rect 24012 10950 24014 11002
rect 24014 10950 24066 11002
rect 24066 10950 24068 11002
rect 24012 10948 24068 10950
rect 22988 10556 23044 10612
rect 24464 10218 24520 10220
rect 24464 10166 24466 10218
rect 24466 10166 24518 10218
rect 24518 10166 24520 10218
rect 24464 10164 24520 10166
rect 24568 10218 24624 10220
rect 24568 10166 24570 10218
rect 24570 10166 24622 10218
rect 24622 10166 24624 10218
rect 24568 10164 24624 10166
rect 24672 10218 24728 10220
rect 24672 10166 24674 10218
rect 24674 10166 24726 10218
rect 24726 10166 24728 10218
rect 24672 10164 24728 10166
rect 22876 9772 22932 9828
rect 22540 8258 22596 8260
rect 22540 8206 22542 8258
rect 22542 8206 22594 8258
rect 22594 8206 22596 8258
rect 22540 8204 22596 8206
rect 25116 9714 25172 9716
rect 25116 9662 25118 9714
rect 25118 9662 25170 9714
rect 25170 9662 25172 9714
rect 25116 9660 25172 9662
rect 23804 9434 23860 9436
rect 23804 9382 23806 9434
rect 23806 9382 23858 9434
rect 23858 9382 23860 9434
rect 23804 9380 23860 9382
rect 23908 9434 23964 9436
rect 23908 9382 23910 9434
rect 23910 9382 23962 9434
rect 23962 9382 23964 9434
rect 23908 9380 23964 9382
rect 24012 9434 24068 9436
rect 24012 9382 24014 9434
rect 24014 9382 24066 9434
rect 24066 9382 24068 9434
rect 24012 9380 24068 9382
rect 24464 8650 24520 8652
rect 24464 8598 24466 8650
rect 24466 8598 24518 8650
rect 24518 8598 24520 8650
rect 24464 8596 24520 8598
rect 24568 8650 24624 8652
rect 24568 8598 24570 8650
rect 24570 8598 24622 8650
rect 24622 8598 24624 8650
rect 24568 8596 24624 8598
rect 24672 8650 24728 8652
rect 24672 8598 24674 8650
rect 24674 8598 24726 8650
rect 24726 8598 24728 8650
rect 24672 8596 24728 8598
rect 22876 8204 22932 8260
rect 23804 7866 23860 7868
rect 23804 7814 23806 7866
rect 23806 7814 23858 7866
rect 23858 7814 23860 7866
rect 23804 7812 23860 7814
rect 23908 7866 23964 7868
rect 23908 7814 23910 7866
rect 23910 7814 23962 7866
rect 23962 7814 23964 7866
rect 23908 7812 23964 7814
rect 24012 7866 24068 7868
rect 24012 7814 24014 7866
rect 24014 7814 24066 7866
rect 24066 7814 24068 7866
rect 24012 7812 24068 7814
rect 22652 7532 22708 7588
rect 22540 7420 22596 7476
rect 24464 7082 24520 7084
rect 24464 7030 24466 7082
rect 24466 7030 24518 7082
rect 24518 7030 24520 7082
rect 24464 7028 24520 7030
rect 24568 7082 24624 7084
rect 24568 7030 24570 7082
rect 24570 7030 24622 7082
rect 24622 7030 24624 7082
rect 24568 7028 24624 7030
rect 24672 7082 24728 7084
rect 24672 7030 24674 7082
rect 24674 7030 24726 7082
rect 24726 7030 24728 7082
rect 24672 7028 24728 7030
rect 23324 6636 23380 6692
rect 23804 6298 23860 6300
rect 23804 6246 23806 6298
rect 23806 6246 23858 6298
rect 23858 6246 23860 6298
rect 23804 6244 23860 6246
rect 23908 6298 23964 6300
rect 23908 6246 23910 6298
rect 23910 6246 23962 6298
rect 23962 6246 23964 6298
rect 23908 6244 23964 6246
rect 24012 6298 24068 6300
rect 24012 6246 24014 6298
rect 24014 6246 24066 6298
rect 24066 6246 24068 6298
rect 24012 6244 24068 6246
rect 24892 5852 24948 5908
rect 24464 5514 24520 5516
rect 24464 5462 24466 5514
rect 24466 5462 24518 5514
rect 24518 5462 24520 5514
rect 24464 5460 24520 5462
rect 24568 5514 24624 5516
rect 24568 5462 24570 5514
rect 24570 5462 24622 5514
rect 24622 5462 24624 5514
rect 24568 5460 24624 5462
rect 24672 5514 24728 5516
rect 24672 5462 24674 5514
rect 24674 5462 24726 5514
rect 24726 5462 24728 5514
rect 24672 5460 24728 5462
rect 23804 4730 23860 4732
rect 23804 4678 23806 4730
rect 23806 4678 23858 4730
rect 23858 4678 23860 4730
rect 23804 4676 23860 4678
rect 23908 4730 23964 4732
rect 23908 4678 23910 4730
rect 23910 4678 23962 4730
rect 23962 4678 23964 4730
rect 23908 4676 23964 4678
rect 24012 4730 24068 4732
rect 24012 4678 24014 4730
rect 24014 4678 24066 4730
rect 24066 4678 24068 4730
rect 24012 4676 24068 4678
rect 24464 3946 24520 3948
rect 24464 3894 24466 3946
rect 24466 3894 24518 3946
rect 24518 3894 24520 3946
rect 24464 3892 24520 3894
rect 24568 3946 24624 3948
rect 24568 3894 24570 3946
rect 24570 3894 24622 3946
rect 24622 3894 24624 3946
rect 24568 3892 24624 3894
rect 24672 3946 24728 3948
rect 24672 3894 24674 3946
rect 24674 3894 24726 3946
rect 24726 3894 24728 3946
rect 24672 3892 24728 3894
rect 23804 3162 23860 3164
rect 23804 3110 23806 3162
rect 23806 3110 23858 3162
rect 23858 3110 23860 3162
rect 23804 3108 23860 3110
rect 23908 3162 23964 3164
rect 23908 3110 23910 3162
rect 23910 3110 23962 3162
rect 23962 3110 23964 3162
rect 23908 3108 23964 3110
rect 24012 3162 24068 3164
rect 24012 3110 24014 3162
rect 24014 3110 24066 3162
rect 24066 3110 24068 3162
rect 24012 3108 24068 3110
rect 24464 2378 24520 2380
rect 24464 2326 24466 2378
rect 24466 2326 24518 2378
rect 24518 2326 24520 2378
rect 24464 2324 24520 2326
rect 24568 2378 24624 2380
rect 24568 2326 24570 2378
rect 24570 2326 24622 2378
rect 24622 2326 24624 2378
rect 24568 2324 24624 2326
rect 24672 2378 24728 2380
rect 24672 2326 24674 2378
rect 24674 2326 24726 2378
rect 24726 2326 24728 2378
rect 24672 2324 24728 2326
rect 23324 2156 23380 2212
rect 23804 1594 23860 1596
rect 23804 1542 23806 1594
rect 23806 1542 23858 1594
rect 23858 1542 23860 1594
rect 23804 1540 23860 1542
rect 23908 1594 23964 1596
rect 23908 1542 23910 1594
rect 23910 1542 23962 1594
rect 23962 1542 23964 1594
rect 23908 1540 23964 1542
rect 24012 1594 24068 1596
rect 24012 1542 24014 1594
rect 24014 1542 24066 1594
rect 24066 1542 24068 1594
rect 24012 1540 24068 1542
rect 22428 1372 22484 1428
rect 25340 11676 25396 11732
rect 25676 26236 25732 26292
rect 25676 24892 25732 24948
rect 25564 23996 25620 24052
rect 25676 23100 25732 23156
rect 25564 22876 25620 22932
rect 25676 21756 25732 21812
rect 25564 20076 25620 20132
rect 25452 11452 25508 11508
rect 25340 11340 25396 11396
rect 25340 7420 25396 7476
rect 25676 14476 25732 14532
rect 25676 9996 25732 10052
rect 25676 9212 25732 9268
rect 25564 5740 25620 5796
rect 26012 41692 26068 41748
rect 26236 42754 26292 42756
rect 26236 42702 26238 42754
rect 26238 42702 26290 42754
rect 26290 42702 26292 42754
rect 26236 42700 26292 42702
rect 26236 41858 26292 41860
rect 26236 41806 26238 41858
rect 26238 41806 26290 41858
rect 26290 41806 26292 41858
rect 26236 41804 26292 41806
rect 26124 41356 26180 41412
rect 26236 40402 26292 40404
rect 26236 40350 26238 40402
rect 26238 40350 26290 40402
rect 26290 40350 26292 40402
rect 26236 40348 26292 40350
rect 26236 39004 26292 39060
rect 26236 38722 26292 38724
rect 26236 38670 26238 38722
rect 26238 38670 26290 38722
rect 26290 38670 26292 38722
rect 26236 38668 26292 38670
rect 26236 38050 26292 38052
rect 26236 37998 26238 38050
rect 26238 37998 26290 38050
rect 26290 37998 26292 38050
rect 26236 37996 26292 37998
rect 26124 36316 26180 36372
rect 26236 35868 26292 35924
rect 26236 34636 26292 34692
rect 26124 34300 26180 34356
rect 26124 32732 26180 32788
rect 26236 32620 26292 32676
rect 26460 34972 26516 35028
rect 26460 32562 26516 32564
rect 26460 32510 26462 32562
rect 26462 32510 26514 32562
rect 26514 32510 26516 32562
rect 26460 32508 26516 32510
rect 26460 31778 26516 31780
rect 26460 31726 26462 31778
rect 26462 31726 26514 31778
rect 26514 31726 26516 31778
rect 26460 31724 26516 31726
rect 26348 31388 26404 31444
rect 26236 30380 26292 30436
rect 26236 29426 26292 29428
rect 26236 29374 26238 29426
rect 26238 29374 26290 29426
rect 26290 29374 26292 29426
rect 26236 29372 26292 29374
rect 26348 29260 26404 29316
rect 26236 28642 26292 28644
rect 26236 28590 26238 28642
rect 26238 28590 26290 28642
rect 26290 28590 26292 28642
rect 26236 28588 26292 28590
rect 26124 28476 26180 28532
rect 26124 27916 26180 27972
rect 26236 27746 26292 27748
rect 26236 27694 26238 27746
rect 26238 27694 26290 27746
rect 26290 27694 26292 27746
rect 26236 27692 26292 27694
rect 26236 27074 26292 27076
rect 26236 27022 26238 27074
rect 26238 27022 26290 27074
rect 26290 27022 26292 27074
rect 26236 27020 26292 27022
rect 26236 26178 26292 26180
rect 26236 26126 26238 26178
rect 26238 26126 26290 26178
rect 26290 26126 26292 26178
rect 26236 26124 26292 26126
rect 26236 25676 26292 25732
rect 26236 23938 26292 23940
rect 26236 23886 26238 23938
rect 26238 23886 26290 23938
rect 26290 23886 26292 23938
rect 26236 23884 26292 23886
rect 25900 21644 25956 21700
rect 26124 23772 26180 23828
rect 25900 21308 25956 21364
rect 26236 23042 26292 23044
rect 26236 22990 26238 23042
rect 26238 22990 26290 23042
rect 26290 22990 26292 23042
rect 26236 22988 26292 22990
rect 26236 22540 26292 22596
rect 26236 21586 26292 21588
rect 26236 21534 26238 21586
rect 26238 21534 26290 21586
rect 26290 21534 26292 21586
rect 26236 21532 26292 21534
rect 25900 20802 25956 20804
rect 25900 20750 25902 20802
rect 25902 20750 25954 20802
rect 25954 20750 25956 20802
rect 25900 20748 25956 20750
rect 26012 20018 26068 20020
rect 26012 19966 26014 20018
rect 26014 19966 26066 20018
rect 26066 19966 26068 20018
rect 26012 19964 26068 19966
rect 26012 19740 26068 19796
rect 25900 19346 25956 19348
rect 25900 19294 25902 19346
rect 25902 19294 25954 19346
rect 25954 19294 25956 19346
rect 25900 19292 25956 19294
rect 25900 18620 25956 18676
rect 26012 17778 26068 17780
rect 26012 17726 26014 17778
rect 26014 17726 26066 17778
rect 26066 17726 26068 17778
rect 26012 17724 26068 17726
rect 26012 16994 26068 16996
rect 26012 16942 26014 16994
rect 26014 16942 26066 16994
rect 26066 16942 26068 16994
rect 26012 16940 26068 16942
rect 26012 15820 26068 15876
rect 26012 15148 26068 15204
rect 26236 15148 26292 15204
rect 27244 52220 27300 52276
rect 27132 51324 27188 51380
rect 27244 50876 27300 50932
rect 27020 49980 27076 50036
rect 27244 49084 27300 49140
rect 27132 48188 27188 48244
rect 27244 47740 27300 47796
rect 27356 48412 27412 48468
rect 27020 46844 27076 46900
rect 27244 45948 27300 46004
rect 27132 45052 27188 45108
rect 27244 44604 27300 44660
rect 27020 43708 27076 43764
rect 26908 41916 26964 41972
rect 27020 40572 27076 40628
rect 27020 38892 27076 38948
rect 26572 22428 26628 22484
rect 26684 37324 26740 37380
rect 27244 42812 27300 42868
rect 27244 41468 27300 41524
rect 27468 41132 27524 41188
rect 27244 39676 27300 39732
rect 27244 38332 27300 38388
rect 27020 37436 27076 37492
rect 26908 36540 26964 36596
rect 27132 35644 27188 35700
rect 27244 35196 27300 35252
rect 27020 34300 27076 34356
rect 27244 33404 27300 33460
rect 27132 32508 27188 32564
rect 27132 32284 27188 32340
rect 27244 32060 27300 32116
rect 27020 31164 27076 31220
rect 27132 30268 27188 30324
rect 27020 29820 27076 29876
rect 26908 29484 26964 29540
rect 27132 29372 27188 29428
rect 27020 28924 27076 28980
rect 27132 28530 27188 28532
rect 27132 28478 27134 28530
rect 27134 28478 27186 28530
rect 27186 28478 27188 28530
rect 27132 28476 27188 28478
rect 27132 28028 27188 28084
rect 27020 27580 27076 27636
rect 27244 26684 27300 26740
rect 27132 25564 27188 25620
rect 27244 25788 27300 25844
rect 27132 25340 27188 25396
rect 27468 32284 27524 32340
rect 27356 24556 27412 24612
rect 27468 31724 27524 31780
rect 27244 24444 27300 24500
rect 27132 23548 27188 23604
rect 27244 22652 27300 22708
rect 27132 22204 27188 22260
rect 27692 30940 27748 30996
rect 26684 20860 26740 20916
rect 26908 20802 26964 20804
rect 26908 20750 26910 20802
rect 26910 20750 26962 20802
rect 26962 20750 26964 20802
rect 26908 20748 26964 20750
rect 26572 20412 26628 20468
rect 26796 20188 26852 20244
rect 26460 19346 26516 19348
rect 26460 19294 26462 19346
rect 26462 19294 26514 19346
rect 26514 19294 26516 19346
rect 26460 19292 26516 19294
rect 26908 19906 26964 19908
rect 26908 19854 26910 19906
rect 26910 19854 26962 19906
rect 26962 19854 26964 19906
rect 26908 19852 26964 19854
rect 26908 18956 26964 19012
rect 26572 18450 26628 18452
rect 26572 18398 26574 18450
rect 26574 18398 26626 18450
rect 26626 18398 26628 18450
rect 26572 18396 26628 18398
rect 26908 18338 26964 18340
rect 26908 18286 26910 18338
rect 26910 18286 26962 18338
rect 26962 18286 26964 18338
rect 26908 18284 26964 18286
rect 26908 17836 26964 17892
rect 26572 17778 26628 17780
rect 26572 17726 26574 17778
rect 26574 17726 26626 17778
rect 26626 17726 26628 17778
rect 26572 17724 26628 17726
rect 26908 17500 26964 17556
rect 26572 16882 26628 16884
rect 26572 16830 26574 16882
rect 26574 16830 26626 16882
rect 26626 16830 26628 16882
rect 26572 16828 26628 16830
rect 26908 16210 26964 16212
rect 26908 16158 26910 16210
rect 26910 16158 26962 16210
rect 26962 16158 26964 16210
rect 26908 16156 26964 16158
rect 26572 15932 26628 15988
rect 26908 15484 26964 15540
rect 26684 15372 26740 15428
rect 26572 15090 26628 15092
rect 26572 15038 26574 15090
rect 26574 15038 26626 15090
rect 26626 15038 26628 15090
rect 26572 15036 26628 15038
rect 26348 14476 26404 14532
rect 26348 14306 26404 14308
rect 26348 14254 26350 14306
rect 26350 14254 26402 14306
rect 26402 14254 26404 14306
rect 26348 14252 26404 14254
rect 26572 13746 26628 13748
rect 26572 13694 26574 13746
rect 26574 13694 26626 13746
rect 26626 13694 26628 13746
rect 26572 13692 26628 13694
rect 26572 13468 26628 13524
rect 26012 12348 26068 12404
rect 26012 12178 26068 12180
rect 26012 12126 26014 12178
rect 26014 12126 26066 12178
rect 26066 12126 26068 12178
rect 26012 12124 26068 12126
rect 25900 11676 25956 11732
rect 26012 11564 26068 11620
rect 26236 11228 26292 11284
rect 26012 9100 26068 9156
rect 25900 8818 25956 8820
rect 25900 8766 25902 8818
rect 25902 8766 25954 8818
rect 25954 8766 25956 8818
rect 25900 8764 25956 8766
rect 26012 8428 26068 8484
rect 26124 7420 26180 7476
rect 26012 6802 26068 6804
rect 26012 6750 26014 6802
rect 26014 6750 26066 6802
rect 26066 6750 26068 6802
rect 26012 6748 26068 6750
rect 25900 5682 25956 5684
rect 25900 5630 25902 5682
rect 25902 5630 25954 5682
rect 25954 5630 25956 5682
rect 25900 5628 25956 5630
rect 26348 9884 26404 9940
rect 26572 12796 26628 12852
rect 26572 11954 26628 11956
rect 26572 11902 26574 11954
rect 26574 11902 26626 11954
rect 26626 11902 26628 11954
rect 26572 11900 26628 11902
rect 26572 11004 26628 11060
rect 26572 10108 26628 10164
rect 26572 9660 26628 9716
rect 26460 8988 26516 9044
rect 27020 14476 27076 14532
rect 27020 13858 27076 13860
rect 27020 13806 27022 13858
rect 27022 13806 27074 13858
rect 27074 13806 27076 13858
rect 27020 13804 27076 13806
rect 26908 12066 26964 12068
rect 26908 12014 26910 12066
rect 26910 12014 26962 12066
rect 26962 12014 26964 12066
rect 26908 12012 26964 12014
rect 26908 11506 26964 11508
rect 26908 11454 26910 11506
rect 26910 11454 26962 11506
rect 26962 11454 26964 11506
rect 26908 11452 26964 11454
rect 26908 10892 26964 10948
rect 27132 12572 27188 12628
rect 26684 7420 26740 7476
rect 26908 7644 26964 7700
rect 26572 6524 26628 6580
rect 27020 7586 27076 7588
rect 27020 7534 27022 7586
rect 27022 7534 27074 7586
rect 27074 7534 27076 7586
rect 27020 7532 27076 7534
rect 26684 6076 26740 6132
rect 25564 2716 25620 2772
rect 26684 5234 26740 5236
rect 26684 5182 26686 5234
rect 26686 5182 26738 5234
rect 26738 5182 26740 5234
rect 26684 5180 26740 5182
rect 26908 4226 26964 4228
rect 26908 4174 26910 4226
rect 26910 4174 26962 4226
rect 26962 4174 26964 4226
rect 26908 4172 26964 4174
rect 26908 3666 26964 3668
rect 26908 3614 26910 3666
rect 26910 3614 26962 3666
rect 26962 3614 26964 3666
rect 26908 3612 26964 3614
rect 26572 2940 26628 2996
rect 27468 21308 27524 21364
rect 27356 20914 27412 20916
rect 27356 20862 27358 20914
rect 27358 20862 27410 20914
rect 27410 20862 27412 20914
rect 27356 20860 27412 20862
rect 27580 20860 27636 20916
rect 27356 19516 27412 19572
rect 27580 19068 27636 19124
rect 27356 18172 27412 18228
rect 27692 18284 27748 18340
rect 27804 25564 27860 25620
rect 27580 17276 27636 17332
rect 27356 16380 27412 16436
rect 27580 15484 27636 15540
rect 27692 15260 27748 15316
rect 27356 14588 27412 14644
rect 27468 14140 27524 14196
rect 27356 13244 27412 13300
rect 27468 12908 27524 12964
rect 27468 12236 27524 12292
rect 27580 12348 27636 12404
rect 27356 11452 27412 11508
rect 27692 10892 27748 10948
rect 27580 10556 27636 10612
rect 28028 23660 28084 23716
rect 27916 20748 27972 20804
rect 27244 9324 27300 9380
rect 27468 9548 27524 9604
rect 27244 8316 27300 8372
rect 27244 8092 27300 8148
rect 27580 8204 27636 8260
rect 27692 9324 27748 9380
rect 27356 7420 27412 7476
rect 27468 7362 27524 7364
rect 27468 7310 27470 7362
rect 27470 7310 27522 7362
rect 27522 7310 27524 7362
rect 27468 7308 27524 7310
rect 27468 6972 27524 7028
rect 27356 5180 27412 5236
rect 27468 4732 27524 4788
rect 27244 4284 27300 4340
rect 27468 4338 27524 4340
rect 27468 4286 27470 4338
rect 27470 4286 27522 4338
rect 27522 4286 27524 4338
rect 27468 4284 27524 4286
rect 27468 3836 27524 3892
rect 28252 20524 28308 20580
rect 28028 16156 28084 16212
rect 28140 16940 28196 16996
rect 28028 15820 28084 15876
rect 28028 12572 28084 12628
rect 27692 5292 27748 5348
rect 28028 12236 28084 12292
rect 28140 9548 28196 9604
rect 28140 7532 28196 7588
rect 27804 4844 27860 4900
rect 28252 4508 28308 4564
rect 27580 3612 27636 3668
rect 27692 4396 27748 4452
rect 27468 3388 27524 3444
rect 25228 1874 25284 1876
rect 25228 1822 25230 1874
rect 25230 1822 25282 1874
rect 25282 1822 25284 1874
rect 25228 1820 25284 1822
rect 25788 2044 25844 2100
rect 26572 2546 26628 2548
rect 26572 2494 26574 2546
rect 26574 2494 26626 2546
rect 26626 2494 26628 2546
rect 26572 2492 26628 2494
rect 27468 2156 27524 2212
rect 26012 1260 26068 1316
rect 26572 1372 26628 1428
rect 25564 1148 25620 1204
rect 23548 1036 23604 1092
rect 24464 810 24520 812
rect 24464 758 24466 810
rect 24466 758 24518 810
rect 24518 758 24520 810
rect 24464 756 24520 758
rect 24568 810 24624 812
rect 24568 758 24570 810
rect 24570 758 24622 810
rect 24622 758 24624 810
rect 24568 756 24624 758
rect 24672 810 24728 812
rect 24672 758 24674 810
rect 24674 758 24726 810
rect 24726 758 24728 810
rect 24672 756 24728 758
rect 25340 700 25396 756
rect 26236 588 26292 644
rect 24892 364 24948 420
rect 26348 252 26404 308
rect 27132 1596 27188 1652
rect 26908 140 26964 196
<< metal3 >>
rect 19506 57260 19516 57316
rect 19572 57260 19852 57316
rect 19908 57260 19918 57316
rect 25890 57260 25900 57316
rect 25956 57260 26236 57316
rect 26292 57260 26302 57316
rect 28448 57204 28560 57232
rect 24994 57148 25004 57204
rect 25060 57148 28560 57204
rect 28448 57120 28560 57148
rect 28448 56756 28560 56784
rect 25778 56700 25788 56756
rect 25844 56700 28560 56756
rect 28448 56672 28560 56700
rect 24322 56588 24332 56644
rect 24388 56588 27580 56644
rect 27636 56588 27646 56644
rect 3794 56420 3804 56476
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 4068 56420 4078 56476
rect 23794 56420 23804 56476
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 24068 56420 24078 56476
rect 28448 56308 28560 56336
rect 15474 56252 15484 56308
rect 15540 56252 16492 56308
rect 16548 56252 16558 56308
rect 20850 56252 20860 56308
rect 20916 56252 22204 56308
rect 22260 56252 22270 56308
rect 23538 56252 23548 56308
rect 23604 56252 24444 56308
rect 24500 56252 24510 56308
rect 24882 56252 24892 56308
rect 24948 56252 26012 56308
rect 26068 56252 26078 56308
rect 26236 56252 28560 56308
rect 26236 56196 26292 56252
rect 28448 56224 28560 56252
rect 22530 56140 22540 56196
rect 22596 56140 26292 56196
rect 3014 55916 3052 55972
rect 3108 55916 3118 55972
rect 14018 55916 14028 55972
rect 14084 55916 19628 55972
rect 19684 55916 19694 55972
rect 21270 55916 21308 55972
rect 21364 55916 21374 55972
rect 24210 55916 24220 55972
rect 24276 55916 25452 55972
rect 25508 55916 25518 55972
rect 28448 55860 28560 55888
rect 6178 55804 6188 55860
rect 6244 55804 14700 55860
rect 14756 55804 14766 55860
rect 21634 55804 21644 55860
rect 21700 55804 28560 55860
rect 28448 55776 28560 55804
rect 4454 55636 4464 55692
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4728 55636 4738 55692
rect 24454 55636 24464 55692
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24728 55636 24738 55692
rect 28448 55412 28560 55440
rect 23538 55356 23548 55412
rect 23604 55356 28560 55412
rect 28448 55328 28560 55356
rect 1362 55244 1372 55300
rect 1428 55244 10220 55300
rect 10276 55244 10286 55300
rect 18274 55244 18284 55300
rect 18340 55244 20524 55300
rect 20580 55244 20590 55300
rect 22390 55244 22428 55300
rect 22484 55244 22494 55300
rect 24882 55244 24892 55300
rect 24948 55244 25340 55300
rect 25396 55244 25406 55300
rect 26114 55244 26124 55300
rect 26180 55244 26236 55300
rect 26292 55244 26302 55300
rect 0 55188 112 55216
rect 0 55132 1036 55188
rect 1092 55132 1102 55188
rect 6066 55132 6076 55188
rect 6132 55132 6860 55188
rect 6916 55132 6926 55188
rect 11442 55132 11452 55188
rect 11508 55132 11900 55188
rect 11956 55132 11966 55188
rect 0 55104 112 55132
rect 28448 54964 28560 54992
rect 26124 54908 28560 54964
rect 3794 54852 3804 54908
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 4068 54852 4078 54908
rect 23794 54852 23804 54908
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 24068 54852 24078 54908
rect 26124 54740 26180 54908
rect 28448 54880 28560 54908
rect 23762 54684 23772 54740
rect 23828 54684 26180 54740
rect 28448 54516 28560 54544
rect 11554 54460 11564 54516
rect 11620 54460 21196 54516
rect 21252 54460 21262 54516
rect 21746 54460 21756 54516
rect 21812 54460 24108 54516
rect 24164 54460 24174 54516
rect 25666 54460 25676 54516
rect 25732 54460 28560 54516
rect 28448 54432 28560 54460
rect 0 54292 112 54320
rect 0 54236 1036 54292
rect 1092 54236 1102 54292
rect 11890 54236 11900 54292
rect 11956 54236 20636 54292
rect 20692 54236 20702 54292
rect 0 54208 112 54236
rect 4454 54068 4464 54124
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4728 54068 4738 54124
rect 24454 54068 24464 54124
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24728 54068 24738 54124
rect 28448 54068 28560 54096
rect 21970 54012 21980 54068
rect 22036 54012 23660 54068
rect 23716 54012 23726 54068
rect 27234 54012 27244 54068
rect 27300 54012 28560 54068
rect 28448 53984 28560 54012
rect 12562 53900 12572 53956
rect 12628 53900 24892 53956
rect 24948 53900 24958 53956
rect 14354 53788 14364 53844
rect 14420 53788 20860 53844
rect 20916 53788 20926 53844
rect 16818 53676 16828 53732
rect 16884 53676 22764 53732
rect 22820 53676 22830 53732
rect 28448 53620 28560 53648
rect 17266 53564 17276 53620
rect 17332 53564 24668 53620
rect 24724 53564 24734 53620
rect 25666 53564 25676 53620
rect 25732 53564 28560 53620
rect 28448 53536 28560 53564
rect 0 53396 112 53424
rect 0 53340 1036 53396
rect 1092 53340 1102 53396
rect 0 53312 112 53340
rect 3794 53284 3804 53340
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 4068 53284 4078 53340
rect 23794 53284 23804 53340
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 24068 53284 24078 53340
rect 28448 53172 28560 53200
rect 11106 53116 11116 53172
rect 11172 53116 26236 53172
rect 26292 53116 26302 53172
rect 27010 53116 27020 53172
rect 27076 53116 28560 53172
rect 28448 53088 28560 53116
rect 12562 52780 12572 52836
rect 12628 52780 24668 52836
rect 24724 52780 24734 52836
rect 28448 52724 28560 52752
rect 23650 52668 23660 52724
rect 23716 52668 25004 52724
rect 25060 52668 25070 52724
rect 25442 52668 25452 52724
rect 25508 52668 28560 52724
rect 28448 52640 28560 52668
rect 0 52500 112 52528
rect 4454 52500 4464 52556
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4728 52500 4738 52556
rect 24454 52500 24464 52556
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24728 52500 24738 52556
rect 0 52444 1036 52500
rect 1092 52444 1102 52500
rect 0 52416 112 52444
rect 10882 52332 10892 52388
rect 10948 52332 26236 52388
rect 26292 52332 26302 52388
rect 28448 52276 28560 52304
rect 27234 52220 27244 52276
rect 27300 52220 28560 52276
rect 28448 52192 28560 52220
rect 1586 52108 1596 52164
rect 1652 52108 9100 52164
rect 9156 52108 9166 52164
rect 20850 52108 20860 52164
rect 20916 52108 21420 52164
rect 21476 52108 21486 52164
rect 22726 52108 22764 52164
rect 22820 52108 22830 52164
rect 24882 52108 24892 52164
rect 24948 52108 26572 52164
rect 26628 52108 26638 52164
rect 28448 51828 28560 51856
rect 25666 51772 25676 51828
rect 25732 51772 28560 51828
rect 3794 51716 3804 51772
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 4068 51716 4078 51772
rect 23794 51716 23804 51772
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 24068 51716 24078 51772
rect 28448 51744 28560 51772
rect 0 51604 112 51632
rect 0 51548 1036 51604
rect 1092 51548 1102 51604
rect 0 51520 112 51548
rect 28448 51380 28560 51408
rect 27122 51324 27132 51380
rect 27188 51324 28560 51380
rect 28448 51296 28560 51324
rect 1586 51212 1596 51268
rect 1652 51212 5852 51268
rect 5908 51212 5918 51268
rect 7746 51212 7756 51268
rect 7812 51212 24668 51268
rect 24724 51212 24734 51268
rect 14130 51100 14140 51156
rect 14196 51100 26236 51156
rect 26292 51100 26302 51156
rect 4454 50932 4464 50988
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4728 50932 4738 50988
rect 24454 50932 24464 50988
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24728 50932 24738 50988
rect 28448 50932 28560 50960
rect 27234 50876 27244 50932
rect 27300 50876 28560 50932
rect 28448 50848 28560 50876
rect 22418 50764 22428 50820
rect 22484 50764 27020 50820
rect 27076 50764 27086 50820
rect 0 50708 112 50736
rect 0 50652 924 50708
rect 980 50652 990 50708
rect 10770 50652 10780 50708
rect 10836 50652 26236 50708
rect 26292 50652 26302 50708
rect 0 50624 112 50652
rect 18386 50540 18396 50596
rect 18452 50540 23884 50596
rect 23940 50540 23950 50596
rect 28448 50484 28560 50512
rect 1586 50428 1596 50484
rect 1652 50428 2380 50484
rect 2436 50428 2446 50484
rect 16034 50428 16044 50484
rect 16100 50428 24668 50484
rect 24724 50428 24734 50484
rect 25666 50428 25676 50484
rect 25732 50428 28560 50484
rect 28448 50400 28560 50428
rect 3794 50148 3804 50204
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 4068 50148 4078 50204
rect 23794 50148 23804 50204
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 24068 50148 24078 50204
rect 28448 50036 28560 50064
rect 27010 49980 27020 50036
rect 27076 49980 28560 50036
rect 28448 49952 28560 49980
rect 0 49812 112 49840
rect 0 49756 1036 49812
rect 1092 49756 1102 49812
rect 0 49728 112 49756
rect 9202 49644 9212 49700
rect 9268 49644 24668 49700
rect 24724 49644 24734 49700
rect 28448 49588 28560 49616
rect 25666 49532 25676 49588
rect 25732 49532 28560 49588
rect 28448 49504 28560 49532
rect 4454 49364 4464 49420
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4728 49364 4738 49420
rect 24454 49364 24464 49420
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24728 49364 24738 49420
rect 16258 49196 16268 49252
rect 16324 49196 26236 49252
rect 26292 49196 26302 49252
rect 28448 49140 28560 49168
rect 27234 49084 27244 49140
rect 27300 49084 28560 49140
rect 28448 49056 28560 49084
rect 6290 48972 6300 49028
rect 6356 48972 24668 49028
rect 24724 48972 24734 49028
rect 0 48916 112 48944
rect 0 48860 1036 48916
rect 1092 48860 1102 48916
rect 14802 48860 14812 48916
rect 14868 48860 26236 48916
rect 26292 48860 26302 48916
rect 0 48832 112 48860
rect 28448 48692 28560 48720
rect 25666 48636 25676 48692
rect 25732 48636 28560 48692
rect 3794 48580 3804 48636
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 4068 48580 4078 48636
rect 23794 48580 23804 48636
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 24068 48580 24078 48636
rect 28448 48608 28560 48636
rect 1138 48412 1148 48468
rect 1204 48412 5628 48468
rect 5684 48412 5694 48468
rect 26450 48412 26460 48468
rect 26516 48412 27356 48468
rect 27412 48412 27422 48468
rect 28448 48244 28560 48272
rect 27122 48188 27132 48244
rect 27188 48188 28560 48244
rect 28448 48160 28560 48188
rect 802 48076 812 48132
rect 868 48076 1596 48132
rect 1652 48076 1662 48132
rect 16706 48076 16716 48132
rect 16772 48076 19964 48132
rect 20020 48076 20030 48132
rect 0 48020 112 48048
rect 0 47964 1036 48020
rect 1092 47964 1102 48020
rect 0 47936 112 47964
rect 4454 47796 4464 47852
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4728 47796 4738 47852
rect 24454 47796 24464 47852
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24728 47796 24738 47852
rect 28448 47796 28560 47824
rect 27234 47740 27244 47796
rect 27300 47740 28560 47796
rect 28448 47712 28560 47740
rect 19282 47404 19292 47460
rect 19348 47404 24668 47460
rect 24724 47404 24734 47460
rect 24892 47404 26236 47460
rect 26292 47404 26302 47460
rect 24892 47348 24948 47404
rect 28448 47348 28560 47376
rect 19730 47292 19740 47348
rect 19796 47292 24948 47348
rect 25666 47292 25676 47348
rect 25732 47292 28560 47348
rect 28448 47264 28560 47292
rect 0 47124 112 47152
rect 0 47068 1036 47124
rect 1092 47068 1102 47124
rect 0 47040 112 47068
rect 3794 47012 3804 47068
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 4068 47012 4078 47068
rect 23794 47012 23804 47068
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 24068 47012 24078 47068
rect 12450 46956 12460 47012
rect 12516 46956 16828 47012
rect 16884 46956 16894 47012
rect 28448 46900 28560 46928
rect 27010 46844 27020 46900
rect 27076 46844 28560 46900
rect 28448 46816 28560 46844
rect 1586 46508 1596 46564
rect 1652 46508 8876 46564
rect 8932 46508 8942 46564
rect 17938 46508 17948 46564
rect 18004 46508 24668 46564
rect 24724 46508 24734 46564
rect 28448 46452 28560 46480
rect 25666 46396 25676 46452
rect 25732 46396 28560 46452
rect 28448 46368 28560 46396
rect 1446 46284 1484 46340
rect 1540 46284 1550 46340
rect 0 46228 112 46256
rect 4454 46228 4464 46284
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4728 46228 4738 46284
rect 24454 46228 24464 46284
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24728 46228 24738 46284
rect 0 46172 1932 46228
rect 1988 46172 1998 46228
rect 0 46144 112 46172
rect 16930 46060 16940 46116
rect 16996 46060 26236 46116
rect 26292 46060 26302 46116
rect 28448 46004 28560 46032
rect 27234 45948 27244 46004
rect 27300 45948 28560 46004
rect 28448 45920 28560 45948
rect 15698 45836 15708 45892
rect 15764 45836 24668 45892
rect 24724 45836 24734 45892
rect 1586 45724 1596 45780
rect 1652 45724 7644 45780
rect 7700 45724 7710 45780
rect 28448 45556 28560 45584
rect 25666 45500 25676 45556
rect 25732 45500 28560 45556
rect 3794 45444 3804 45500
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 4068 45444 4078 45500
rect 23794 45444 23804 45500
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 24068 45444 24078 45500
rect 28448 45472 28560 45500
rect 0 45332 112 45360
rect 0 45276 924 45332
rect 980 45276 990 45332
rect 9090 45276 9100 45332
rect 9156 45276 13692 45332
rect 13748 45276 13758 45332
rect 0 45248 112 45276
rect 28448 45108 28560 45136
rect 27122 45052 27132 45108
rect 27188 45052 28560 45108
rect 28448 45024 28560 45052
rect 8530 44940 8540 44996
rect 8596 44940 26236 44996
rect 26292 44940 26302 44996
rect 4454 44660 4464 44716
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4728 44660 4738 44716
rect 24454 44660 24464 44716
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24728 44660 24738 44716
rect 28448 44660 28560 44688
rect 27234 44604 27244 44660
rect 27300 44604 28560 44660
rect 28448 44576 28560 44604
rect 0 44436 112 44464
rect 0 44380 1148 44436
rect 1204 44380 1214 44436
rect 1558 44380 1596 44436
rect 1652 44380 1662 44436
rect 0 44352 112 44380
rect 20178 44268 20188 44324
rect 20244 44268 24668 44324
rect 24724 44268 24734 44324
rect 25554 44268 25564 44324
rect 25620 44268 26236 44324
rect 26292 44268 26302 44324
rect 28448 44212 28560 44240
rect 25666 44156 25676 44212
rect 25732 44156 28560 44212
rect 28448 44128 28560 44156
rect 3794 43876 3804 43932
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 4068 43876 4078 43932
rect 23794 43876 23804 43932
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 24068 43876 24078 43932
rect 28448 43764 28560 43792
rect 1586 43708 1596 43764
rect 1652 43708 1708 43764
rect 1764 43708 1774 43764
rect 27010 43708 27020 43764
rect 27076 43708 28560 43764
rect 28448 43680 28560 43708
rect 802 43596 812 43652
rect 868 43596 10780 43652
rect 10836 43596 10846 43652
rect 0 43540 112 43568
rect 0 43484 924 43540
rect 980 43484 990 43540
rect 0 43456 112 43484
rect 1586 43372 1596 43428
rect 1652 43372 2604 43428
rect 2660 43372 2670 43428
rect 28448 43316 28560 43344
rect 25666 43260 25676 43316
rect 25732 43260 28560 43316
rect 28448 43232 28560 43260
rect 4454 43092 4464 43148
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4728 43092 4738 43148
rect 24454 43092 24464 43148
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24728 43092 24738 43148
rect 2370 42924 2380 42980
rect 2436 42924 6748 42980
rect 6804 42924 6814 42980
rect 28448 42868 28560 42896
rect 1698 42812 1708 42868
rect 1764 42812 3388 42868
rect 8082 42812 8092 42868
rect 8148 42812 23324 42868
rect 23380 42812 23390 42868
rect 27234 42812 27244 42868
rect 27300 42812 28560 42868
rect 0 42644 112 42672
rect 0 42588 1148 42644
rect 1204 42588 1214 42644
rect 1698 42588 1708 42644
rect 1764 42588 2380 42644
rect 2436 42588 2446 42644
rect 0 42560 112 42588
rect 3332 42532 3388 42812
rect 28448 42784 28560 42812
rect 9762 42700 9772 42756
rect 9828 42700 26236 42756
rect 26292 42700 26302 42756
rect 9874 42588 9884 42644
rect 9940 42588 24668 42644
rect 24724 42588 24734 42644
rect 3332 42476 8652 42532
rect 8708 42476 8718 42532
rect 28448 42420 28560 42448
rect 25666 42364 25676 42420
rect 25732 42364 28560 42420
rect 3794 42308 3804 42364
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 4068 42308 4078 42364
rect 23794 42308 23804 42364
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 24068 42308 24078 42364
rect 28448 42336 28560 42364
rect 1372 42140 1596 42196
rect 1652 42140 1662 42196
rect 2034 42140 2044 42196
rect 2100 42140 8316 42196
rect 8372 42140 8382 42196
rect 1372 42084 1428 42140
rect 1362 42028 1372 42084
rect 1428 42028 1438 42084
rect 5506 42028 5516 42084
rect 5572 42028 8540 42084
rect 8596 42028 8606 42084
rect 28448 41972 28560 42000
rect 3042 41916 3052 41972
rect 3108 41916 10892 41972
rect 10948 41916 10958 41972
rect 14690 41916 14700 41972
rect 14756 41916 19852 41972
rect 19908 41916 19918 41972
rect 26898 41916 26908 41972
rect 26964 41916 28560 41972
rect 28448 41888 28560 41916
rect 1586 41804 1596 41860
rect 1652 41804 11228 41860
rect 11284 41804 11294 41860
rect 16706 41804 16716 41860
rect 16772 41804 26236 41860
rect 26292 41804 26302 41860
rect 0 41748 112 41776
rect 0 41692 1932 41748
rect 1988 41692 1998 41748
rect 15586 41692 15596 41748
rect 15652 41692 26012 41748
rect 26068 41692 26078 41748
rect 0 41664 112 41692
rect 1698 41580 1708 41636
rect 1764 41580 2268 41636
rect 2324 41580 2334 41636
rect 4454 41524 4464 41580
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4728 41524 4738 41580
rect 24454 41524 24464 41580
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24728 41524 24738 41580
rect 28448 41524 28560 41552
rect 5506 41468 5516 41524
rect 5572 41468 14364 41524
rect 14420 41468 14430 41524
rect 27234 41468 27244 41524
rect 27300 41468 28560 41524
rect 28448 41440 28560 41468
rect 5842 41356 5852 41412
rect 5908 41356 13244 41412
rect 13300 41356 13310 41412
rect 15026 41356 15036 41412
rect 15092 41356 26124 41412
rect 26180 41356 26190 41412
rect 1586 41244 1596 41300
rect 1652 41244 8428 41300
rect 10098 41244 10108 41300
rect 10164 41244 10892 41300
rect 10948 41244 10958 41300
rect 11116 41244 20076 41300
rect 20132 41244 20142 41300
rect 8372 41188 8428 41244
rect 11116 41188 11172 41244
rect 8372 41132 11172 41188
rect 11778 41132 11788 41188
rect 11844 41132 27468 41188
rect 27524 41132 27534 41188
rect 28448 41076 28560 41104
rect 242 41020 252 41076
rect 308 41020 1596 41076
rect 1652 41020 1662 41076
rect 7858 41020 7868 41076
rect 7924 41020 12124 41076
rect 12180 41020 13916 41076
rect 13972 41020 14364 41076
rect 14420 41020 14430 41076
rect 25666 41020 25676 41076
rect 25732 41020 28560 41076
rect 28448 40992 28560 41020
rect 0 40852 112 40880
rect 0 40796 1820 40852
rect 1876 40796 1886 40852
rect 0 40768 112 40796
rect 3794 40740 3804 40796
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 4068 40740 4078 40796
rect 23794 40740 23804 40796
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 24068 40740 24078 40796
rect 28448 40628 28560 40656
rect 1362 40572 1372 40628
rect 1428 40572 13468 40628
rect 13524 40572 13534 40628
rect 27010 40572 27020 40628
rect 27076 40572 28560 40628
rect 28448 40544 28560 40572
rect 2482 40460 2492 40516
rect 2548 40460 16044 40516
rect 16100 40460 16110 40516
rect 14578 40348 14588 40404
rect 14644 40348 26236 40404
rect 26292 40348 26302 40404
rect 690 40236 700 40292
rect 756 40236 1596 40292
rect 1652 40236 1662 40292
rect 2146 40236 2156 40292
rect 2212 40236 5964 40292
rect 6020 40236 6030 40292
rect 12226 40236 12236 40292
rect 12292 40236 25788 40292
rect 25844 40236 25854 40292
rect 28448 40180 28560 40208
rect 6066 40124 6076 40180
rect 6132 40124 6300 40180
rect 6356 40124 6366 40180
rect 12114 40124 12124 40180
rect 12180 40124 14252 40180
rect 14308 40124 14318 40180
rect 18386 40124 18396 40180
rect 18452 40124 24780 40180
rect 24836 40124 24846 40180
rect 25666 40124 25676 40180
rect 25732 40124 28560 40180
rect 28448 40096 28560 40124
rect 12898 40012 12908 40068
rect 12964 40012 21084 40068
rect 21140 40012 21150 40068
rect 0 39956 112 39984
rect 4454 39956 4464 40012
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4728 39956 4738 40012
rect 24454 39956 24464 40012
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24728 39956 24738 40012
rect 0 39900 2044 39956
rect 2100 39900 2110 39956
rect 9538 39900 9548 39956
rect 9604 39900 24332 39956
rect 24388 39900 24398 39956
rect 0 39872 112 39900
rect 2258 39788 2268 39844
rect 2324 39788 2492 39844
rect 2548 39788 5852 39844
rect 5908 39788 5918 39844
rect 7298 39788 7308 39844
rect 7364 39788 12572 39844
rect 12628 39788 12638 39844
rect 28448 39732 28560 39760
rect 3490 39676 3500 39732
rect 3556 39676 7308 39732
rect 7364 39676 7374 39732
rect 9986 39676 9996 39732
rect 10052 39676 26908 39732
rect 26964 39676 26974 39732
rect 27234 39676 27244 39732
rect 27300 39676 28560 39732
rect 28448 39648 28560 39676
rect 3938 39564 3948 39620
rect 4004 39564 8428 39620
rect 8484 39564 8494 39620
rect 22306 39564 22316 39620
rect 22372 39564 24668 39620
rect 24724 39564 24734 39620
rect 6402 39452 6412 39508
rect 6468 39452 11788 39508
rect 11844 39452 14476 39508
rect 14532 39452 14542 39508
rect 3490 39340 3500 39396
rect 3556 39340 5180 39396
rect 5236 39340 6636 39396
rect 6692 39340 10444 39396
rect 10500 39340 10510 39396
rect 28448 39284 28560 39312
rect 5394 39228 5404 39284
rect 5460 39228 14140 39284
rect 14196 39228 14206 39284
rect 25666 39228 25676 39284
rect 25732 39228 28560 39284
rect 3794 39172 3804 39228
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 4068 39172 4078 39228
rect 23794 39172 23804 39228
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 24068 39172 24078 39228
rect 28448 39200 28560 39228
rect 8754 39116 8764 39172
rect 8820 39116 15596 39172
rect 15652 39116 15662 39172
rect 0 39060 112 39088
rect 0 39004 364 39060
rect 420 39004 430 39060
rect 7858 39004 7868 39060
rect 7924 39004 8204 39060
rect 8260 39004 10108 39060
rect 10164 39004 10174 39060
rect 17378 39004 17388 39060
rect 17444 39004 26236 39060
rect 26292 39004 26302 39060
rect 0 38976 112 39004
rect 1586 38892 1596 38948
rect 1652 38892 12572 38948
rect 12628 38892 12638 38948
rect 27010 38892 27020 38948
rect 27076 38892 27086 38948
rect 27020 38836 27076 38892
rect 28448 38836 28560 38864
rect 6850 38780 6860 38836
rect 6916 38780 8764 38836
rect 8820 38780 8830 38836
rect 10098 38780 10108 38836
rect 10164 38780 13580 38836
rect 13636 38780 13646 38836
rect 13906 38780 13916 38836
rect 13972 38780 14812 38836
rect 14868 38780 14878 38836
rect 15250 38780 15260 38836
rect 15316 38780 15820 38836
rect 15876 38780 15886 38836
rect 27020 38780 28560 38836
rect 28448 38752 28560 38780
rect 6290 38668 6300 38724
rect 6356 38668 7980 38724
rect 8036 38668 8046 38724
rect 9202 38668 9212 38724
rect 9268 38668 9884 38724
rect 9940 38668 11004 38724
rect 11060 38668 11070 38724
rect 13346 38668 13356 38724
rect 13412 38668 13804 38724
rect 13860 38668 13870 38724
rect 19954 38668 19964 38724
rect 20020 38668 26236 38724
rect 26292 38668 26302 38724
rect 1698 38556 1708 38612
rect 1764 38556 2156 38612
rect 2212 38556 6860 38612
rect 6916 38556 6926 38612
rect 10434 38556 10444 38612
rect 10500 38556 10892 38612
rect 10948 38556 15148 38612
rect 15204 38556 15214 38612
rect 2706 38444 2716 38500
rect 2772 38444 4172 38500
rect 4228 38444 4238 38500
rect 13570 38444 13580 38500
rect 13636 38444 14924 38500
rect 14980 38444 14990 38500
rect 4454 38388 4464 38444
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4728 38388 4738 38444
rect 24454 38388 24464 38444
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24728 38388 24738 38444
rect 28448 38388 28560 38416
rect 27234 38332 27244 38388
rect 27300 38332 28560 38388
rect 28448 38304 28560 38332
rect 8194 38220 8204 38276
rect 8260 38220 13132 38276
rect 13188 38220 13198 38276
rect 15092 38220 24892 38276
rect 24948 38220 24958 38276
rect 0 38164 112 38192
rect 15092 38164 15148 38220
rect 0 38108 2828 38164
rect 2884 38108 2894 38164
rect 9538 38108 9548 38164
rect 9604 38108 15148 38164
rect 0 38080 112 38108
rect 1810 37996 1820 38052
rect 1876 37996 2492 38052
rect 2548 37996 2558 38052
rect 20738 37996 20748 38052
rect 20804 37996 26236 38052
rect 26292 37996 26302 38052
rect 28448 37940 28560 37968
rect 1922 37884 1932 37940
rect 1988 37884 2828 37940
rect 2884 37884 4732 37940
rect 4788 37884 4798 37940
rect 6514 37884 6524 37940
rect 6580 37884 23660 37940
rect 23716 37884 23726 37940
rect 25666 37884 25676 37940
rect 25732 37884 28560 37940
rect 28448 37856 28560 37884
rect 4386 37772 4396 37828
rect 4452 37772 5068 37828
rect 5124 37772 5404 37828
rect 5460 37772 5470 37828
rect 3794 37604 3804 37660
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 4068 37604 4078 37660
rect 23794 37604 23804 37660
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 24068 37604 24078 37660
rect 28448 37492 28560 37520
rect 27010 37436 27020 37492
rect 27076 37436 28560 37492
rect 28448 37408 28560 37436
rect 2706 37324 2716 37380
rect 2772 37324 4844 37380
rect 4900 37324 6524 37380
rect 6580 37324 10668 37380
rect 10724 37324 10734 37380
rect 12002 37324 12012 37380
rect 12068 37324 13020 37380
rect 13076 37324 17164 37380
rect 17220 37324 17230 37380
rect 17490 37324 17500 37380
rect 17556 37324 26684 37380
rect 26740 37324 26750 37380
rect 0 37268 112 37296
rect 0 37212 476 37268
rect 532 37212 542 37268
rect 8642 37212 8652 37268
rect 8708 37212 9660 37268
rect 9716 37212 9726 37268
rect 11778 37212 11788 37268
rect 11844 37212 12796 37268
rect 12852 37212 15932 37268
rect 15988 37212 15998 37268
rect 0 37184 112 37212
rect 1698 37100 1708 37156
rect 1764 37100 3388 37156
rect 4162 37100 4172 37156
rect 4228 37100 13580 37156
rect 13636 37100 13646 37156
rect 16482 37100 16492 37156
rect 16548 37100 24668 37156
rect 24724 37100 24734 37156
rect 3332 37044 3388 37100
rect 28448 37044 28560 37072
rect 3332 36988 13804 37044
rect 13860 36988 13870 37044
rect 25442 36988 25452 37044
rect 25508 36988 28560 37044
rect 28448 36960 28560 36988
rect 1474 36876 1484 36932
rect 1540 36876 1708 36932
rect 1764 36876 1774 36932
rect 4454 36820 4464 36876
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4728 36820 4738 36876
rect 24454 36820 24464 36876
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24728 36820 24738 36876
rect 354 36764 364 36820
rect 420 36764 812 36820
rect 868 36764 878 36820
rect 2258 36652 2268 36708
rect 2324 36652 2604 36708
rect 2660 36652 2670 36708
rect 16146 36652 16156 36708
rect 16212 36652 16716 36708
rect 16772 36652 16782 36708
rect 28448 36596 28560 36624
rect 3042 36540 3052 36596
rect 3108 36540 8764 36596
rect 8820 36540 8830 36596
rect 12562 36540 12572 36596
rect 12628 36540 17500 36596
rect 17556 36540 18284 36596
rect 18340 36540 18350 36596
rect 26898 36540 26908 36596
rect 26964 36540 28560 36596
rect 28448 36512 28560 36540
rect 3154 36428 3164 36484
rect 3220 36428 6412 36484
rect 6468 36428 6478 36484
rect 0 36372 112 36400
rect 0 36316 588 36372
rect 644 36316 654 36372
rect 2146 36316 2156 36372
rect 2212 36316 26124 36372
rect 26180 36316 26190 36372
rect 0 36288 112 36316
rect 19394 36204 19404 36260
rect 19460 36204 19852 36260
rect 19908 36204 19918 36260
rect 20076 36204 24892 36260
rect 24948 36204 24958 36260
rect 20076 36148 20132 36204
rect 28448 36148 28560 36176
rect 5394 36092 5404 36148
rect 5460 36092 20132 36148
rect 25666 36092 25676 36148
rect 25732 36092 28560 36148
rect 3794 36036 3804 36092
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 4068 36036 4078 36092
rect 23794 36036 23804 36092
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 24068 36036 24078 36092
rect 28448 36064 28560 36092
rect 8306 35868 8316 35924
rect 8372 35868 26236 35924
rect 26292 35868 26302 35924
rect 578 35756 588 35812
rect 644 35756 1372 35812
rect 1428 35756 2716 35812
rect 2772 35756 2782 35812
rect 6514 35756 6524 35812
rect 6580 35756 7980 35812
rect 8036 35756 8046 35812
rect 17266 35756 17276 35812
rect 17332 35756 25564 35812
rect 25620 35756 25630 35812
rect 28448 35700 28560 35728
rect 1222 35644 1260 35700
rect 1316 35644 1326 35700
rect 1586 35644 1596 35700
rect 1652 35644 3164 35700
rect 3220 35644 3230 35700
rect 4386 35644 4396 35700
rect 4452 35644 20188 35700
rect 20244 35644 20254 35700
rect 27122 35644 27132 35700
rect 27188 35644 28560 35700
rect 28448 35616 28560 35644
rect 2258 35532 2268 35588
rect 2324 35532 4844 35588
rect 4900 35532 4910 35588
rect 0 35476 112 35504
rect 0 35420 364 35476
rect 420 35420 430 35476
rect 2146 35420 2156 35476
rect 2212 35420 5292 35476
rect 5348 35420 5358 35476
rect 8642 35420 8652 35476
rect 8708 35420 9324 35476
rect 9380 35420 9390 35476
rect 0 35392 112 35420
rect 2594 35308 2604 35364
rect 2660 35308 3724 35364
rect 3780 35308 3790 35364
rect 9874 35308 9884 35364
rect 9940 35308 11116 35364
rect 11172 35308 11182 35364
rect 17490 35308 17500 35364
rect 17556 35308 18060 35364
rect 18116 35308 18126 35364
rect 4454 35252 4464 35308
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4728 35252 4738 35308
rect 24454 35252 24464 35308
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24728 35252 24738 35308
rect 28448 35252 28560 35280
rect 1922 35196 1932 35252
rect 1988 35196 2268 35252
rect 2324 35196 2334 35252
rect 2818 35196 2828 35252
rect 2884 35196 2940 35252
rect 2996 35196 3006 35252
rect 10434 35196 10444 35252
rect 10500 35196 16604 35252
rect 16660 35196 16670 35252
rect 27234 35196 27244 35252
rect 27300 35196 28560 35252
rect 28448 35168 28560 35196
rect 1334 35084 1372 35140
rect 1428 35084 1438 35140
rect 3602 35084 3612 35140
rect 3668 35084 9212 35140
rect 9268 35084 10668 35140
rect 10724 35084 10734 35140
rect 12674 35084 12684 35140
rect 12740 35084 25788 35140
rect 25844 35084 25854 35140
rect 1250 34972 1260 35028
rect 1316 34972 3948 35028
rect 4004 34972 4014 35028
rect 9314 34972 9324 35028
rect 9380 34972 26460 35028
rect 26516 34972 26526 35028
rect 5282 34860 5292 34916
rect 5348 34860 5852 34916
rect 5908 34860 5918 34916
rect 10854 34860 10892 34916
rect 10948 34860 10958 34916
rect 16258 34860 16268 34916
rect 16324 34860 19068 34916
rect 19124 34860 19134 34916
rect 28448 34804 28560 34832
rect 1586 34748 1596 34804
rect 1652 34748 10444 34804
rect 10500 34748 10510 34804
rect 15586 34748 15596 34804
rect 15652 34748 18284 34804
rect 18340 34748 18350 34804
rect 25666 34748 25676 34804
rect 25732 34748 28560 34804
rect 28448 34720 28560 34748
rect 8194 34636 8204 34692
rect 8260 34636 9100 34692
rect 9156 34636 9166 34692
rect 17042 34636 17052 34692
rect 17108 34636 26236 34692
rect 26292 34636 26302 34692
rect 0 34580 112 34608
rect 0 34524 1148 34580
rect 1204 34524 1214 34580
rect 7522 34524 7532 34580
rect 7588 34524 21868 34580
rect 21924 34524 21934 34580
rect 0 34496 112 34524
rect 3794 34468 3804 34524
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 4068 34468 4078 34524
rect 23794 34468 23804 34524
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 24068 34468 24078 34524
rect 1558 34412 1596 34468
rect 1652 34412 1662 34468
rect 2258 34412 2268 34468
rect 2324 34412 2334 34468
rect 4274 34412 4284 34468
rect 4340 34412 5292 34468
rect 5348 34412 5358 34468
rect 7074 34412 7084 34468
rect 7140 34412 8204 34468
rect 8260 34412 8270 34468
rect 8838 34412 8876 34468
rect 8932 34412 8942 34468
rect 14018 34412 14028 34468
rect 14084 34412 19964 34468
rect 20020 34412 20030 34468
rect 1362 34076 1372 34132
rect 1428 34076 1484 34132
rect 1540 34076 1550 34132
rect 2268 34020 2324 34412
rect 28448 34356 28560 34384
rect 4162 34300 4172 34356
rect 4228 34300 26124 34356
rect 26180 34300 26190 34356
rect 27010 34300 27020 34356
rect 27076 34300 28560 34356
rect 28448 34272 28560 34300
rect 2482 34188 2492 34244
rect 2548 34188 17836 34244
rect 17892 34188 17902 34244
rect 3378 34076 3388 34132
rect 3444 34076 4844 34132
rect 4900 34076 4910 34132
rect 5618 34076 5628 34132
rect 5684 34076 6300 34132
rect 6356 34076 6366 34132
rect 8082 34076 8092 34132
rect 8148 34076 10220 34132
rect 10276 34076 10286 34132
rect 11778 34076 11788 34132
rect 11844 34076 13356 34132
rect 13412 34076 21308 34132
rect 21364 34076 21374 34132
rect 2268 33964 2492 34020
rect 2548 33964 2558 34020
rect 8642 33964 8652 34020
rect 8708 33964 9660 34020
rect 9716 33964 9726 34020
rect 28448 33908 28560 33936
rect 1922 33852 1932 33908
rect 1988 33852 3612 33908
rect 3668 33852 3678 33908
rect 5058 33852 5068 33908
rect 5124 33852 5516 33908
rect 5572 33852 5582 33908
rect 6178 33852 6188 33908
rect 6244 33852 6972 33908
rect 7028 33852 7756 33908
rect 7812 33852 7822 33908
rect 15092 33852 24668 33908
rect 24724 33852 24734 33908
rect 25666 33852 25676 33908
rect 25732 33852 28560 33908
rect 15092 33796 15148 33852
rect 28448 33824 28560 33852
rect 6412 33740 15148 33796
rect 17714 33740 17724 33796
rect 17780 33740 18284 33796
rect 18340 33740 18350 33796
rect 0 33684 112 33712
rect 4454 33684 4464 33740
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4728 33684 4738 33740
rect 6412 33684 6468 33740
rect 24454 33684 24464 33740
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24728 33684 24738 33740
rect 0 33628 812 33684
rect 868 33628 878 33684
rect 1250 33628 1260 33684
rect 1316 33628 1484 33684
rect 1540 33628 1550 33684
rect 1698 33628 1708 33684
rect 1764 33628 2044 33684
rect 2100 33628 2110 33684
rect 2930 33628 2940 33684
rect 2996 33628 3052 33684
rect 3108 33628 3118 33684
rect 6402 33628 6412 33684
rect 6468 33628 6478 33684
rect 8642 33628 8652 33684
rect 8708 33628 8876 33684
rect 8932 33628 8942 33684
rect 9314 33628 9324 33684
rect 9380 33628 9660 33684
rect 9716 33628 9726 33684
rect 12674 33628 12684 33684
rect 12740 33628 13132 33684
rect 13188 33628 13198 33684
rect 17490 33628 17500 33684
rect 17556 33628 17836 33684
rect 17892 33628 18788 33684
rect 0 33600 112 33628
rect 18732 33572 18788 33628
rect 1138 33516 1148 33572
rect 1204 33516 2268 33572
rect 2324 33516 2716 33572
rect 2772 33516 15148 33572
rect 18722 33516 18732 33572
rect 18788 33516 19292 33572
rect 19348 33516 19358 33572
rect 2594 33404 2604 33460
rect 2660 33404 4284 33460
rect 4340 33404 4350 33460
rect 6738 33404 6748 33460
rect 6804 33404 6860 33460
rect 6916 33404 7644 33460
rect 7700 33404 8876 33460
rect 8932 33404 8942 33460
rect 578 33292 588 33348
rect 644 33292 1148 33348
rect 1204 33292 1214 33348
rect 3332 33292 7196 33348
rect 7252 33292 10892 33348
rect 10948 33292 10958 33348
rect 3332 33236 3388 33292
rect 1586 33180 1596 33236
rect 1652 33180 3388 33236
rect 15092 33236 15148 33516
rect 28448 33460 28560 33488
rect 27234 33404 27244 33460
rect 27300 33404 28560 33460
rect 28448 33376 28560 33404
rect 15092 33180 18956 33236
rect 19012 33180 19022 33236
rect 578 33068 588 33124
rect 644 33068 21532 33124
rect 21588 33068 21598 33124
rect 28448 33012 28560 33040
rect 11666 32956 11676 33012
rect 11732 32956 12684 33012
rect 12740 32956 12750 33012
rect 25666 32956 25676 33012
rect 25732 32956 28560 33012
rect 3794 32900 3804 32956
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 4068 32900 4078 32956
rect 23794 32900 23804 32956
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 24068 32900 24078 32956
rect 28448 32928 28560 32956
rect 8754 32844 8764 32900
rect 8820 32844 10220 32900
rect 10276 32844 10286 32900
rect 12002 32844 12012 32900
rect 12068 32844 12908 32900
rect 12964 32844 12974 32900
rect 0 32788 112 32816
rect 0 32732 1820 32788
rect 1876 32732 1886 32788
rect 4918 32732 4956 32788
rect 5012 32732 5022 32788
rect 8530 32732 8540 32788
rect 8596 32732 8606 32788
rect 11218 32732 11228 32788
rect 11284 32732 26124 32788
rect 26180 32732 26190 32788
rect 0 32704 112 32732
rect 8540 32676 8596 32732
rect 8540 32620 8764 32676
rect 8820 32620 8830 32676
rect 12562 32620 12572 32676
rect 12628 32620 15596 32676
rect 15652 32620 15662 32676
rect 22082 32620 22092 32676
rect 22148 32620 26236 32676
rect 26292 32620 26302 32676
rect 28448 32564 28560 32592
rect 13206 32508 13244 32564
rect 13300 32508 13310 32564
rect 13794 32508 13804 32564
rect 13860 32508 26460 32564
rect 26516 32508 26526 32564
rect 27122 32508 27132 32564
rect 27188 32508 28560 32564
rect 28448 32480 28560 32508
rect 1222 32396 1260 32452
rect 1316 32396 1708 32452
rect 1764 32396 1774 32452
rect 4274 32396 4284 32452
rect 4340 32396 7644 32452
rect 7700 32396 7710 32452
rect 1138 32284 1148 32340
rect 1204 32284 5516 32340
rect 5572 32284 5582 32340
rect 8866 32284 8876 32340
rect 8932 32284 15820 32340
rect 15876 32284 15886 32340
rect 27122 32284 27132 32340
rect 27188 32284 27468 32340
rect 27524 32284 27534 32340
rect 10882 32172 10892 32228
rect 10948 32172 14924 32228
rect 14980 32172 16380 32228
rect 16436 32172 16446 32228
rect 4454 32116 4464 32172
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4728 32116 4738 32172
rect 24454 32116 24464 32172
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24728 32116 24738 32172
rect 28448 32116 28560 32144
rect 12114 32060 12124 32116
rect 12180 32060 12908 32116
rect 12964 32060 12974 32116
rect 13430 32060 13468 32116
rect 13524 32060 13534 32116
rect 14130 32060 14140 32116
rect 14196 32060 15036 32116
rect 15092 32060 15102 32116
rect 27234 32060 27244 32116
rect 27300 32060 28560 32116
rect 28448 32032 28560 32060
rect 12786 31948 12796 32004
rect 12852 31948 13356 32004
rect 13412 31948 13422 32004
rect 15138 31948 15148 32004
rect 15204 31948 15932 32004
rect 15988 31948 15998 32004
rect 18050 31948 18060 32004
rect 18116 31948 18508 32004
rect 18564 31948 18574 32004
rect 21410 31948 21420 32004
rect 21476 31948 24220 32004
rect 24276 31948 24286 32004
rect 0 31892 112 31920
rect 0 31836 924 31892
rect 980 31836 990 31892
rect 2034 31836 2044 31892
rect 2100 31836 2492 31892
rect 2548 31836 2558 31892
rect 2706 31836 2716 31892
rect 2772 31836 4956 31892
rect 5012 31836 5022 31892
rect 5954 31836 5964 31892
rect 6020 31836 9660 31892
rect 9716 31836 9726 31892
rect 11106 31836 11116 31892
rect 11172 31836 12460 31892
rect 12516 31836 12526 31892
rect 13122 31836 13132 31892
rect 13188 31836 24780 31892
rect 24836 31836 24846 31892
rect 0 31808 112 31836
rect 1138 31724 1148 31780
rect 1204 31724 1260 31780
rect 1316 31724 1708 31780
rect 1764 31724 1774 31780
rect 3266 31724 3276 31780
rect 3332 31724 3612 31780
rect 3668 31724 3678 31780
rect 9090 31724 9100 31780
rect 9156 31724 14476 31780
rect 14532 31724 14542 31780
rect 16818 31724 16828 31780
rect 16884 31724 18060 31780
rect 18116 31724 18396 31780
rect 18452 31724 18462 31780
rect 20962 31724 20972 31780
rect 21028 31724 21532 31780
rect 21588 31724 21598 31780
rect 26450 31724 26460 31780
rect 26516 31724 27468 31780
rect 27524 31724 27534 31780
rect 5058 31612 5068 31668
rect 5124 31612 5628 31668
rect 5684 31612 5694 31668
rect 7382 31612 7420 31668
rect 7476 31612 7486 31668
rect 7970 31612 7980 31668
rect 8036 31612 8204 31668
rect 8260 31612 9884 31668
rect 9940 31612 9950 31668
rect 10630 31612 10668 31668
rect 10724 31612 10734 31668
rect 11330 31612 11340 31668
rect 11396 31612 12236 31668
rect 12292 31612 13580 31668
rect 13636 31612 13646 31668
rect 14476 31556 14532 31724
rect 28448 31668 28560 31696
rect 25666 31612 25676 31668
rect 25732 31612 28560 31668
rect 28448 31584 28560 31612
rect 14476 31500 20524 31556
rect 20580 31500 21308 31556
rect 21364 31500 21374 31556
rect 7298 31388 7308 31444
rect 7364 31388 23212 31444
rect 23268 31388 23660 31444
rect 23716 31388 23726 31444
rect 26310 31388 26348 31444
rect 26404 31388 26414 31444
rect 3794 31332 3804 31388
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 4068 31332 4078 31388
rect 23794 31332 23804 31388
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 24068 31332 24078 31388
rect 9996 31276 13244 31332
rect 13300 31276 13468 31332
rect 13524 31276 13534 31332
rect 4274 31164 4284 31220
rect 4340 31164 5404 31220
rect 5460 31164 5470 31220
rect 0 30996 112 31024
rect 9996 30996 10052 31276
rect 28448 31220 28560 31248
rect 10210 31164 10220 31220
rect 10276 31164 11228 31220
rect 11284 31164 11294 31220
rect 12226 31164 12236 31220
rect 12292 31164 13916 31220
rect 13972 31164 13982 31220
rect 15092 31164 24892 31220
rect 24948 31164 24958 31220
rect 27010 31164 27020 31220
rect 27076 31164 28560 31220
rect 15092 31108 15148 31164
rect 28448 31136 28560 31164
rect 11116 31052 15148 31108
rect 19954 31052 19964 31108
rect 20020 31052 20972 31108
rect 21028 31052 21038 31108
rect 0 30940 1036 30996
rect 1092 30940 1102 30996
rect 5516 30940 9996 30996
rect 10052 30940 10062 30996
rect 10546 30940 10556 30996
rect 10612 30940 10622 30996
rect 0 30912 112 30940
rect 5516 30884 5572 30940
rect 10556 30884 10612 30940
rect 5506 30828 5516 30884
rect 5572 30828 5582 30884
rect 5730 30828 5740 30884
rect 5796 30828 7308 30884
rect 7364 30828 7374 30884
rect 10098 30828 10108 30884
rect 10164 30828 10612 30884
rect 130 30716 140 30772
rect 196 30716 364 30772
rect 420 30716 3164 30772
rect 3220 30716 10892 30772
rect 10948 30716 10958 30772
rect 11116 30660 11172 31052
rect 11442 30940 11452 30996
rect 11508 30940 15708 30996
rect 15764 30940 18508 30996
rect 18564 30940 18574 30996
rect 19730 30940 19740 30996
rect 19796 30940 22092 30996
rect 22148 30940 22158 30996
rect 23650 30940 23660 30996
rect 23716 30940 27692 30996
rect 27748 30940 27758 30996
rect 13570 30828 13580 30884
rect 13636 30828 14364 30884
rect 14420 30828 14430 30884
rect 15026 30828 15036 30884
rect 15092 30828 16940 30884
rect 16996 30828 17006 30884
rect 18508 30772 18564 30940
rect 20178 30828 20188 30884
rect 20244 30828 20636 30884
rect 20692 30828 20702 30884
rect 28448 30772 28560 30800
rect 13682 30716 13692 30772
rect 13748 30716 14588 30772
rect 14644 30716 14654 30772
rect 18508 30716 22428 30772
rect 22484 30716 22494 30772
rect 25442 30716 25452 30772
rect 25508 30716 28560 30772
rect 28448 30688 28560 30716
rect 4946 30604 4956 30660
rect 5012 30604 5292 30660
rect 5348 30604 5358 30660
rect 10322 30604 10332 30660
rect 10388 30604 11172 30660
rect 13906 30604 13916 30660
rect 13972 30604 13982 30660
rect 4454 30548 4464 30604
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4728 30548 4738 30604
rect 13916 30548 13972 30604
rect 24454 30548 24464 30604
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24728 30548 24738 30604
rect 6860 30492 13972 30548
rect 17490 30492 17500 30548
rect 17556 30492 18508 30548
rect 18564 30492 18574 30548
rect 4386 30380 4396 30436
rect 4452 30380 6300 30436
rect 6356 30380 6366 30436
rect 6860 30324 6916 30492
rect 10994 30380 11004 30436
rect 11060 30380 11340 30436
rect 11396 30380 11406 30436
rect 12786 30380 12796 30436
rect 12852 30380 26236 30436
rect 26292 30380 26302 30436
rect 28448 30324 28560 30352
rect 1250 30268 1260 30324
rect 1316 30268 2716 30324
rect 2772 30268 2782 30324
rect 4162 30268 4172 30324
rect 4228 30268 6916 30324
rect 8082 30268 8092 30324
rect 8148 30268 12236 30324
rect 12292 30268 12302 30324
rect 13346 30268 13356 30324
rect 13412 30268 14308 30324
rect 17714 30268 17724 30324
rect 17780 30268 21644 30324
rect 21700 30268 21710 30324
rect 27122 30268 27132 30324
rect 27188 30268 28560 30324
rect 14252 30212 14308 30268
rect 28448 30240 28560 30268
rect 2258 30156 2268 30212
rect 2324 30156 2604 30212
rect 2660 30156 2670 30212
rect 4498 30156 4508 30212
rect 4564 30156 5068 30212
rect 5124 30156 5134 30212
rect 6514 30156 6524 30212
rect 6580 30156 9100 30212
rect 9156 30156 9166 30212
rect 9650 30156 9660 30212
rect 9716 30156 11676 30212
rect 11732 30156 11742 30212
rect 12114 30156 12124 30212
rect 12180 30156 14028 30212
rect 14084 30156 14094 30212
rect 14242 30156 14252 30212
rect 14308 30156 14318 30212
rect 17042 30156 17052 30212
rect 17108 30156 19292 30212
rect 19348 30156 20412 30212
rect 20468 30156 21420 30212
rect 21476 30156 21486 30212
rect 21746 30156 21756 30212
rect 21812 30156 23100 30212
rect 23156 30156 23166 30212
rect 0 30100 112 30128
rect 0 30044 1036 30100
rect 1092 30044 1102 30100
rect 1922 30044 1932 30100
rect 1988 30044 3164 30100
rect 3220 30044 4284 30100
rect 4340 30044 4350 30100
rect 8530 30044 8540 30100
rect 8596 30044 12908 30100
rect 12964 30044 12974 30100
rect 19058 30044 19068 30100
rect 19124 30044 19740 30100
rect 19796 30044 19806 30100
rect 20066 30044 20076 30100
rect 20132 30044 23548 30100
rect 23604 30044 23614 30100
rect 0 30016 112 30044
rect 3378 29932 3388 29988
rect 3444 29932 5068 29988
rect 5124 29932 5134 29988
rect 9426 29932 9436 29988
rect 9492 29932 9884 29988
rect 9940 29932 11340 29988
rect 11396 29932 17388 29988
rect 17444 29932 17454 29988
rect 17714 29932 17724 29988
rect 17780 29932 18620 29988
rect 18676 29932 18686 29988
rect 18946 29932 18956 29988
rect 19012 29932 19292 29988
rect 19348 29932 19358 29988
rect 28448 29876 28560 29904
rect 2930 29820 2940 29876
rect 2996 29820 3052 29876
rect 3108 29820 3118 29876
rect 14354 29820 14364 29876
rect 14420 29820 17052 29876
rect 17108 29820 17118 29876
rect 27010 29820 27020 29876
rect 27076 29820 28560 29876
rect 3794 29764 3804 29820
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 4068 29764 4078 29820
rect 14364 29764 14420 29820
rect 23794 29764 23804 29820
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 24068 29764 24078 29820
rect 28448 29792 28560 29820
rect 6962 29708 6972 29764
rect 7028 29708 7756 29764
rect 7812 29708 8092 29764
rect 8148 29708 10556 29764
rect 10612 29708 14420 29764
rect 15092 29708 21028 29764
rect 15092 29652 15148 29708
rect 20972 29652 21028 29708
rect 4274 29596 4284 29652
rect 4340 29596 4956 29652
rect 5012 29596 5022 29652
rect 6402 29596 6412 29652
rect 6468 29596 7196 29652
rect 7252 29596 7262 29652
rect 11554 29596 11564 29652
rect 11620 29596 11900 29652
rect 11956 29596 15148 29652
rect 15474 29596 15484 29652
rect 15540 29596 16716 29652
rect 16772 29596 16782 29652
rect 20972 29596 26908 29652
rect 4172 29484 7308 29540
rect 7364 29484 8540 29540
rect 8596 29484 8606 29540
rect 8764 29484 16940 29540
rect 16996 29484 17006 29540
rect 26852 29484 26908 29596
rect 26964 29484 26974 29540
rect 4172 29428 4228 29484
rect 8764 29428 8820 29484
rect 28448 29428 28560 29456
rect 2594 29372 2604 29428
rect 2660 29372 4172 29428
rect 4228 29372 4238 29428
rect 4918 29372 4956 29428
rect 5012 29372 5022 29428
rect 5282 29372 5292 29428
rect 5348 29372 5628 29428
rect 5684 29372 8820 29428
rect 10882 29372 10892 29428
rect 10948 29372 11004 29428
rect 11060 29372 11070 29428
rect 15138 29372 15148 29428
rect 15204 29372 15484 29428
rect 15540 29372 15550 29428
rect 15698 29372 15708 29428
rect 15764 29372 16380 29428
rect 16436 29372 16446 29428
rect 25778 29372 25788 29428
rect 25844 29372 26236 29428
rect 26292 29372 26302 29428
rect 27122 29372 27132 29428
rect 27188 29372 28560 29428
rect 28448 29344 28560 29372
rect 7410 29260 7420 29316
rect 7476 29260 8764 29316
rect 8820 29260 18060 29316
rect 18116 29260 18126 29316
rect 26310 29260 26348 29316
rect 26404 29260 26414 29316
rect 0 29204 112 29232
rect 0 29148 1036 29204
rect 1092 29148 1102 29204
rect 10966 29148 11004 29204
rect 11060 29148 11070 29204
rect 18834 29148 18844 29204
rect 18900 29148 25788 29204
rect 25844 29148 25854 29204
rect 0 29120 112 29148
rect 4454 28980 4464 29036
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4728 28980 4738 29036
rect 24454 28980 24464 29036
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24728 28980 24738 29036
rect 28448 28980 28560 29008
rect 1026 28924 1036 28980
rect 1092 28924 2604 28980
rect 2660 28924 2670 28980
rect 5170 28924 5180 28980
rect 5236 28924 6076 28980
rect 6132 28924 6142 28980
rect 13906 28924 13916 28980
rect 13972 28924 22988 28980
rect 23044 28924 23054 28980
rect 27010 28924 27020 28980
rect 27076 28924 28560 28980
rect 28448 28896 28560 28924
rect 3490 28812 3500 28868
rect 3556 28812 11564 28868
rect 11620 28812 11630 28868
rect 15698 28812 15708 28868
rect 15764 28812 16492 28868
rect 16548 28812 16558 28868
rect 17938 28812 17948 28868
rect 18004 28812 18508 28868
rect 18564 28812 18574 28868
rect 2342 28700 2380 28756
rect 2436 28700 2446 28756
rect 5170 28700 5180 28756
rect 5236 28700 5852 28756
rect 5908 28700 5918 28756
rect 8866 28700 8876 28756
rect 8932 28700 9100 28756
rect 9156 28700 9884 28756
rect 9940 28700 9950 28756
rect 11330 28700 11340 28756
rect 11396 28700 13804 28756
rect 13860 28700 13870 28756
rect 11106 28588 11116 28644
rect 11172 28588 11900 28644
rect 11956 28588 11966 28644
rect 13570 28588 13580 28644
rect 13636 28588 13916 28644
rect 13972 28588 13982 28644
rect 16034 28588 16044 28644
rect 16100 28588 26236 28644
rect 26292 28588 26302 28644
rect 28448 28532 28560 28560
rect 1474 28476 1484 28532
rect 1540 28476 2044 28532
rect 2100 28476 8092 28532
rect 8148 28476 8158 28532
rect 10546 28476 10556 28532
rect 10612 28476 11676 28532
rect 11732 28476 17388 28532
rect 17444 28476 17454 28532
rect 19170 28476 19180 28532
rect 19236 28476 26124 28532
rect 26180 28476 26190 28532
rect 27122 28476 27132 28532
rect 27188 28476 28560 28532
rect 28448 28448 28560 28476
rect 3332 28364 5628 28420
rect 5684 28364 5694 28420
rect 6514 28364 6524 28420
rect 6580 28364 7308 28420
rect 7364 28364 8876 28420
rect 8932 28364 8942 28420
rect 12114 28364 12124 28420
rect 12180 28364 13020 28420
rect 13076 28364 13086 28420
rect 16034 28364 16044 28420
rect 16100 28364 18732 28420
rect 18788 28364 18798 28420
rect 0 28308 112 28336
rect 3332 28308 3388 28364
rect 0 28252 3388 28308
rect 5954 28252 5964 28308
rect 6020 28252 7420 28308
rect 7476 28252 7486 28308
rect 7942 28252 7980 28308
rect 8036 28252 8046 28308
rect 12674 28252 12684 28308
rect 12740 28252 13580 28308
rect 13636 28252 13646 28308
rect 0 28224 112 28252
rect 3794 28196 3804 28252
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 4068 28196 4078 28252
rect 23794 28196 23804 28252
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 24068 28196 24078 28252
rect 5730 28140 5740 28196
rect 5796 28140 7644 28196
rect 7700 28140 7710 28196
rect 28448 28084 28560 28112
rect 7410 28028 7420 28084
rect 7476 28028 9548 28084
rect 9604 28028 10444 28084
rect 10500 28028 10510 28084
rect 10658 28028 10668 28084
rect 10724 28028 25004 28084
rect 25060 28028 25070 28084
rect 27122 28028 27132 28084
rect 27188 28028 28560 28084
rect 28448 28000 28560 28028
rect 11666 27916 11676 27972
rect 11732 27916 26124 27972
rect 26180 27916 26190 27972
rect 4946 27804 4956 27860
rect 5012 27804 5796 27860
rect 16594 27804 16604 27860
rect 16660 27804 17836 27860
rect 17892 27804 18172 27860
rect 18228 27804 18238 27860
rect 5740 27748 5796 27804
rect 5730 27692 5740 27748
rect 5796 27692 5806 27748
rect 8642 27692 8652 27748
rect 8708 27692 9548 27748
rect 9604 27692 11004 27748
rect 11060 27692 11070 27748
rect 13570 27692 13580 27748
rect 13636 27692 15148 27748
rect 26198 27692 26236 27748
rect 26292 27692 26302 27748
rect 15092 27524 15148 27692
rect 28448 27636 28560 27664
rect 17154 27580 17164 27636
rect 17220 27580 18060 27636
rect 18116 27580 18126 27636
rect 27010 27580 27020 27636
rect 27076 27580 28560 27636
rect 28448 27552 28560 27580
rect 15092 27468 16604 27524
rect 16660 27468 21532 27524
rect 21588 27468 21598 27524
rect 0 27412 112 27440
rect 4454 27412 4464 27468
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4728 27412 4738 27468
rect 24454 27412 24464 27468
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24728 27412 24738 27468
rect 0 27356 140 27412
rect 196 27356 206 27412
rect 5506 27356 5516 27412
rect 5572 27356 15148 27412
rect 0 27328 112 27356
rect 15092 27300 15148 27356
rect 1698 27244 1708 27300
rect 1764 27244 3164 27300
rect 3220 27244 3230 27300
rect 4274 27244 4284 27300
rect 4340 27244 4956 27300
rect 5012 27244 5022 27300
rect 10070 27244 10108 27300
rect 10164 27244 10174 27300
rect 11218 27244 11228 27300
rect 11284 27244 12012 27300
rect 12068 27244 12908 27300
rect 12964 27244 12974 27300
rect 13122 27244 13132 27300
rect 13188 27244 13916 27300
rect 13972 27244 13982 27300
rect 15092 27244 24892 27300
rect 24948 27244 24958 27300
rect 28448 27188 28560 27216
rect 2818 27132 2828 27188
rect 2884 27132 3276 27188
rect 3332 27132 3342 27188
rect 4050 27132 4060 27188
rect 4116 27132 5964 27188
rect 6020 27132 6030 27188
rect 13458 27132 13468 27188
rect 13524 27132 14140 27188
rect 14196 27132 14206 27188
rect 16706 27132 16716 27188
rect 16772 27132 17388 27188
rect 17444 27132 17454 27188
rect 21298 27132 21308 27188
rect 21364 27132 21532 27188
rect 21588 27132 21598 27188
rect 25666 27132 25676 27188
rect 25732 27132 28560 27188
rect 13916 27076 13972 27132
rect 28448 27104 28560 27132
rect 130 27020 140 27076
rect 196 27020 1036 27076
rect 1092 27020 1102 27076
rect 1250 27020 1260 27076
rect 1316 27020 1820 27076
rect 1876 27020 1886 27076
rect 5254 27020 5292 27076
rect 5348 27020 5358 27076
rect 13906 27020 13916 27076
rect 13972 27020 13982 27076
rect 14252 27020 26236 27076
rect 26292 27020 26302 27076
rect 14252 26964 14308 27020
rect 3266 26908 3276 26964
rect 3332 26908 5404 26964
rect 5460 26908 5470 26964
rect 7970 26908 7980 26964
rect 8036 26908 11564 26964
rect 11620 26908 11630 26964
rect 14242 26908 14252 26964
rect 14308 26908 14318 26964
rect 14690 26908 14700 26964
rect 14756 26908 15596 26964
rect 15652 26908 15662 26964
rect 22082 26908 22092 26964
rect 22148 26908 22316 26964
rect 22372 26908 22382 26964
rect 12002 26796 12012 26852
rect 12068 26796 15932 26852
rect 15988 26796 15998 26852
rect 16258 26796 16268 26852
rect 16324 26796 20188 26852
rect 20244 26796 20254 26852
rect 28448 26740 28560 26768
rect 5506 26684 5516 26740
rect 5572 26684 13132 26740
rect 13188 26684 13198 26740
rect 13990 26684 14028 26740
rect 14084 26684 14094 26740
rect 16268 26684 17500 26740
rect 17556 26684 17566 26740
rect 27234 26684 27244 26740
rect 27300 26684 28560 26740
rect 3794 26628 3804 26684
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 4068 26628 4078 26684
rect 16268 26628 16324 26684
rect 23794 26628 23804 26684
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 24068 26628 24078 26684
rect 28448 26656 28560 26684
rect 6402 26572 6412 26628
rect 6468 26572 6478 26628
rect 11106 26572 11116 26628
rect 11172 26572 16324 26628
rect 0 26516 112 26544
rect 6412 26516 6468 26572
rect 0 26460 1260 26516
rect 1316 26460 1326 26516
rect 3042 26460 3052 26516
rect 3108 26460 6468 26516
rect 13346 26460 13356 26516
rect 13412 26460 25116 26516
rect 25172 26460 25182 26516
rect 0 26432 112 26460
rect 466 26348 476 26404
rect 532 26348 6188 26404
rect 6244 26348 6254 26404
rect 6402 26348 6412 26404
rect 6468 26348 7756 26404
rect 7812 26348 7822 26404
rect 12450 26348 12460 26404
rect 12516 26348 16884 26404
rect 17042 26348 17052 26404
rect 17108 26348 18396 26404
rect 18452 26348 18462 26404
rect 16828 26292 16884 26348
rect 28448 26292 28560 26320
rect 1922 26236 1932 26292
rect 1988 26236 9884 26292
rect 9940 26236 10892 26292
rect 10948 26236 10958 26292
rect 14578 26236 14588 26292
rect 14644 26236 15260 26292
rect 15316 26236 15326 26292
rect 16828 26236 25228 26292
rect 25284 26236 25294 26292
rect 25666 26236 25676 26292
rect 25732 26236 28560 26292
rect 28448 26208 28560 26236
rect 6178 26124 6188 26180
rect 6244 26124 10220 26180
rect 10276 26124 11676 26180
rect 11732 26124 11742 26180
rect 15810 26124 15820 26180
rect 15876 26124 24332 26180
rect 24388 26124 24398 26180
rect 25218 26124 25228 26180
rect 25284 26124 26236 26180
rect 26292 26124 26302 26180
rect 6710 26012 6748 26068
rect 6804 26012 6814 26068
rect 7410 26012 7420 26068
rect 7476 26012 7980 26068
rect 8036 26012 8046 26068
rect 9874 26012 9884 26068
rect 9940 26012 10108 26068
rect 10164 26012 10174 26068
rect 14578 26012 14588 26068
rect 14644 26012 16828 26068
rect 16884 26012 16894 26068
rect 17378 26012 17388 26068
rect 17444 26012 18284 26068
rect 18340 26012 18350 26068
rect 21298 26012 21308 26068
rect 21364 26012 21868 26068
rect 21924 26012 21934 26068
rect 13794 25900 13804 25956
rect 13860 25900 14252 25956
rect 14308 25900 14318 25956
rect 15922 25900 15932 25956
rect 15988 25900 20524 25956
rect 20580 25900 21084 25956
rect 21140 25900 21150 25956
rect 4454 25844 4464 25900
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4728 25844 4738 25900
rect 24454 25844 24464 25900
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24728 25844 24738 25900
rect 28448 25844 28560 25872
rect 2258 25788 2268 25844
rect 2324 25788 3052 25844
rect 3108 25788 3118 25844
rect 6860 25788 13244 25844
rect 13300 25788 13310 25844
rect 27234 25788 27244 25844
rect 27300 25788 28560 25844
rect 6860 25732 6916 25788
rect 28448 25760 28560 25788
rect 3602 25676 3612 25732
rect 3668 25676 4956 25732
rect 5012 25676 5022 25732
rect 5730 25676 5740 25732
rect 5796 25676 6860 25732
rect 6916 25676 6926 25732
rect 12674 25676 12684 25732
rect 12740 25676 13132 25732
rect 13188 25676 14924 25732
rect 14980 25676 14990 25732
rect 15092 25676 17276 25732
rect 17332 25676 18732 25732
rect 18788 25676 18798 25732
rect 18946 25676 18956 25732
rect 19012 25676 26236 25732
rect 26292 25676 26302 25732
rect 0 25620 112 25648
rect 15092 25620 15148 25676
rect 0 25564 5516 25620
rect 5572 25564 5582 25620
rect 11442 25564 11452 25620
rect 11508 25564 15148 25620
rect 17490 25564 17500 25620
rect 17556 25564 21812 25620
rect 27122 25564 27132 25620
rect 27188 25564 27804 25620
rect 27860 25564 27870 25620
rect 0 25536 112 25564
rect 1810 25452 1820 25508
rect 1876 25452 5572 25508
rect 5730 25452 5740 25508
rect 5796 25452 8652 25508
rect 8708 25452 9996 25508
rect 10052 25452 10062 25508
rect 10210 25452 10220 25508
rect 10276 25452 10668 25508
rect 10724 25452 10734 25508
rect 12898 25452 12908 25508
rect 12964 25452 13132 25508
rect 13188 25452 13198 25508
rect 5516 25396 5572 25452
rect 3378 25340 3388 25396
rect 3444 25340 4228 25396
rect 5516 25340 8988 25396
rect 9044 25340 10556 25396
rect 10612 25340 10622 25396
rect 13234 25340 13244 25396
rect 13300 25340 14476 25396
rect 14532 25340 14542 25396
rect 18386 25340 18396 25396
rect 18452 25340 19740 25396
rect 19796 25340 20524 25396
rect 20580 25340 20590 25396
rect 20738 25340 20748 25396
rect 20804 25340 21308 25396
rect 21364 25340 21374 25396
rect 4172 25172 4228 25340
rect 21756 25284 21812 25564
rect 28448 25396 28560 25424
rect 27122 25340 27132 25396
rect 27188 25340 28560 25396
rect 28448 25312 28560 25340
rect 6178 25228 6188 25284
rect 6244 25228 7084 25284
rect 7140 25228 8876 25284
rect 8932 25228 8942 25284
rect 20178 25228 20188 25284
rect 20244 25228 21420 25284
rect 21476 25228 21486 25284
rect 21746 25228 21756 25284
rect 21812 25228 21822 25284
rect 4162 25116 4172 25172
rect 4228 25116 5852 25172
rect 5908 25116 7756 25172
rect 7812 25116 7822 25172
rect 11442 25116 11452 25172
rect 11508 25116 13692 25172
rect 13748 25116 13758 25172
rect 15586 25116 15596 25172
rect 15652 25116 15876 25172
rect 3794 25060 3804 25116
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 4068 25060 4078 25116
rect 15820 25060 15876 25116
rect 23794 25060 23804 25116
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 24068 25060 24078 25116
rect 5366 25004 5404 25060
rect 5460 25004 5470 25060
rect 8978 25004 8988 25060
rect 9044 25004 9660 25060
rect 9716 25004 12012 25060
rect 12068 25004 12078 25060
rect 15810 25004 15820 25060
rect 15876 25004 15886 25060
rect 28448 24948 28560 24976
rect 1362 24892 1372 24948
rect 1428 24892 9324 24948
rect 9380 24892 9390 24948
rect 13654 24892 13692 24948
rect 13748 24892 13758 24948
rect 25666 24892 25676 24948
rect 25732 24892 28560 24948
rect 28448 24864 28560 24892
rect 2594 24780 2604 24836
rect 2660 24780 6972 24836
rect 7028 24780 7038 24836
rect 7196 24780 26236 24836
rect 26292 24780 26302 24836
rect 0 24724 112 24752
rect 7196 24724 7252 24780
rect 0 24668 3724 24724
rect 3780 24668 3790 24724
rect 5282 24668 5292 24724
rect 5348 24668 7252 24724
rect 8194 24668 8204 24724
rect 8260 24668 8428 24724
rect 8484 24668 8494 24724
rect 10098 24668 10108 24724
rect 10164 24668 10556 24724
rect 10612 24668 10622 24724
rect 13570 24668 13580 24724
rect 13636 24668 14140 24724
rect 14196 24668 15372 24724
rect 15428 24668 15438 24724
rect 0 24640 112 24668
rect 2342 24556 2380 24612
rect 2436 24556 2446 24612
rect 4610 24556 4620 24612
rect 4676 24556 9212 24612
rect 9268 24556 9278 24612
rect 23090 24556 23100 24612
rect 23156 24556 27356 24612
rect 27412 24556 27422 24612
rect 28448 24500 28560 24528
rect 7970 24444 7980 24500
rect 8036 24444 8316 24500
rect 8372 24444 8382 24500
rect 14354 24444 14364 24500
rect 14420 24444 15540 24500
rect 16034 24444 16044 24500
rect 16100 24444 24668 24500
rect 24724 24444 24734 24500
rect 27234 24444 27244 24500
rect 27300 24444 28560 24500
rect 15484 24388 15540 24444
rect 28448 24416 28560 24444
rect 2370 24332 2380 24388
rect 2436 24332 4172 24388
rect 4228 24332 4238 24388
rect 6962 24332 6972 24388
rect 7028 24332 15260 24388
rect 15316 24332 15326 24388
rect 15484 24332 17388 24388
rect 17444 24332 17454 24388
rect 4454 24276 4464 24332
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4728 24276 4738 24332
rect 24454 24276 24464 24332
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24728 24276 24738 24332
rect 9202 24220 9212 24276
rect 9268 24220 17500 24276
rect 17556 24220 17566 24276
rect 1586 24108 1596 24164
rect 1652 24108 6748 24164
rect 6804 24108 6814 24164
rect 12226 24108 12236 24164
rect 12292 24108 12796 24164
rect 12852 24108 12862 24164
rect 15586 24108 15596 24164
rect 15652 24108 16828 24164
rect 16884 24108 16894 24164
rect 21074 24108 21084 24164
rect 21140 24108 22092 24164
rect 22148 24108 22158 24164
rect 6524 24052 6580 24108
rect 28448 24052 28560 24080
rect 3490 23996 3500 24052
rect 3556 23996 3724 24052
rect 3780 23996 3790 24052
rect 5842 23996 5852 24052
rect 5908 23996 6300 24052
rect 6356 23996 6366 24052
rect 6514 23996 6524 24052
rect 6580 23996 6590 24052
rect 10182 23996 10220 24052
rect 10276 23996 10286 24052
rect 17154 23996 17164 24052
rect 17220 23996 19068 24052
rect 19124 23996 20972 24052
rect 21028 23996 22540 24052
rect 22596 23996 22606 24052
rect 25554 23996 25564 24052
rect 25620 23996 28560 24052
rect 28448 23968 28560 23996
rect 690 23884 700 23940
rect 756 23884 2380 23940
rect 2436 23884 2446 23940
rect 5506 23884 5516 23940
rect 5572 23884 7196 23940
rect 7252 23884 7262 23940
rect 12562 23884 12572 23940
rect 12628 23884 13468 23940
rect 13524 23884 13534 23940
rect 18946 23884 18956 23940
rect 19012 23884 19404 23940
rect 19460 23884 19470 23940
rect 20626 23884 20636 23940
rect 20692 23884 26236 23940
rect 26292 23884 26302 23940
rect 0 23828 112 23856
rect 0 23772 1036 23828
rect 1092 23772 1102 23828
rect 1922 23772 1932 23828
rect 1988 23772 3164 23828
rect 3220 23772 3230 23828
rect 10210 23772 10220 23828
rect 10276 23772 11004 23828
rect 11060 23772 11228 23828
rect 11284 23772 11294 23828
rect 16706 23772 16716 23828
rect 16772 23772 26124 23828
rect 26180 23772 26190 23828
rect 0 23744 112 23772
rect 4162 23660 4172 23716
rect 4228 23660 13804 23716
rect 13860 23660 13870 23716
rect 15138 23660 15148 23716
rect 15204 23660 15372 23716
rect 15428 23660 15438 23716
rect 17490 23660 17500 23716
rect 17556 23660 18284 23716
rect 18340 23660 28028 23716
rect 28084 23660 28094 23716
rect 28448 23604 28560 23632
rect 1586 23548 1596 23604
rect 1652 23548 3388 23604
rect 3444 23548 3454 23604
rect 4610 23548 4620 23604
rect 4676 23548 5292 23604
rect 5348 23548 5684 23604
rect 11778 23548 11788 23604
rect 11844 23548 16268 23604
rect 16324 23548 16334 23604
rect 27122 23548 27132 23604
rect 27188 23548 28560 23604
rect 3794 23492 3804 23548
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 4068 23492 4078 23548
rect 5628 23380 5684 23548
rect 23794 23492 23804 23548
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 24068 23492 24078 23548
rect 28448 23520 28560 23548
rect 10098 23436 10108 23492
rect 10164 23436 20188 23492
rect 20244 23436 23548 23492
rect 23604 23436 23614 23492
rect 5618 23324 5628 23380
rect 5684 23324 5694 23380
rect 13458 23324 13468 23380
rect 13524 23324 13692 23380
rect 13748 23324 13758 23380
rect 15092 23324 15148 23436
rect 15204 23324 15214 23380
rect 16258 23324 16268 23380
rect 16324 23324 17052 23380
rect 17108 23324 17118 23380
rect 1474 23212 1484 23268
rect 1540 23212 2268 23268
rect 2324 23212 2334 23268
rect 7074 23212 7084 23268
rect 7140 23212 7756 23268
rect 7812 23212 7822 23268
rect 9650 23212 9660 23268
rect 9716 23212 24892 23268
rect 24948 23212 24958 23268
rect 28448 23156 28560 23184
rect 2706 23100 2716 23156
rect 2772 23100 3276 23156
rect 3332 23100 6076 23156
rect 6132 23100 6142 23156
rect 6290 23100 6300 23156
rect 6356 23100 10332 23156
rect 10388 23100 10398 23156
rect 14690 23100 14700 23156
rect 14756 23100 18396 23156
rect 18452 23100 18462 23156
rect 20038 23100 20076 23156
rect 20132 23100 20142 23156
rect 25666 23100 25676 23156
rect 25732 23100 28560 23156
rect 28448 23072 28560 23100
rect 1698 22988 1708 23044
rect 1764 22988 2268 23044
rect 2324 22988 2334 23044
rect 2930 22988 2940 23044
rect 2996 22988 14140 23044
rect 14196 22988 14206 23044
rect 18610 22988 18620 23044
rect 18676 22988 26236 23044
rect 26292 22988 26302 23044
rect 0 22932 112 22960
rect 0 22876 5516 22932
rect 5572 22876 5582 22932
rect 5730 22876 5740 22932
rect 5796 22876 7532 22932
rect 7588 22876 7598 22932
rect 9426 22876 9436 22932
rect 9492 22876 20636 22932
rect 20692 22876 20702 22932
rect 23426 22876 23436 22932
rect 23492 22876 25564 22932
rect 25620 22876 25630 22932
rect 0 22848 112 22876
rect 2034 22764 2044 22820
rect 2100 22764 2604 22820
rect 2660 22764 2670 22820
rect 6850 22764 6860 22820
rect 6916 22764 9324 22820
rect 9380 22764 9548 22820
rect 9604 22764 9614 22820
rect 13346 22764 13356 22820
rect 13412 22764 15148 22820
rect 4454 22708 4464 22764
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4728 22708 4738 22764
rect 15092 22708 15148 22764
rect 24454 22708 24464 22764
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24728 22708 24738 22764
rect 28448 22708 28560 22736
rect 11666 22652 11676 22708
rect 11732 22652 11742 22708
rect 15092 22652 18340 22708
rect 27234 22652 27244 22708
rect 27300 22652 28560 22708
rect 11676 22596 11732 22652
rect 18284 22596 18340 22652
rect 28448 22624 28560 22652
rect 11218 22540 11228 22596
rect 11284 22540 12236 22596
rect 12292 22540 12302 22596
rect 13346 22540 13356 22596
rect 13412 22540 18060 22596
rect 18116 22540 18126 22596
rect 18284 22540 26236 22596
rect 26292 22540 26302 22596
rect 1586 22428 1596 22484
rect 1652 22428 3052 22484
rect 3108 22428 3118 22484
rect 8530 22428 8540 22484
rect 8596 22428 9996 22484
rect 10052 22428 10062 22484
rect 10770 22428 10780 22484
rect 10836 22428 14812 22484
rect 14868 22428 14878 22484
rect 17938 22428 17948 22484
rect 18004 22428 21868 22484
rect 21924 22428 22876 22484
rect 22932 22428 22942 22484
rect 23426 22428 23436 22484
rect 23492 22428 26572 22484
rect 26628 22428 26638 22484
rect 1138 22316 1148 22372
rect 1204 22316 13468 22372
rect 13524 22316 13534 22372
rect 19058 22316 19068 22372
rect 19124 22316 19628 22372
rect 19684 22316 20188 22372
rect 20244 22316 20254 22372
rect 28448 22260 28560 22288
rect 1250 22204 1260 22260
rect 1316 22204 1484 22260
rect 1540 22204 1708 22260
rect 1764 22204 1774 22260
rect 5618 22204 5628 22260
rect 5684 22204 10444 22260
rect 10500 22204 11788 22260
rect 11844 22204 11854 22260
rect 15362 22204 15372 22260
rect 15428 22204 20076 22260
rect 20132 22204 21420 22260
rect 21476 22204 21486 22260
rect 27122 22204 27132 22260
rect 27188 22204 28560 22260
rect 28448 22176 28560 22204
rect 354 22092 364 22148
rect 420 22092 1596 22148
rect 1652 22092 1662 22148
rect 16146 22092 16156 22148
rect 16212 22092 16828 22148
rect 16884 22092 16894 22148
rect 17378 22092 17388 22148
rect 17444 22092 18396 22148
rect 18452 22092 18462 22148
rect 19282 22092 19292 22148
rect 19348 22092 19516 22148
rect 19572 22092 19582 22148
rect 19842 22092 19852 22148
rect 19908 22092 19964 22148
rect 20020 22092 20030 22148
rect 23538 22092 23548 22148
rect 23604 22092 24332 22148
rect 24388 22092 24398 22148
rect 0 22036 112 22064
rect 0 21980 1484 22036
rect 1540 21980 1550 22036
rect 13346 21980 13356 22036
rect 13412 21980 15372 22036
rect 15428 21980 15438 22036
rect 19730 21980 19740 22036
rect 19796 21980 19806 22036
rect 0 21952 112 21980
rect 3794 21924 3804 21980
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 4068 21924 4078 21980
rect 7746 21868 7756 21924
rect 7812 21868 11564 21924
rect 11620 21868 11630 21924
rect 12002 21868 12012 21924
rect 12068 21868 12124 21924
rect 12180 21868 12190 21924
rect 16034 21868 16044 21924
rect 16100 21868 19068 21924
rect 19124 21868 19134 21924
rect 19740 21812 19796 21980
rect 23794 21924 23804 21980
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 24068 21924 24078 21980
rect 28448 21812 28560 21840
rect 2716 21756 3388 21812
rect 4946 21756 4956 21812
rect 5012 21756 15148 21812
rect 17490 21756 17500 21812
rect 17556 21756 18284 21812
rect 18340 21756 18350 21812
rect 19740 21756 21980 21812
rect 22036 21756 22046 21812
rect 22204 21756 25004 21812
rect 25060 21756 25070 21812
rect 25666 21756 25676 21812
rect 25732 21756 28560 21812
rect 2716 21700 2772 21756
rect 3332 21700 3388 21756
rect 15092 21700 15148 21756
rect 22204 21700 22260 21756
rect 28448 21728 28560 21756
rect 2146 21644 2156 21700
rect 2212 21644 2716 21700
rect 2772 21644 2782 21700
rect 3332 21644 5628 21700
rect 5684 21644 5694 21700
rect 15092 21644 22260 21700
rect 23986 21644 23996 21700
rect 24052 21644 25900 21700
rect 25956 21644 25966 21700
rect 2370 21532 2380 21588
rect 2436 21532 4956 21588
rect 5012 21532 5022 21588
rect 6514 21532 6524 21588
rect 6580 21532 6860 21588
rect 6916 21532 6926 21588
rect 10434 21532 10444 21588
rect 10500 21532 10510 21588
rect 12114 21532 12124 21588
rect 12180 21532 14812 21588
rect 14868 21532 14878 21588
rect 17378 21532 17388 21588
rect 17444 21532 19292 21588
rect 19348 21532 19358 21588
rect 19506 21532 19516 21588
rect 19572 21532 21084 21588
rect 21140 21532 21150 21588
rect 23538 21532 23548 21588
rect 23604 21532 26236 21588
rect 26292 21532 26302 21588
rect 10444 21476 10500 21532
rect 5282 21420 5292 21476
rect 5348 21420 8540 21476
rect 8596 21420 9100 21476
rect 9156 21420 9166 21476
rect 10444 21420 10892 21476
rect 10948 21420 10958 21476
rect 14466 21420 14476 21476
rect 14532 21420 27132 21476
rect 27188 21420 27198 21476
rect 28448 21364 28560 21392
rect 9538 21308 9548 21364
rect 9604 21308 10444 21364
rect 10500 21308 10510 21364
rect 10994 21308 11004 21364
rect 11060 21308 17052 21364
rect 17108 21308 17118 21364
rect 19618 21308 19628 21364
rect 19684 21308 20636 21364
rect 20692 21308 20702 21364
rect 21186 21308 21196 21364
rect 21252 21308 25900 21364
rect 25956 21308 25966 21364
rect 27458 21308 27468 21364
rect 27524 21308 28560 21364
rect 28448 21280 28560 21308
rect 5180 21196 8876 21252
rect 8932 21196 9996 21252
rect 10052 21196 11116 21252
rect 11172 21196 11182 21252
rect 16034 21196 16044 21252
rect 16100 21196 17276 21252
rect 17332 21196 18508 21252
rect 18564 21196 19068 21252
rect 19124 21196 20748 21252
rect 20804 21196 20814 21252
rect 21970 21196 21980 21252
rect 22036 21196 22652 21252
rect 22708 21196 22718 21252
rect 0 21140 112 21168
rect 4454 21140 4464 21196
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4728 21140 4738 21196
rect 0 21084 1652 21140
rect 0 21056 112 21084
rect 1596 20804 1652 21084
rect 5180 21028 5236 21196
rect 24454 21140 24464 21196
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24728 21140 24738 21196
rect 5394 21084 5404 21140
rect 5460 21084 8540 21140
rect 8596 21084 12348 21140
rect 12404 21084 12414 21140
rect 15092 21084 19292 21140
rect 19348 21084 19516 21140
rect 19572 21084 19582 21140
rect 19926 21084 19964 21140
rect 20020 21084 20030 21140
rect 15092 21028 15148 21084
rect 3042 20972 3052 21028
rect 3108 20972 5236 21028
rect 5842 20972 5852 21028
rect 5908 20972 10332 21028
rect 10388 20972 15148 21028
rect 15362 20972 15372 21028
rect 15428 20972 15932 21028
rect 15988 20972 15998 21028
rect 17938 20972 17948 21028
rect 18004 20972 18844 21028
rect 18900 20972 18910 21028
rect 19394 20972 19404 21028
rect 19460 20972 20076 21028
rect 20132 20972 20142 21028
rect 28448 20916 28560 20944
rect 1810 20860 1820 20916
rect 1876 20860 3164 20916
rect 3220 20860 3230 20916
rect 4946 20860 4956 20916
rect 5012 20860 6972 20916
rect 7028 20860 7038 20916
rect 7186 20860 7196 20916
rect 7252 20860 8428 20916
rect 8484 20860 8494 20916
rect 10210 20860 10220 20916
rect 10276 20860 10286 20916
rect 26674 20860 26684 20916
rect 26740 20860 27356 20916
rect 27412 20860 27422 20916
rect 27570 20860 27580 20916
rect 27636 20860 28560 20916
rect 1596 20748 6188 20804
rect 6244 20748 6254 20804
rect 7970 20748 7980 20804
rect 8036 20748 8876 20804
rect 8932 20748 8942 20804
rect 354 20636 364 20692
rect 420 20636 2156 20692
rect 2212 20636 2222 20692
rect 4386 20636 4396 20692
rect 4452 20636 6860 20692
rect 6916 20636 6926 20692
rect 2156 20580 2212 20636
rect 2156 20524 5684 20580
rect 5842 20524 5852 20580
rect 5908 20524 6524 20580
rect 6580 20524 6590 20580
rect 5628 20468 5684 20524
rect 10220 20468 10276 20860
rect 28448 20832 28560 20860
rect 14354 20748 14364 20804
rect 14420 20748 14924 20804
rect 14980 20748 14990 20804
rect 15586 20748 15596 20804
rect 15652 20748 16268 20804
rect 16324 20748 16334 20804
rect 21746 20748 21756 20804
rect 21812 20748 22092 20804
rect 22148 20748 22158 20804
rect 25862 20748 25900 20804
rect 25956 20748 25966 20804
rect 26898 20748 26908 20804
rect 26964 20748 27916 20804
rect 27972 20748 27982 20804
rect 16268 20636 25228 20692
rect 25284 20636 25294 20692
rect 16268 20580 16324 20636
rect 16258 20524 16268 20580
rect 16324 20524 16334 20580
rect 25330 20524 25340 20580
rect 25396 20524 28252 20580
rect 28308 20524 28318 20580
rect 28448 20468 28560 20496
rect 5628 20412 11228 20468
rect 11284 20412 11294 20468
rect 12450 20412 12460 20468
rect 12516 20412 20972 20468
rect 21028 20412 21196 20468
rect 21252 20412 21262 20468
rect 26562 20412 26572 20468
rect 26628 20412 28560 20468
rect 3794 20356 3804 20412
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 4068 20356 4078 20412
rect 23794 20356 23804 20412
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 24068 20356 24078 20412
rect 28448 20384 28560 20412
rect 13122 20300 13132 20356
rect 13188 20300 13468 20356
rect 13524 20300 13534 20356
rect 15138 20300 15148 20356
rect 15204 20300 21140 20356
rect 21298 20300 21308 20356
rect 21364 20300 21644 20356
rect 21700 20300 21710 20356
rect 0 20244 112 20272
rect 21084 20244 21140 20300
rect 0 20188 4844 20244
rect 4900 20188 4910 20244
rect 6962 20188 6972 20244
rect 7028 20188 7756 20244
rect 7812 20188 7822 20244
rect 11106 20188 11116 20244
rect 11172 20188 14700 20244
rect 14756 20188 14766 20244
rect 19394 20188 19404 20244
rect 19460 20188 19740 20244
rect 19796 20188 19806 20244
rect 19954 20188 19964 20244
rect 20020 20188 20860 20244
rect 20916 20188 20926 20244
rect 21084 20188 26796 20244
rect 26852 20188 26862 20244
rect 0 20160 112 20188
rect 7522 20076 7532 20132
rect 7588 20076 7868 20132
rect 7924 20076 19572 20132
rect 4274 19964 4284 20020
rect 4340 19964 7308 20020
rect 7364 19964 7374 20020
rect 9996 19964 12796 20020
rect 12852 19964 12862 20020
rect 13094 19964 13132 20020
rect 13188 19964 13198 20020
rect 14130 19964 14140 20020
rect 14196 19964 14924 20020
rect 14980 19964 16492 20020
rect 16548 19964 16558 20020
rect 18694 19964 18732 20020
rect 18788 19964 18798 20020
rect 9996 19908 10052 19964
rect 9986 19852 9996 19908
rect 10052 19852 10062 19908
rect 10882 19852 10892 19908
rect 10948 19852 13692 19908
rect 13748 19852 14028 19908
rect 14084 19852 14094 19908
rect 15026 19852 15036 19908
rect 15092 19852 17612 19908
rect 17668 19852 17678 19908
rect 17826 19852 17836 19908
rect 17892 19852 18620 19908
rect 18676 19852 18686 19908
rect 19516 19796 19572 20076
rect 19852 20076 20188 20132
rect 20244 20076 20254 20132
rect 20962 20076 20972 20132
rect 21028 20076 22204 20132
rect 22260 20076 22270 20132
rect 25554 20076 25564 20132
rect 25620 20076 26908 20132
rect 19852 20020 19908 20076
rect 26852 20020 26908 20076
rect 28448 20020 28560 20048
rect 19842 19964 19852 20020
rect 19908 19964 19918 20020
rect 20066 19964 20076 20020
rect 20132 19964 21308 20020
rect 21364 19964 21374 20020
rect 22754 19964 22764 20020
rect 22820 19964 26012 20020
rect 26068 19964 26078 20020
rect 26852 19964 28560 20020
rect 28448 19936 28560 19964
rect 19730 19852 19740 19908
rect 19796 19852 20860 19908
rect 20916 19852 20926 19908
rect 21074 19852 21084 19908
rect 21140 19852 26908 19908
rect 26964 19852 26974 19908
rect 10210 19740 10220 19796
rect 10276 19740 15148 19796
rect 19516 19740 26012 19796
rect 26068 19740 26078 19796
rect 7410 19628 7420 19684
rect 7476 19628 11004 19684
rect 11060 19628 11070 19684
rect 12674 19628 12684 19684
rect 12740 19628 13356 19684
rect 13412 19628 13422 19684
rect 14018 19628 14028 19684
rect 14084 19628 14924 19684
rect 14980 19628 14990 19684
rect 4454 19572 4464 19628
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4728 19572 4738 19628
rect 2258 19516 2268 19572
rect 2324 19516 3388 19572
rect 3444 19516 3454 19572
rect 9426 19516 9436 19572
rect 9492 19516 9884 19572
rect 9940 19516 9950 19572
rect 12562 19516 12572 19572
rect 12628 19516 12638 19572
rect 0 19348 112 19376
rect 12572 19348 12628 19516
rect 15092 19460 15148 19740
rect 18834 19628 18844 19684
rect 18900 19628 19516 19684
rect 19572 19628 19582 19684
rect 24454 19572 24464 19628
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24728 19572 24738 19628
rect 28448 19572 28560 19600
rect 15810 19516 15820 19572
rect 15876 19516 18620 19572
rect 18676 19516 20412 19572
rect 20468 19516 20478 19572
rect 27346 19516 27356 19572
rect 27412 19516 28560 19572
rect 28448 19488 28560 19516
rect 12786 19404 12796 19460
rect 12852 19404 12862 19460
rect 15092 19404 24220 19460
rect 24276 19404 24286 19460
rect 0 19292 1148 19348
rect 1204 19292 1214 19348
rect 9846 19292 9884 19348
rect 9940 19292 9950 19348
rect 12012 19292 12628 19348
rect 0 19264 112 19292
rect 4610 19180 4620 19236
rect 4676 19180 5404 19236
rect 5460 19180 5470 19236
rect 12012 19124 12068 19292
rect 12796 19124 12852 19404
rect 15922 19292 15932 19348
rect 15988 19292 25900 19348
rect 25956 19292 25966 19348
rect 26450 19292 26460 19348
rect 26516 19292 26908 19348
rect 26964 19292 26974 19348
rect 13234 19180 13244 19236
rect 13300 19180 13580 19236
rect 13636 19180 13646 19236
rect 15474 19180 15484 19236
rect 15540 19180 15820 19236
rect 15876 19180 15886 19236
rect 17378 19180 17388 19236
rect 17444 19180 19852 19236
rect 19908 19180 19918 19236
rect 28448 19124 28560 19152
rect 12002 19068 12012 19124
rect 12068 19068 12078 19124
rect 12450 19068 12460 19124
rect 12516 19068 16044 19124
rect 16100 19068 17780 19124
rect 1586 18956 1596 19012
rect 1652 18956 1662 19012
rect 5730 18956 5740 19012
rect 5796 18956 5806 19012
rect 8194 18956 8204 19012
rect 8260 18956 12908 19012
rect 12964 18956 14476 19012
rect 14532 18956 14542 19012
rect 16146 18956 16156 19012
rect 16212 18956 17164 19012
rect 17220 18956 17230 19012
rect 1596 18900 1652 18956
rect 5740 18900 5796 18956
rect 17724 18900 17780 19068
rect 18844 19068 25340 19124
rect 25396 19068 25406 19124
rect 27570 19068 27580 19124
rect 27636 19068 28560 19124
rect 18844 19012 18900 19068
rect 28448 19040 28560 19068
rect 18498 18956 18508 19012
rect 18564 18956 18900 19012
rect 19170 18956 19180 19012
rect 19236 18956 26908 19012
rect 26964 18956 26974 19012
rect 1596 18844 2380 18900
rect 2436 18844 2446 18900
rect 5058 18844 5068 18900
rect 5124 18844 15876 18900
rect 16034 18844 16044 18900
rect 16100 18844 17500 18900
rect 17556 18844 17566 18900
rect 17724 18844 18844 18900
rect 18900 18844 18910 18900
rect 19282 18844 19292 18900
rect 19348 18844 20076 18900
rect 20132 18844 20142 18900
rect 3794 18788 3804 18844
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 4068 18788 4078 18844
rect 15820 18788 15876 18844
rect 23794 18788 23804 18844
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 24068 18788 24078 18844
rect 1586 18732 1596 18788
rect 1652 18732 3388 18788
rect 3444 18732 3612 18788
rect 3668 18732 3678 18788
rect 6066 18732 6076 18788
rect 6132 18732 8316 18788
rect 8372 18732 8382 18788
rect 12114 18732 12124 18788
rect 12180 18732 13132 18788
rect 13188 18732 13198 18788
rect 15820 18732 21140 18788
rect 21084 18676 21140 18732
rect 28448 18676 28560 18704
rect 802 18620 812 18676
rect 868 18620 878 18676
rect 2146 18620 2156 18676
rect 2212 18620 6300 18676
rect 6356 18620 6366 18676
rect 10434 18620 10444 18676
rect 10500 18620 10780 18676
rect 10836 18620 13356 18676
rect 13412 18620 13422 18676
rect 18162 18620 18172 18676
rect 18228 18620 20860 18676
rect 20916 18620 20926 18676
rect 21084 18620 25900 18676
rect 25956 18620 25966 18676
rect 26852 18620 28560 18676
rect 812 18564 868 18620
rect 812 18508 1092 18564
rect 2258 18508 2268 18564
rect 2324 18508 2828 18564
rect 2884 18508 2894 18564
rect 3042 18508 3052 18564
rect 3108 18508 3836 18564
rect 3892 18508 3902 18564
rect 5058 18508 5068 18564
rect 5124 18508 18620 18564
rect 18676 18508 18686 18564
rect 0 18452 112 18480
rect 1036 18452 1092 18508
rect 26852 18452 26908 18620
rect 28448 18592 28560 18620
rect 0 18396 812 18452
rect 868 18396 878 18452
rect 1036 18396 3388 18452
rect 0 18368 112 18396
rect 3332 18228 3388 18396
rect 5068 18396 19012 18452
rect 21634 18396 21644 18452
rect 21700 18396 22372 18452
rect 22530 18396 22540 18452
rect 22596 18396 22876 18452
rect 22932 18396 23660 18452
rect 23716 18396 23726 18452
rect 26562 18396 26572 18452
rect 26628 18396 26908 18452
rect 5068 18340 5124 18396
rect 18956 18340 19012 18396
rect 22316 18340 22372 18396
rect 5058 18284 5068 18340
rect 5124 18284 5134 18340
rect 5394 18284 5404 18340
rect 5460 18284 5964 18340
rect 6020 18284 6030 18340
rect 8082 18284 8092 18340
rect 8148 18284 8764 18340
rect 8820 18284 9436 18340
rect 9492 18284 9502 18340
rect 10210 18284 10220 18340
rect 10276 18284 10444 18340
rect 10500 18284 10510 18340
rect 12870 18284 12908 18340
rect 12964 18284 12974 18340
rect 13318 18284 13356 18340
rect 13412 18284 13422 18340
rect 17378 18284 17388 18340
rect 17444 18284 18284 18340
rect 18340 18284 18350 18340
rect 18956 18284 21980 18340
rect 22036 18284 22046 18340
rect 22316 18284 22652 18340
rect 22708 18284 22718 18340
rect 26898 18284 26908 18340
rect 26964 18284 27692 18340
rect 27748 18284 27758 18340
rect 28448 18228 28560 18256
rect 3332 18172 6524 18228
rect 6580 18172 11676 18228
rect 11732 18172 11742 18228
rect 18806 18172 18844 18228
rect 18900 18172 18910 18228
rect 19282 18172 19292 18228
rect 19348 18172 20524 18228
rect 20580 18172 20972 18228
rect 21028 18172 21532 18228
rect 21588 18172 21598 18228
rect 27346 18172 27356 18228
rect 27412 18172 28560 18228
rect 28448 18144 28560 18172
rect 19030 18060 19068 18116
rect 19124 18060 19134 18116
rect 20290 18060 20300 18116
rect 20356 18060 21420 18116
rect 21476 18060 21486 18116
rect 4454 18004 4464 18060
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4728 18004 4738 18060
rect 24454 18004 24464 18060
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24728 18004 24738 18060
rect 9874 17948 9884 18004
rect 9940 17948 9950 18004
rect 11106 17948 11116 18004
rect 11172 17948 11452 18004
rect 11508 17948 11518 18004
rect 20636 17948 21644 18004
rect 21700 17948 21710 18004
rect 4274 17836 4284 17892
rect 4340 17836 6524 17892
rect 6580 17836 6590 17892
rect 2706 17724 2716 17780
rect 2772 17724 5068 17780
rect 5124 17724 5134 17780
rect 6066 17724 6076 17780
rect 6132 17724 8876 17780
rect 8932 17724 8942 17780
rect 9884 17668 9940 17948
rect 20636 17892 20692 17948
rect 16818 17836 16828 17892
rect 16884 17836 19516 17892
rect 19572 17836 19582 17892
rect 19954 17836 19964 17892
rect 20020 17836 20692 17892
rect 20972 17836 26908 17892
rect 26964 17836 26974 17892
rect 17490 17724 17500 17780
rect 17556 17724 18844 17780
rect 18900 17724 18910 17780
rect 2930 17612 2940 17668
rect 2996 17612 4284 17668
rect 4340 17612 4350 17668
rect 8194 17612 8204 17668
rect 8260 17612 8652 17668
rect 8708 17612 9212 17668
rect 9268 17612 9278 17668
rect 9884 17612 16716 17668
rect 16772 17612 17276 17668
rect 17332 17612 17342 17668
rect 18498 17612 18508 17668
rect 18564 17612 19292 17668
rect 19348 17612 19358 17668
rect 19506 17612 19516 17668
rect 19572 17612 20636 17668
rect 20692 17612 20702 17668
rect 0 17556 112 17584
rect 20972 17556 21028 17836
rect 28448 17780 28560 17808
rect 23314 17724 23324 17780
rect 23380 17724 24556 17780
rect 24612 17724 24622 17780
rect 25218 17724 25228 17780
rect 25284 17724 26012 17780
rect 26068 17724 26078 17780
rect 26562 17724 26572 17780
rect 26628 17724 28560 17780
rect 28448 17696 28560 17724
rect 21522 17612 21532 17668
rect 21588 17612 22652 17668
rect 22708 17612 22718 17668
rect 0 17500 1036 17556
rect 1092 17500 1102 17556
rect 3938 17500 3948 17556
rect 4004 17500 5964 17556
rect 6020 17500 21028 17556
rect 21970 17500 21980 17556
rect 22036 17500 26908 17556
rect 26964 17500 26974 17556
rect 0 17472 112 17500
rect 1810 17388 1820 17444
rect 1876 17388 7756 17444
rect 7812 17388 7822 17444
rect 9986 17388 9996 17444
rect 10052 17388 10332 17444
rect 10388 17388 11116 17444
rect 11172 17388 11182 17444
rect 11554 17388 11564 17444
rect 11620 17388 16156 17444
rect 16212 17388 16222 17444
rect 18050 17388 18060 17444
rect 18116 17388 18126 17444
rect 18274 17388 18284 17444
rect 18340 17388 19404 17444
rect 19460 17388 22092 17444
rect 22148 17388 22158 17444
rect 18060 17332 18116 17388
rect 28448 17332 28560 17360
rect 5170 17276 5180 17332
rect 5236 17276 5516 17332
rect 5572 17276 5582 17332
rect 9762 17276 9772 17332
rect 9828 17276 14924 17332
rect 14980 17276 14990 17332
rect 15810 17276 15820 17332
rect 15876 17276 16940 17332
rect 16996 17276 20972 17332
rect 21028 17276 21038 17332
rect 27570 17276 27580 17332
rect 27636 17276 28560 17332
rect 3794 17220 3804 17276
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 4068 17220 4078 17276
rect 23794 17220 23804 17276
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 24068 17220 24078 17276
rect 28448 17248 28560 17276
rect 4722 17164 4732 17220
rect 4788 17164 7308 17220
rect 7364 17164 12404 17220
rect 12348 17108 12404 17164
rect 15092 17164 19236 17220
rect 19394 17164 19404 17220
rect 19460 17164 19628 17220
rect 19684 17164 19694 17220
rect 15092 17108 15148 17164
rect 19180 17108 19236 17164
rect 1250 17052 1260 17108
rect 1316 17052 1708 17108
rect 1764 17052 9996 17108
rect 10052 17052 10062 17108
rect 11106 17052 11116 17108
rect 11172 17052 12124 17108
rect 12180 17052 12190 17108
rect 12348 17052 15148 17108
rect 15810 17052 15820 17108
rect 15876 17052 16268 17108
rect 16324 17052 16334 17108
rect 17378 17052 17388 17108
rect 17444 17052 18284 17108
rect 18340 17052 18350 17108
rect 18498 17052 18508 17108
rect 18564 17052 18732 17108
rect 18788 17052 18798 17108
rect 19180 17052 23548 17108
rect 23604 17052 26012 17108
rect 26068 17052 26078 17108
rect 3826 16940 3836 16996
rect 3892 16940 4172 16996
rect 4228 16940 4238 16996
rect 7746 16940 7756 16996
rect 7812 16940 8988 16996
rect 9044 16940 9054 16996
rect 9202 16940 9212 16996
rect 9268 16940 14700 16996
rect 14756 16940 14766 16996
rect 14914 16940 14924 16996
rect 14980 16940 26012 16996
rect 26068 16940 26078 16996
rect 26236 16940 28140 16996
rect 28196 16940 28206 16996
rect 26236 16884 26292 16940
rect 28448 16884 28560 16912
rect 1810 16828 1820 16884
rect 1876 16828 3164 16884
rect 3220 16828 4284 16884
rect 4340 16828 5740 16884
rect 5796 16828 5806 16884
rect 8194 16828 8204 16884
rect 8260 16828 9324 16884
rect 9380 16828 9390 16884
rect 9874 16828 9884 16884
rect 9940 16828 9996 16884
rect 10052 16828 10062 16884
rect 12786 16828 12796 16884
rect 12852 16828 15036 16884
rect 15092 16828 15102 16884
rect 17266 16828 17276 16884
rect 17332 16828 19740 16884
rect 19796 16828 19806 16884
rect 20962 16828 20972 16884
rect 21028 16828 26292 16884
rect 26562 16828 26572 16884
rect 26628 16828 28560 16884
rect 28448 16800 28560 16828
rect 1586 16716 1596 16772
rect 1652 16716 2044 16772
rect 2100 16716 2110 16772
rect 3602 16716 3612 16772
rect 3668 16716 13580 16772
rect 13636 16716 13646 16772
rect 13794 16716 13804 16772
rect 13860 16716 26908 16772
rect 26964 16716 26974 16772
rect 0 16660 112 16688
rect 0 16604 5292 16660
rect 5348 16604 5358 16660
rect 12562 16604 12572 16660
rect 12628 16604 14140 16660
rect 14196 16604 14206 16660
rect 18610 16604 18620 16660
rect 18676 16604 20860 16660
rect 20916 16604 20926 16660
rect 0 16576 112 16604
rect 4918 16492 4956 16548
rect 5012 16492 5022 16548
rect 12114 16492 12124 16548
rect 12180 16492 18732 16548
rect 18788 16492 19068 16548
rect 19124 16492 19134 16548
rect 20626 16492 20636 16548
rect 20692 16492 21308 16548
rect 21364 16492 21374 16548
rect 4454 16436 4464 16492
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4728 16436 4738 16492
rect 24454 16436 24464 16492
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24728 16436 24738 16492
rect 28448 16436 28560 16464
rect 8530 16380 8540 16436
rect 8596 16380 14476 16436
rect 14532 16380 14542 16436
rect 17378 16380 17388 16436
rect 17444 16380 17948 16436
rect 18004 16380 18014 16436
rect 18918 16380 18956 16436
rect 19012 16380 19022 16436
rect 19366 16380 19404 16436
rect 19460 16380 19470 16436
rect 19618 16380 19628 16436
rect 19684 16380 19740 16436
rect 19796 16380 19806 16436
rect 27346 16380 27356 16436
rect 27412 16380 28560 16436
rect 28448 16352 28560 16380
rect 1362 16268 1372 16324
rect 1428 16268 3388 16324
rect 4162 16268 4172 16324
rect 4228 16268 4956 16324
rect 5012 16268 5022 16324
rect 5842 16268 5852 16324
rect 5908 16268 5918 16324
rect 7410 16268 7420 16324
rect 7476 16268 13804 16324
rect 13860 16268 13870 16324
rect 15092 16268 22540 16324
rect 22596 16268 22606 16324
rect 3332 16212 3388 16268
rect 5852 16212 5908 16268
rect 1810 16156 1820 16212
rect 1876 16156 2380 16212
rect 2436 16156 2828 16212
rect 2884 16156 2894 16212
rect 3332 16156 5908 16212
rect 6962 16156 6972 16212
rect 7028 16156 9324 16212
rect 9380 16156 9390 16212
rect 10406 16156 10444 16212
rect 10500 16156 10510 16212
rect 9324 16100 9380 16156
rect 15092 16100 15148 16268
rect 17266 16156 17276 16212
rect 17332 16156 20412 16212
rect 20468 16156 20478 16212
rect 26898 16156 26908 16212
rect 26964 16156 28028 16212
rect 28084 16156 28094 16212
rect 3602 16044 3612 16100
rect 3668 16044 7532 16100
rect 7588 16044 7598 16100
rect 9324 16044 13804 16100
rect 13860 16044 15148 16100
rect 16930 16044 16940 16100
rect 16996 16044 18284 16100
rect 18340 16044 18350 16100
rect 18694 16044 18732 16100
rect 18788 16044 18798 16100
rect 18946 16044 18956 16100
rect 19012 16044 19628 16100
rect 19684 16044 19694 16100
rect 28448 15988 28560 16016
rect 5618 15932 5628 15988
rect 5684 15932 6300 15988
rect 6356 15932 6366 15988
rect 6626 15932 6636 15988
rect 6692 15932 8092 15988
rect 8148 15932 8158 15988
rect 9874 15932 9884 15988
rect 9940 15932 10556 15988
rect 10612 15932 10622 15988
rect 14354 15932 14364 15988
rect 14420 15932 19180 15988
rect 19236 15932 19246 15988
rect 21410 15932 21420 15988
rect 21476 15932 26292 15988
rect 26562 15932 26572 15988
rect 26628 15932 28560 15988
rect 26236 15876 26292 15932
rect 28448 15904 28560 15932
rect 7970 15820 7980 15876
rect 8036 15820 9212 15876
rect 9268 15820 9278 15876
rect 13430 15820 13468 15876
rect 13524 15820 13534 15876
rect 15026 15820 15036 15876
rect 15092 15820 16156 15876
rect 16212 15820 16222 15876
rect 17154 15820 17164 15876
rect 17220 15820 18172 15876
rect 18228 15820 18844 15876
rect 18900 15820 18910 15876
rect 19618 15820 19628 15876
rect 19684 15820 26012 15876
rect 26068 15820 26078 15876
rect 26236 15820 28028 15876
rect 28084 15820 28094 15876
rect 0 15764 112 15792
rect 0 15708 2828 15764
rect 2884 15708 2894 15764
rect 6738 15708 6748 15764
rect 6804 15708 7084 15764
rect 7140 15708 7150 15764
rect 18498 15708 18508 15764
rect 18564 15708 21420 15764
rect 21476 15708 21486 15764
rect 0 15680 112 15708
rect 3794 15652 3804 15708
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 4068 15652 4078 15708
rect 23794 15652 23804 15708
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 24068 15652 24078 15708
rect 17714 15596 17724 15652
rect 17780 15596 20636 15652
rect 20692 15596 20702 15652
rect 28448 15540 28560 15568
rect 4050 15484 4060 15540
rect 4116 15484 5180 15540
rect 5236 15484 8316 15540
rect 8372 15484 10556 15540
rect 10612 15484 12572 15540
rect 12628 15484 12638 15540
rect 14466 15484 14476 15540
rect 14532 15484 26908 15540
rect 26964 15484 26974 15540
rect 27570 15484 27580 15540
rect 27636 15484 28560 15540
rect 28448 15456 28560 15484
rect 3332 15372 3500 15428
rect 3556 15372 5908 15428
rect 7858 15372 7868 15428
rect 7924 15372 19628 15428
rect 19684 15372 19694 15428
rect 19842 15372 19852 15428
rect 19908 15372 20076 15428
rect 20132 15372 20142 15428
rect 20626 15372 20636 15428
rect 20692 15372 26684 15428
rect 26740 15372 26750 15428
rect 3332 15316 3388 15372
rect 5852 15316 5908 15372
rect 1362 15260 1372 15316
rect 1428 15260 1820 15316
rect 1876 15260 1886 15316
rect 2594 15260 2604 15316
rect 2660 15260 3388 15316
rect 3948 15260 5404 15316
rect 5460 15260 5470 15316
rect 5842 15260 5852 15316
rect 5908 15260 7532 15316
rect 7588 15260 8876 15316
rect 8932 15260 8942 15316
rect 12450 15260 12460 15316
rect 12516 15260 15148 15316
rect 15204 15260 15214 15316
rect 16818 15260 16828 15316
rect 16884 15260 18396 15316
rect 18452 15260 18462 15316
rect 19730 15260 19740 15316
rect 19796 15260 20524 15316
rect 20580 15260 20590 15316
rect 21186 15260 21196 15316
rect 21252 15260 22092 15316
rect 22148 15260 22158 15316
rect 22978 15260 22988 15316
rect 23044 15260 27692 15316
rect 27748 15260 27758 15316
rect 1586 15148 1596 15204
rect 1652 15148 2268 15204
rect 2324 15148 2334 15204
rect 3042 15148 3052 15204
rect 3108 15148 3724 15204
rect 3780 15148 3790 15204
rect 3948 15092 4004 15260
rect 6962 15148 6972 15204
rect 7028 15148 7420 15204
rect 7476 15148 7486 15204
rect 7634 15148 7644 15204
rect 7700 15148 9100 15204
rect 9156 15148 9166 15204
rect 9538 15148 9548 15204
rect 9604 15148 10892 15204
rect 10948 15148 10958 15204
rect 14690 15148 14700 15204
rect 14756 15148 16492 15204
rect 16548 15148 17836 15204
rect 17892 15148 17902 15204
rect 20066 15148 20076 15204
rect 20132 15148 21644 15204
rect 21700 15148 21710 15204
rect 26002 15148 26012 15204
rect 26068 15148 26236 15204
rect 26292 15148 26302 15204
rect 28448 15092 28560 15120
rect 2146 15036 2156 15092
rect 2212 15036 2716 15092
rect 2772 15036 4004 15092
rect 7074 15036 7084 15092
rect 7140 15036 7756 15092
rect 7812 15036 7822 15092
rect 17490 15036 17500 15092
rect 17556 15036 18396 15092
rect 18452 15036 18462 15092
rect 21074 15036 21084 15092
rect 21140 15036 23660 15092
rect 23716 15036 23726 15092
rect 26562 15036 26572 15092
rect 26628 15036 28560 15092
rect 28448 15008 28560 15036
rect 7410 14924 7420 14980
rect 7476 14924 8764 14980
rect 8820 14924 8830 14980
rect 17042 14924 17052 14980
rect 17108 14924 17276 14980
rect 17332 14924 20524 14980
rect 20580 14924 21196 14980
rect 21252 14924 21262 14980
rect 0 14868 112 14896
rect 4454 14868 4464 14924
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4728 14868 4738 14924
rect 24454 14868 24464 14924
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24728 14868 24738 14924
rect 0 14812 3332 14868
rect 6178 14812 6188 14868
rect 6244 14812 9324 14868
rect 9380 14812 9390 14868
rect 15362 14812 15372 14868
rect 15428 14812 19852 14868
rect 19908 14812 19918 14868
rect 0 14784 112 14812
rect 3276 14644 3332 14812
rect 4162 14700 4172 14756
rect 4228 14700 8540 14756
rect 8596 14700 8606 14756
rect 9202 14700 9212 14756
rect 9268 14700 26908 14756
rect 3276 14588 6412 14644
rect 6468 14588 6478 14644
rect 6850 14588 6860 14644
rect 6916 14588 7756 14644
rect 7812 14588 8876 14644
rect 8932 14588 8942 14644
rect 14690 14588 14700 14644
rect 14756 14588 17052 14644
rect 17108 14588 18620 14644
rect 18676 14588 19292 14644
rect 19348 14588 19358 14644
rect 19730 14588 19740 14644
rect 19796 14588 19852 14644
rect 19908 14588 22764 14644
rect 22820 14588 22830 14644
rect 26852 14532 26908 14700
rect 28448 14644 28560 14672
rect 27346 14588 27356 14644
rect 27412 14588 28560 14644
rect 28448 14560 28560 14588
rect 4274 14476 4284 14532
rect 4340 14476 7308 14532
rect 7364 14476 8036 14532
rect 8194 14476 8204 14532
rect 8260 14476 8764 14532
rect 8820 14476 8830 14532
rect 12002 14476 12012 14532
rect 12068 14476 12460 14532
rect 12516 14476 12526 14532
rect 16706 14476 16716 14532
rect 16772 14476 18060 14532
rect 18116 14476 19180 14532
rect 19236 14476 19246 14532
rect 20738 14476 20748 14532
rect 20804 14476 21084 14532
rect 21140 14476 21150 14532
rect 25666 14476 25676 14532
rect 25732 14476 26348 14532
rect 26404 14476 26414 14532
rect 26852 14476 27020 14532
rect 27076 14476 27086 14532
rect 7980 14308 8036 14476
rect 20748 14420 20804 14476
rect 8306 14364 8316 14420
rect 8372 14364 8428 14420
rect 8484 14364 8494 14420
rect 13122 14364 13132 14420
rect 13188 14364 14364 14420
rect 14420 14364 14430 14420
rect 16818 14364 16828 14420
rect 16884 14364 20804 14420
rect 4722 14252 4732 14308
rect 4788 14252 7308 14308
rect 7364 14252 7374 14308
rect 7980 14252 8204 14308
rect 8260 14252 8270 14308
rect 17938 14252 17948 14308
rect 18004 14252 18396 14308
rect 18452 14252 20076 14308
rect 20132 14252 20972 14308
rect 21028 14252 21420 14308
rect 21476 14252 21486 14308
rect 21858 14252 21868 14308
rect 21924 14252 26348 14308
rect 26404 14252 26414 14308
rect 28448 14196 28560 14224
rect 4386 14140 4396 14196
rect 4452 14140 9212 14196
rect 9268 14140 9278 14196
rect 12002 14140 12012 14196
rect 12068 14140 15372 14196
rect 15428 14140 15438 14196
rect 15586 14140 15596 14196
rect 15652 14140 22204 14196
rect 22260 14140 22270 14196
rect 27458 14140 27468 14196
rect 27524 14140 28560 14196
rect 3794 14084 3804 14140
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 4068 14084 4078 14140
rect 23794 14084 23804 14140
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 24068 14084 24078 14140
rect 28448 14112 28560 14140
rect 4620 14028 9940 14084
rect 17154 14028 17164 14084
rect 17220 14028 19068 14084
rect 19124 14028 19134 14084
rect 0 13972 112 14000
rect 4620 13972 4676 14028
rect 0 13916 1372 13972
rect 1428 13916 1438 13972
rect 3714 13916 3724 13972
rect 3780 13916 4676 13972
rect 4834 13916 4844 13972
rect 4900 13916 5516 13972
rect 5572 13916 5582 13972
rect 0 13888 112 13916
rect 9884 13860 9940 14028
rect 14690 13916 14700 13972
rect 14756 13916 15148 13972
rect 15204 13916 15214 13972
rect 16594 13916 16604 13972
rect 16660 13916 17388 13972
rect 17444 13916 17454 13972
rect 19282 13916 19292 13972
rect 19348 13916 19964 13972
rect 20020 13916 20030 13972
rect 3938 13804 3948 13860
rect 4004 13804 4956 13860
rect 5012 13804 8372 13860
rect 8530 13804 8540 13860
rect 8596 13804 9324 13860
rect 9380 13804 9390 13860
rect 9884 13804 19740 13860
rect 19796 13804 19806 13860
rect 22754 13804 22764 13860
rect 22820 13804 25508 13860
rect 27010 13804 27020 13860
rect 27076 13804 27132 13860
rect 27188 13804 27198 13860
rect 8316 13748 8372 13804
rect 1698 13692 1708 13748
rect 1764 13692 8092 13748
rect 8148 13692 8158 13748
rect 8316 13692 15260 13748
rect 15316 13692 15326 13748
rect 20850 13692 20860 13748
rect 20916 13692 21420 13748
rect 21476 13692 21644 13748
rect 21700 13692 21710 13748
rect 24210 13692 24220 13748
rect 24276 13692 24892 13748
rect 24948 13692 25228 13748
rect 25284 13692 25294 13748
rect 25452 13636 25508 13804
rect 28448 13748 28560 13776
rect 26562 13692 26572 13748
rect 26628 13692 28560 13748
rect 28448 13664 28560 13692
rect 3378 13580 3388 13636
rect 3444 13580 4956 13636
rect 5012 13580 5022 13636
rect 7410 13580 7420 13636
rect 7476 13580 10220 13636
rect 10276 13580 11340 13636
rect 11396 13580 11406 13636
rect 13794 13580 13804 13636
rect 13860 13580 15148 13636
rect 15204 13580 15214 13636
rect 19954 13580 19964 13636
rect 20020 13580 20972 13636
rect 21028 13580 21038 13636
rect 21746 13580 21756 13636
rect 21812 13580 24332 13636
rect 24388 13580 24398 13636
rect 25452 13580 26628 13636
rect 26572 13524 26628 13580
rect 2258 13468 2268 13524
rect 2324 13468 4844 13524
rect 4900 13468 4910 13524
rect 6402 13468 6412 13524
rect 6468 13468 7196 13524
rect 7252 13468 7262 13524
rect 8530 13468 8540 13524
rect 8596 13468 8820 13524
rect 10434 13468 10444 13524
rect 10500 13468 12572 13524
rect 12628 13468 12638 13524
rect 12786 13468 12796 13524
rect 12852 13468 12890 13524
rect 14018 13468 14028 13524
rect 14084 13468 14364 13524
rect 14420 13468 14812 13524
rect 14868 13468 14878 13524
rect 19730 13468 19740 13524
rect 19796 13468 20748 13524
rect 20804 13468 20814 13524
rect 23762 13468 23772 13524
rect 23828 13468 25228 13524
rect 25284 13468 25294 13524
rect 26562 13468 26572 13524
rect 26628 13468 26638 13524
rect 8764 13412 8820 13468
rect 8754 13356 8764 13412
rect 8820 13356 8830 13412
rect 11638 13356 11676 13412
rect 11732 13356 11742 13412
rect 12674 13356 12684 13412
rect 12740 13356 12908 13412
rect 12964 13356 12974 13412
rect 13234 13356 13244 13412
rect 13300 13356 13356 13412
rect 13412 13356 13422 13412
rect 20514 13356 20524 13412
rect 20580 13356 20860 13412
rect 20916 13356 20926 13412
rect 4454 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4738 13356
rect 24454 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24738 13356
rect 28448 13300 28560 13328
rect 1810 13244 1820 13300
rect 1876 13244 2268 13300
rect 2324 13244 2334 13300
rect 5730 13244 5740 13300
rect 5796 13244 19516 13300
rect 19572 13244 19582 13300
rect 21074 13244 21084 13300
rect 21140 13244 21420 13300
rect 21476 13244 21486 13300
rect 27346 13244 27356 13300
rect 27412 13244 28560 13300
rect 28448 13216 28560 13244
rect 578 13132 588 13188
rect 644 13132 3164 13188
rect 3220 13132 3230 13188
rect 7186 13132 7196 13188
rect 7252 13132 7644 13188
rect 7700 13132 8092 13188
rect 8148 13132 8158 13188
rect 8278 13132 8316 13188
rect 8372 13132 8382 13188
rect 12684 13132 22540 13188
rect 22596 13132 23324 13188
rect 23380 13132 23390 13188
rect 0 13076 112 13104
rect 12684 13076 12740 13132
rect 0 13020 3052 13076
rect 3108 13020 3118 13076
rect 8418 13020 8428 13076
rect 8484 13020 9996 13076
rect 10052 13020 10062 13076
rect 11666 13020 11676 13076
rect 11732 13020 12684 13076
rect 12740 13020 12750 13076
rect 17798 13020 17836 13076
rect 17892 13020 18284 13076
rect 18340 13020 18350 13076
rect 19142 13020 19180 13076
rect 19236 13020 19246 13076
rect 0 12992 112 13020
rect 2370 12908 2380 12964
rect 2436 12908 15596 12964
rect 15652 12908 15662 12964
rect 16034 12908 16044 12964
rect 16100 12908 17388 12964
rect 17444 12908 18396 12964
rect 18452 12908 18462 12964
rect 19842 12908 19852 12964
rect 19908 12908 21420 12964
rect 21476 12908 27468 12964
rect 27524 12908 27534 12964
rect 28448 12852 28560 12880
rect 3332 12796 9604 12852
rect 9986 12796 9996 12852
rect 10052 12796 12572 12852
rect 12628 12796 13020 12852
rect 13076 12796 13086 12852
rect 18022 12796 18060 12852
rect 18116 12796 18126 12852
rect 19618 12796 19628 12852
rect 19684 12796 20076 12852
rect 20132 12796 20412 12852
rect 20468 12796 20478 12852
rect 26562 12796 26572 12852
rect 26628 12796 28560 12852
rect 3332 12740 3388 12796
rect 9548 12740 9604 12796
rect 28448 12768 28560 12796
rect 2594 12684 2604 12740
rect 2660 12684 3388 12740
rect 8194 12684 8204 12740
rect 8260 12684 9324 12740
rect 9380 12684 9390 12740
rect 9548 12684 13916 12740
rect 13972 12684 13982 12740
rect 17126 12684 17164 12740
rect 17220 12684 17724 12740
rect 17780 12684 17790 12740
rect 17938 12684 17948 12740
rect 18004 12684 24220 12740
rect 24276 12684 24286 12740
rect 7410 12572 7420 12628
rect 7476 12572 23660 12628
rect 23716 12572 23726 12628
rect 27122 12572 27132 12628
rect 27188 12572 28028 12628
rect 28084 12572 28094 12628
rect 3794 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4078 12572
rect 23794 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24078 12572
rect 4162 12460 4172 12516
rect 4228 12460 4956 12516
rect 5012 12460 7924 12516
rect 9426 12460 9436 12516
rect 9492 12460 9660 12516
rect 9716 12460 9726 12516
rect 10322 12460 10332 12516
rect 10388 12460 10780 12516
rect 10836 12460 10846 12516
rect 11974 12460 12012 12516
rect 12068 12460 12078 12516
rect 12758 12460 12796 12516
rect 12852 12460 12862 12516
rect 13682 12460 13692 12516
rect 13748 12460 18228 12516
rect 20514 12460 20524 12516
rect 20580 12460 20860 12516
rect 20916 12460 21532 12516
rect 21588 12460 21598 12516
rect 7868 12404 7924 12460
rect 18172 12404 18228 12460
rect 28448 12404 28560 12432
rect 3602 12348 3612 12404
rect 3668 12348 5068 12404
rect 5124 12348 5134 12404
rect 6962 12348 6972 12404
rect 7028 12348 7038 12404
rect 7868 12348 14924 12404
rect 14980 12348 14990 12404
rect 15092 12348 17948 12404
rect 18004 12348 18014 12404
rect 18172 12348 26012 12404
rect 26068 12348 26078 12404
rect 27570 12348 27580 12404
rect 27636 12348 28560 12404
rect 6972 12292 7028 12348
rect 15092 12292 15148 12348
rect 28448 12320 28560 12348
rect 2482 12236 2492 12292
rect 2548 12236 5628 12292
rect 5684 12236 5694 12292
rect 6972 12236 9436 12292
rect 9492 12236 12236 12292
rect 12292 12236 12302 12292
rect 12450 12236 12460 12292
rect 12516 12236 15148 12292
rect 16146 12236 16156 12292
rect 16212 12236 17612 12292
rect 17668 12236 19628 12292
rect 19684 12236 19694 12292
rect 27458 12236 27468 12292
rect 27524 12236 28028 12292
rect 28084 12236 28094 12292
rect 0 12180 112 12208
rect 0 12124 1148 12180
rect 1204 12124 1214 12180
rect 2034 12124 2044 12180
rect 2100 12124 2268 12180
rect 2324 12124 3164 12180
rect 3220 12124 6412 12180
rect 6468 12124 6478 12180
rect 9062 12124 9100 12180
rect 9156 12124 15148 12180
rect 16482 12124 16492 12180
rect 16548 12124 18508 12180
rect 18564 12124 19964 12180
rect 20020 12124 20030 12180
rect 25974 12124 26012 12180
rect 26068 12124 26078 12180
rect 0 12096 112 12124
rect 15092 12068 15148 12124
rect 4162 12012 4172 12068
rect 4228 12012 6748 12068
rect 6804 12012 6814 12068
rect 8306 12012 8316 12068
rect 8372 12012 8382 12068
rect 8530 12012 8540 12068
rect 8596 12012 8988 12068
rect 9044 12012 9054 12068
rect 15092 12012 26908 12068
rect 26964 12012 26974 12068
rect 8316 11956 8372 12012
rect 28448 11956 28560 11984
rect 3602 11900 3612 11956
rect 3668 11900 5404 11956
rect 5460 11900 5470 11956
rect 7298 11900 7308 11956
rect 7364 11900 8764 11956
rect 8820 11900 12460 11956
rect 12516 11900 12526 11956
rect 17042 11900 17052 11956
rect 17108 11900 18844 11956
rect 18900 11900 18910 11956
rect 19478 11900 19516 11956
rect 19572 11900 19582 11956
rect 19730 11900 19740 11956
rect 19796 11900 21084 11956
rect 21140 11900 21150 11956
rect 21410 11900 21420 11956
rect 21476 11900 25900 11956
rect 25956 11900 25966 11956
rect 26562 11900 26572 11956
rect 26628 11900 28560 11956
rect 4454 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4738 11788
rect 7308 11732 7364 11900
rect 28448 11872 28560 11900
rect 8306 11788 8316 11844
rect 8372 11788 8652 11844
rect 8708 11788 8718 11844
rect 9314 11788 9324 11844
rect 9380 11788 9772 11844
rect 9828 11788 9838 11844
rect 17798 11788 17836 11844
rect 17892 11788 17902 11844
rect 18022 11788 18060 11844
rect 18116 11788 18126 11844
rect 19170 11788 19180 11844
rect 19236 11788 19292 11844
rect 19348 11788 19358 11844
rect 20178 11788 20188 11844
rect 20244 11788 20636 11844
rect 20692 11788 20702 11844
rect 22642 11788 22652 11844
rect 22708 11788 23212 11844
rect 23268 11788 23660 11844
rect 23716 11788 23726 11844
rect 24454 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24738 11788
rect 6514 11676 6524 11732
rect 6580 11676 7364 11732
rect 11106 11676 11116 11732
rect 11172 11676 11452 11732
rect 11508 11676 13356 11732
rect 13412 11676 13422 11732
rect 15092 11676 21868 11732
rect 21924 11676 21934 11732
rect 25330 11676 25340 11732
rect 25396 11676 25900 11732
rect 25956 11676 25966 11732
rect 15092 11620 15148 11676
rect 1586 11564 1596 11620
rect 1652 11564 1932 11620
rect 1988 11564 1998 11620
rect 2370 11564 2380 11620
rect 2436 11564 15148 11620
rect 15586 11564 15596 11620
rect 15652 11564 15662 11620
rect 16370 11564 16380 11620
rect 16436 11564 26012 11620
rect 26068 11564 26078 11620
rect 15596 11508 15652 11564
rect 28448 11508 28560 11536
rect 2706 11452 2716 11508
rect 2772 11452 5404 11508
rect 5460 11452 5852 11508
rect 5908 11452 5918 11508
rect 6626 11452 6636 11508
rect 6692 11452 6972 11508
rect 7028 11452 8204 11508
rect 8260 11452 9212 11508
rect 9268 11452 9278 11508
rect 9874 11452 9884 11508
rect 9940 11452 15652 11508
rect 17154 11452 17164 11508
rect 17220 11452 18396 11508
rect 18452 11452 19180 11508
rect 19236 11452 19246 11508
rect 20850 11452 20860 11508
rect 20916 11452 22204 11508
rect 22260 11452 22270 11508
rect 23762 11452 23772 11508
rect 23828 11452 25452 11508
rect 25508 11452 25518 11508
rect 26870 11452 26908 11508
rect 26964 11452 26974 11508
rect 27346 11452 27356 11508
rect 27412 11452 28560 11508
rect 15596 11396 15652 11452
rect 28448 11424 28560 11452
rect 11666 11340 11676 11396
rect 11732 11340 11742 11396
rect 15596 11340 17220 11396
rect 18498 11340 18508 11396
rect 18564 11340 20076 11396
rect 20132 11340 25340 11396
rect 25396 11340 25406 11396
rect 0 11284 112 11312
rect 11676 11284 11732 11340
rect 17164 11284 17220 11340
rect 0 11228 3276 11284
rect 3332 11228 3342 11284
rect 8306 11228 8316 11284
rect 8372 11228 16828 11284
rect 16884 11228 16894 11284
rect 17154 11228 17164 11284
rect 17220 11228 26236 11284
rect 26292 11228 26302 11284
rect 0 11200 112 11228
rect 4274 11116 4284 11172
rect 4340 11116 10780 11172
rect 10836 11116 10846 11172
rect 11638 11116 11676 11172
rect 11732 11116 11742 11172
rect 13010 11116 13020 11172
rect 13076 11116 13244 11172
rect 13300 11116 19404 11172
rect 19460 11116 25004 11172
rect 25060 11116 25070 11172
rect 28448 11060 28560 11088
rect 9062 11004 9100 11060
rect 9156 11004 9166 11060
rect 11106 11004 11116 11060
rect 11172 11004 11340 11060
rect 11396 11004 11406 11060
rect 11778 11004 11788 11060
rect 11844 11004 12012 11060
rect 12068 11004 12078 11060
rect 17938 11004 17948 11060
rect 18004 11004 18508 11060
rect 18564 11004 18574 11060
rect 26562 11004 26572 11060
rect 26628 11004 28560 11060
rect 3794 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4078 11004
rect 23794 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24078 11004
rect 28448 10976 28560 11004
rect 7186 10892 7196 10948
rect 7252 10892 8092 10948
rect 8148 10892 8158 10948
rect 8754 10892 8764 10948
rect 8820 10892 9212 10948
rect 9268 10892 9278 10948
rect 10882 10892 10892 10948
rect 10948 10892 11564 10948
rect 11620 10892 11630 10948
rect 26898 10892 26908 10948
rect 26964 10892 27692 10948
rect 27748 10892 27758 10948
rect 4946 10780 4956 10836
rect 5012 10780 5180 10836
rect 5236 10780 8820 10836
rect 12114 10780 12124 10836
rect 12180 10780 12796 10836
rect 12852 10780 12862 10836
rect 17266 10780 17276 10836
rect 17332 10780 18284 10836
rect 18340 10780 19964 10836
rect 20020 10780 20030 10836
rect 8764 10724 8820 10780
rect 1922 10668 1932 10724
rect 1988 10668 7980 10724
rect 8036 10668 8046 10724
rect 8726 10668 8764 10724
rect 8820 10668 8830 10724
rect 10658 10668 10668 10724
rect 10724 10668 10948 10724
rect 11106 10668 11116 10724
rect 11172 10668 13244 10724
rect 13300 10668 13310 10724
rect 17714 10668 17724 10724
rect 17780 10668 18620 10724
rect 18676 10668 18686 10724
rect 7858 10556 7868 10612
rect 7924 10556 9436 10612
rect 9492 10556 9502 10612
rect 2034 10444 2044 10500
rect 2100 10444 6524 10500
rect 6580 10444 6590 10500
rect 6738 10444 6748 10500
rect 6804 10444 7756 10500
rect 7812 10444 9660 10500
rect 9716 10444 9726 10500
rect 0 10388 112 10416
rect 10892 10388 10948 10668
rect 28448 10612 28560 10640
rect 12226 10556 12236 10612
rect 12292 10556 13020 10612
rect 13076 10556 13086 10612
rect 14018 10556 14028 10612
rect 14084 10556 14812 10612
rect 14868 10556 19852 10612
rect 19908 10556 22988 10612
rect 23044 10556 23054 10612
rect 27570 10556 27580 10612
rect 27636 10556 28560 10612
rect 28448 10528 28560 10556
rect 11974 10444 12012 10500
rect 12068 10444 12078 10500
rect 0 10332 5180 10388
rect 5236 10332 5246 10388
rect 8082 10332 8092 10388
rect 8148 10332 9548 10388
rect 9604 10332 9614 10388
rect 10882 10332 10892 10388
rect 10948 10332 10958 10388
rect 11218 10332 11228 10388
rect 11284 10332 13692 10388
rect 13748 10332 13758 10388
rect 0 10304 112 10332
rect 6178 10220 6188 10276
rect 6244 10220 8204 10276
rect 8260 10220 8270 10276
rect 11442 10220 11452 10276
rect 11508 10220 12348 10276
rect 12404 10220 12414 10276
rect 16818 10220 16828 10276
rect 16884 10220 17724 10276
rect 17780 10220 20860 10276
rect 20916 10220 20926 10276
rect 4454 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4738 10220
rect 24454 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24738 10220
rect 28448 10164 28560 10192
rect 7074 10108 7084 10164
rect 7140 10108 7644 10164
rect 7700 10108 7710 10164
rect 8306 10108 8316 10164
rect 8372 10108 10108 10164
rect 10164 10108 10174 10164
rect 11666 10108 11676 10164
rect 11732 10108 15148 10164
rect 15204 10108 16044 10164
rect 16100 10108 16110 10164
rect 16258 10108 16268 10164
rect 16324 10108 18060 10164
rect 18116 10108 19404 10164
rect 19460 10108 19470 10164
rect 26562 10108 26572 10164
rect 26628 10108 28560 10164
rect 28448 10080 28560 10108
rect 2482 9996 2492 10052
rect 2548 9996 2716 10052
rect 2772 9996 2940 10052
rect 2996 9996 3006 10052
rect 6514 9996 6524 10052
rect 6580 9996 6972 10052
rect 7028 9996 7532 10052
rect 7588 9996 8988 10052
rect 9044 9996 9054 10052
rect 14578 9996 14588 10052
rect 14644 9996 15036 10052
rect 15092 9996 15102 10052
rect 16482 9996 16492 10052
rect 16548 9996 17276 10052
rect 17332 9996 17342 10052
rect 17826 9996 17836 10052
rect 17892 9996 18956 10052
rect 19012 9996 19022 10052
rect 21858 9996 21868 10052
rect 21924 9996 25676 10052
rect 25732 9996 25742 10052
rect 2940 9940 2996 9996
rect 2940 9884 5292 9940
rect 5348 9884 5358 9940
rect 7858 9884 7868 9940
rect 7924 9884 8876 9940
rect 8932 9884 8942 9940
rect 11890 9884 11900 9940
rect 11956 9884 12124 9940
rect 12180 9884 13132 9940
rect 13188 9884 13804 9940
rect 13860 9884 13870 9940
rect 15092 9884 16940 9940
rect 16996 9884 17006 9940
rect 17602 9884 17612 9940
rect 17668 9884 19292 9940
rect 19348 9884 26348 9940
rect 26404 9884 26414 9940
rect 15092 9828 15148 9884
rect 3826 9772 3836 9828
rect 3892 9772 15148 9828
rect 15372 9772 17052 9828
rect 17108 9772 17118 9828
rect 17266 9772 17276 9828
rect 17332 9772 17724 9828
rect 17780 9772 17790 9828
rect 21074 9772 21084 9828
rect 21140 9772 22876 9828
rect 22932 9772 22942 9828
rect 15372 9716 15428 9772
rect 28448 9716 28560 9744
rect 15138 9660 15148 9716
rect 15204 9660 15372 9716
rect 15428 9660 15438 9716
rect 15586 9660 15596 9716
rect 15652 9660 16044 9716
rect 16100 9660 25116 9716
rect 25172 9660 25182 9716
rect 26562 9660 26572 9716
rect 26628 9660 28560 9716
rect 28448 9632 28560 9660
rect 9986 9548 9996 9604
rect 10052 9548 10332 9604
rect 10388 9548 10398 9604
rect 12338 9548 12348 9604
rect 12404 9548 14028 9604
rect 14084 9548 14094 9604
rect 15474 9548 15484 9604
rect 15540 9548 15708 9604
rect 15764 9548 16604 9604
rect 16660 9548 16670 9604
rect 27458 9548 27468 9604
rect 27524 9548 28140 9604
rect 28196 9548 28206 9604
rect 0 9492 112 9520
rect 0 9436 2940 9492
rect 2996 9436 3006 9492
rect 12226 9436 12236 9492
rect 12292 9436 16156 9492
rect 16212 9436 17836 9492
rect 17892 9436 17902 9492
rect 0 9408 112 9436
rect 3794 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4078 9436
rect 23794 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24078 9436
rect 6850 9324 6860 9380
rect 6916 9324 7308 9380
rect 7364 9324 17612 9380
rect 17668 9324 17678 9380
rect 27234 9324 27244 9380
rect 27300 9324 27692 9380
rect 27748 9324 27758 9380
rect 28448 9268 28560 9296
rect 802 9212 812 9268
rect 868 9212 1260 9268
rect 1316 9212 1326 9268
rect 12450 9212 12460 9268
rect 12516 9212 13244 9268
rect 13300 9212 13310 9268
rect 25666 9212 25676 9268
rect 25732 9212 28560 9268
rect 28448 9184 28560 9212
rect 5478 9100 5516 9156
rect 5572 9100 5582 9156
rect 6374 9100 6412 9156
rect 6468 9100 6478 9156
rect 7410 9100 7420 9156
rect 7476 9100 9884 9156
rect 9940 9100 9950 9156
rect 11330 9100 11340 9156
rect 11396 9100 26012 9156
rect 26068 9100 26078 9156
rect 9314 8988 9324 9044
rect 9380 8988 10444 9044
rect 10500 8988 12796 9044
rect 12852 8988 12862 9044
rect 13020 8988 18172 9044
rect 18228 8988 18238 9044
rect 20850 8988 20860 9044
rect 20916 8988 26460 9044
rect 26516 8988 26526 9044
rect 12114 8876 12124 8932
rect 12180 8876 12348 8932
rect 12404 8876 12414 8932
rect 13020 8820 13076 8988
rect 28448 8820 28560 8848
rect 10882 8764 10892 8820
rect 10948 8764 13076 8820
rect 15092 8764 15372 8820
rect 15428 8764 15438 8820
rect 25890 8764 25900 8820
rect 25956 8764 28560 8820
rect 15092 8708 15148 8764
rect 28448 8736 28560 8764
rect 2146 8652 2156 8708
rect 2212 8652 3164 8708
rect 3220 8652 3230 8708
rect 7186 8652 7196 8708
rect 7252 8652 8540 8708
rect 8596 8652 11564 8708
rect 11620 8652 15148 8708
rect 0 8596 112 8624
rect 4454 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4738 8652
rect 24454 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24738 8652
rect 0 8540 1428 8596
rect 8082 8540 8092 8596
rect 8148 8540 9380 8596
rect 9650 8540 9660 8596
rect 9716 8540 13356 8596
rect 13412 8540 13422 8596
rect 0 8512 112 8540
rect 1372 8260 1428 8540
rect 9324 8484 9380 8540
rect 5506 8428 5516 8484
rect 5572 8428 8428 8484
rect 8484 8428 8494 8484
rect 9314 8428 9324 8484
rect 9380 8428 9996 8484
rect 10052 8428 12964 8484
rect 13906 8428 13916 8484
rect 13972 8428 14924 8484
rect 14980 8428 14990 8484
rect 17826 8428 17836 8484
rect 17892 8428 19516 8484
rect 19572 8428 26012 8484
rect 26068 8428 26078 8484
rect 12908 8372 12964 8428
rect 28448 8372 28560 8400
rect 6178 8316 6188 8372
rect 6244 8316 6860 8372
rect 6916 8316 9772 8372
rect 9828 8316 9838 8372
rect 10210 8316 10220 8372
rect 10276 8316 11116 8372
rect 11172 8316 11182 8372
rect 12898 8316 12908 8372
rect 12964 8316 12974 8372
rect 13458 8316 13468 8372
rect 13524 8316 15596 8372
rect 15652 8316 18844 8372
rect 18900 8316 20300 8372
rect 20356 8316 20366 8372
rect 27234 8316 27244 8372
rect 27300 8316 28560 8372
rect 28448 8288 28560 8316
rect 1372 8204 1596 8260
rect 1652 8204 1662 8260
rect 7074 8204 7084 8260
rect 7140 8204 14252 8260
rect 14308 8204 14812 8260
rect 14868 8204 14878 8260
rect 15250 8204 15260 8260
rect 15316 8204 16940 8260
rect 16996 8204 17006 8260
rect 20066 8204 20076 8260
rect 20132 8204 21308 8260
rect 21364 8204 21644 8260
rect 21700 8204 21710 8260
rect 22530 8204 22540 8260
rect 22596 8204 22876 8260
rect 22932 8204 22942 8260
rect 27570 8204 27580 8260
rect 27636 8204 27646 8260
rect 27580 8148 27636 8204
rect 7746 8092 7756 8148
rect 7812 8092 21868 8148
rect 21924 8092 21934 8148
rect 27234 8092 27244 8148
rect 27300 8092 27636 8148
rect 2258 7980 2268 8036
rect 2324 7980 5068 8036
rect 5124 7980 5134 8036
rect 15026 7980 15036 8036
rect 15092 7980 15372 8036
rect 15428 7980 15438 8036
rect 16146 7980 16156 8036
rect 16212 7980 16716 8036
rect 16772 7980 16782 8036
rect 19058 7980 19068 8036
rect 19124 7980 26124 8036
rect 26180 7980 26190 8036
rect 28448 7924 28560 7952
rect 14802 7868 14812 7924
rect 14868 7868 16660 7924
rect 27458 7868 27468 7924
rect 27524 7868 28560 7924
rect 3794 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4078 7868
rect 16604 7812 16660 7868
rect 23794 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24078 7868
rect 28448 7840 28560 7868
rect 16594 7756 16604 7812
rect 16660 7756 17052 7812
rect 17108 7756 17118 7812
rect 0 7700 112 7728
rect 0 7644 1316 7700
rect 2370 7644 2380 7700
rect 2436 7644 3388 7700
rect 7270 7644 7308 7700
rect 7364 7644 7374 7700
rect 16706 7644 16716 7700
rect 16772 7644 17388 7700
rect 17444 7644 17454 7700
rect 20290 7644 20300 7700
rect 20356 7644 26908 7700
rect 26964 7644 26974 7700
rect 0 7616 112 7644
rect 1260 7588 1316 7644
rect 3332 7588 3388 7644
rect 1260 7532 2492 7588
rect 2548 7532 2558 7588
rect 3332 7532 22652 7588
rect 22708 7532 22718 7588
rect 27010 7532 27020 7588
rect 27076 7532 28140 7588
rect 28196 7532 28206 7588
rect 28448 7476 28560 7504
rect 3826 7420 3836 7476
rect 3892 7420 13580 7476
rect 13636 7420 13646 7476
rect 14578 7420 14588 7476
rect 14644 7420 15484 7476
rect 15540 7420 16156 7476
rect 16212 7420 16222 7476
rect 16930 7420 16940 7476
rect 16996 7420 17388 7476
rect 17444 7420 22540 7476
rect 22596 7420 25340 7476
rect 25396 7420 25406 7476
rect 26114 7420 26124 7476
rect 26180 7420 26684 7476
rect 26740 7420 26750 7476
rect 27346 7420 27356 7476
rect 27412 7420 28560 7476
rect 28448 7392 28560 7420
rect 9762 7308 9772 7364
rect 9828 7308 10668 7364
rect 10724 7308 11004 7364
rect 11060 7308 11070 7364
rect 14914 7308 14924 7364
rect 14980 7308 15596 7364
rect 15652 7308 16380 7364
rect 16436 7308 16446 7364
rect 27430 7308 27468 7364
rect 27524 7308 27534 7364
rect 11218 7196 11228 7252
rect 11284 7196 15708 7252
rect 15764 7196 20076 7252
rect 20132 7196 20142 7252
rect 13234 7084 13244 7140
rect 13300 7084 14812 7140
rect 14868 7084 14878 7140
rect 4454 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4738 7084
rect 24454 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24738 7084
rect 28448 7028 28560 7056
rect 13010 6972 13020 7028
rect 13076 6972 13356 7028
rect 13412 6972 13422 7028
rect 27458 6972 27468 7028
rect 27524 6972 28560 7028
rect 28448 6944 28560 6972
rect 0 6804 112 6832
rect 0 6748 1484 6804
rect 1540 6748 1550 6804
rect 10994 6748 11004 6804
rect 11060 6748 12684 6804
rect 12740 6748 12750 6804
rect 21634 6748 21644 6804
rect 21700 6748 26012 6804
rect 26068 6748 26078 6804
rect 0 6720 112 6748
rect 11554 6636 11564 6692
rect 11620 6636 19292 6692
rect 19348 6636 19358 6692
rect 21298 6636 21308 6692
rect 21364 6636 23324 6692
rect 23380 6636 23390 6692
rect 28448 6580 28560 6608
rect 3826 6524 3836 6580
rect 3892 6524 16492 6580
rect 16548 6524 16558 6580
rect 18498 6524 18508 6580
rect 18564 6524 22428 6580
rect 22484 6524 22494 6580
rect 26562 6524 26572 6580
rect 26628 6524 28560 6580
rect 28448 6496 28560 6524
rect 3490 6412 3500 6468
rect 3556 6412 22764 6468
rect 22820 6412 22830 6468
rect 3794 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4078 6300
rect 23794 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24078 6300
rect 28448 6132 28560 6160
rect 6066 6076 6076 6132
rect 6132 6076 7756 6132
rect 7812 6076 7822 6132
rect 26674 6076 26684 6132
rect 26740 6076 28560 6132
rect 28448 6048 28560 6076
rect 0 5908 112 5936
rect 0 5852 2828 5908
rect 2884 5852 2894 5908
rect 12226 5852 12236 5908
rect 12292 5852 24892 5908
rect 24948 5852 24958 5908
rect 0 5824 112 5852
rect 3154 5740 3164 5796
rect 3220 5740 25564 5796
rect 25620 5740 25630 5796
rect 28448 5684 28560 5712
rect 14802 5628 14812 5684
rect 14868 5628 15372 5684
rect 15428 5628 15438 5684
rect 25890 5628 25900 5684
rect 25956 5628 28560 5684
rect 28448 5600 28560 5628
rect 690 5516 700 5572
rect 756 5516 1596 5572
rect 1652 5516 1662 5572
rect 4454 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4738 5516
rect 24454 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24738 5516
rect 8306 5404 8316 5460
rect 8372 5404 19068 5460
rect 19124 5404 19134 5460
rect 7746 5292 7756 5348
rect 7812 5292 8876 5348
rect 8932 5292 11116 5348
rect 11172 5292 11182 5348
rect 11554 5292 11564 5348
rect 11620 5292 13804 5348
rect 13860 5292 14476 5348
rect 14532 5292 14542 5348
rect 15922 5292 15932 5348
rect 15988 5292 27692 5348
rect 27748 5292 27758 5348
rect 28448 5236 28560 5264
rect 17938 5180 17948 5236
rect 18004 5180 26684 5236
rect 26740 5180 26750 5236
rect 27346 5180 27356 5236
rect 27412 5180 28560 5236
rect 28448 5152 28560 5180
rect 4050 5068 4060 5124
rect 4116 5068 6636 5124
rect 6692 5068 6702 5124
rect 8754 5068 8764 5124
rect 8820 5068 15708 5124
rect 15764 5068 15774 5124
rect 0 5012 112 5040
rect 0 4956 1036 5012
rect 1092 4956 1102 5012
rect 6514 4956 6524 5012
rect 6580 4956 7980 5012
rect 8036 4956 8046 5012
rect 0 4928 112 4956
rect 15474 4844 15484 4900
rect 15540 4844 27804 4900
rect 27860 4844 27870 4900
rect 28448 4788 28560 4816
rect 27458 4732 27468 4788
rect 27524 4732 28560 4788
rect 3794 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4078 4732
rect 23794 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24078 4732
rect 28448 4704 28560 4732
rect 11554 4508 11564 4564
rect 11620 4508 28252 4564
rect 28308 4508 28318 4564
rect 6626 4396 6636 4452
rect 6692 4396 27692 4452
rect 27748 4396 27758 4452
rect 28448 4340 28560 4368
rect 2034 4284 2044 4340
rect 2100 4284 27244 4340
rect 27300 4284 27310 4340
rect 27458 4284 27468 4340
rect 27524 4284 28560 4340
rect 28448 4256 28560 4284
rect 2258 4172 2268 4228
rect 2324 4172 17500 4228
rect 17556 4172 17566 4228
rect 18834 4172 18844 4228
rect 18900 4172 26908 4228
rect 26964 4172 26974 4228
rect 0 4116 112 4144
rect 0 4060 1484 4116
rect 1540 4060 1550 4116
rect 0 4032 112 4060
rect 4454 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4738 3948
rect 24454 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24738 3948
rect 28448 3892 28560 3920
rect 27458 3836 27468 3892
rect 27524 3836 28560 3892
rect 28448 3808 28560 3836
rect 26898 3612 26908 3668
rect 26964 3612 27580 3668
rect 27636 3612 27646 3668
rect 2258 3500 2268 3556
rect 2324 3500 21980 3556
rect 22036 3500 22046 3556
rect 28448 3444 28560 3472
rect 27458 3388 27468 3444
rect 27524 3388 28560 3444
rect 28448 3360 28560 3388
rect 0 3220 112 3248
rect 0 3164 1260 3220
rect 1316 3164 1326 3220
rect 0 3136 112 3164
rect 3794 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4078 3164
rect 23794 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24078 3164
rect 28448 2996 28560 3024
rect 26562 2940 26572 2996
rect 26628 2940 28560 2996
rect 28448 2912 28560 2940
rect 354 2828 364 2884
rect 420 2828 1484 2884
rect 1540 2828 1550 2884
rect 18050 2716 18060 2772
rect 18116 2716 25564 2772
rect 25620 2716 25630 2772
rect 28448 2548 28560 2576
rect 26562 2492 26572 2548
rect 26628 2492 28560 2548
rect 28448 2464 28560 2492
rect 0 2324 112 2352
rect 4454 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4738 2380
rect 24454 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24738 2380
rect 0 2268 1036 2324
rect 1092 2268 1102 2324
rect 0 2240 112 2268
rect 23314 2156 23324 2212
rect 23380 2156 27468 2212
rect 27524 2156 27534 2212
rect 28448 2100 28560 2128
rect 13234 2044 13244 2100
rect 13300 2044 18508 2100
rect 18564 2044 18574 2100
rect 25778 2044 25788 2100
rect 25844 2044 28560 2100
rect 28448 2016 28560 2044
rect 13794 1932 13804 1988
rect 13860 1932 22204 1988
rect 22260 1932 22270 1988
rect 21634 1820 21644 1876
rect 21700 1820 25228 1876
rect 25284 1820 25294 1876
rect 28448 1652 28560 1680
rect 914 1596 924 1652
rect 980 1596 3388 1652
rect 3444 1596 3454 1652
rect 16706 1596 16716 1652
rect 16772 1596 16828 1652
rect 16884 1596 16894 1652
rect 20822 1596 20860 1652
rect 20916 1596 20926 1652
rect 27122 1596 27132 1652
rect 27188 1596 28560 1652
rect 3794 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4078 1596
rect 23794 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24078 1596
rect 28448 1568 28560 1596
rect 22418 1372 22428 1428
rect 22484 1372 26572 1428
rect 26628 1372 26638 1428
rect 12786 1260 12796 1316
rect 12852 1260 16044 1316
rect 16100 1260 16110 1316
rect 18162 1260 18172 1316
rect 18228 1260 26012 1316
rect 26068 1260 26078 1316
rect 28448 1204 28560 1232
rect 25554 1148 25564 1204
rect 25620 1148 28560 1204
rect 28448 1120 28560 1148
rect 23538 1036 23548 1092
rect 23604 1036 27020 1092
rect 27076 1036 27086 1092
rect 10098 924 10108 980
rect 10164 924 11900 980
rect 11956 924 11966 980
rect 14130 924 14140 980
rect 14196 924 21420 980
rect 21476 924 21486 980
rect 4454 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4738 812
rect 24454 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24738 812
rect 28448 756 28560 784
rect 25330 700 25340 756
rect 25396 700 28560 756
rect 28448 672 28560 700
rect 690 588 700 644
rect 756 588 10892 644
rect 10948 588 10958 644
rect 12002 588 12012 644
rect 12068 588 26236 644
rect 26292 588 26302 644
rect 4722 364 4732 420
rect 4788 364 8428 420
rect 8484 364 8494 420
rect 18386 364 18396 420
rect 18452 364 24892 420
rect 24948 364 24958 420
rect 28448 308 28560 336
rect 26338 252 26348 308
rect 26404 252 28560 308
rect 28448 224 28560 252
rect 19506 140 19516 196
rect 19572 140 26908 196
rect 26964 140 26974 196
<< via3 >>
rect 3804 56420 3860 56476
rect 3908 56420 3964 56476
rect 4012 56420 4068 56476
rect 23804 56420 23860 56476
rect 23908 56420 23964 56476
rect 24012 56420 24068 56476
rect 3052 55916 3108 55972
rect 21308 55916 21364 55972
rect 4464 55636 4520 55692
rect 4568 55636 4624 55692
rect 4672 55636 4728 55692
rect 24464 55636 24520 55692
rect 24568 55636 24624 55692
rect 24672 55636 24728 55692
rect 22428 55244 22484 55300
rect 26124 55244 26180 55300
rect 3804 54852 3860 54908
rect 3908 54852 3964 54908
rect 4012 54852 4068 54908
rect 23804 54852 23860 54908
rect 23908 54852 23964 54908
rect 24012 54852 24068 54908
rect 21756 54460 21812 54516
rect 4464 54068 4520 54124
rect 4568 54068 4624 54124
rect 4672 54068 4728 54124
rect 24464 54068 24520 54124
rect 24568 54068 24624 54124
rect 24672 54068 24728 54124
rect 12572 53900 12628 53956
rect 3804 53284 3860 53340
rect 3908 53284 3964 53340
rect 4012 53284 4068 53340
rect 23804 53284 23860 53340
rect 23908 53284 23964 53340
rect 24012 53284 24068 53340
rect 4464 52500 4520 52556
rect 4568 52500 4624 52556
rect 4672 52500 4728 52556
rect 24464 52500 24520 52556
rect 24568 52500 24624 52556
rect 24672 52500 24728 52556
rect 20860 52108 20916 52164
rect 22764 52108 22820 52164
rect 3804 51716 3860 51772
rect 3908 51716 3964 51772
rect 4012 51716 4068 51772
rect 23804 51716 23860 51772
rect 23908 51716 23964 51772
rect 24012 51716 24068 51772
rect 14140 51100 14196 51156
rect 4464 50932 4520 50988
rect 4568 50932 4624 50988
rect 4672 50932 4728 50988
rect 24464 50932 24520 50988
rect 24568 50932 24624 50988
rect 24672 50932 24728 50988
rect 27020 50764 27076 50820
rect 10780 50652 10836 50708
rect 18396 50540 18452 50596
rect 3804 50148 3860 50204
rect 3908 50148 3964 50204
rect 4012 50148 4068 50204
rect 23804 50148 23860 50204
rect 23908 50148 23964 50204
rect 24012 50148 24068 50204
rect 9212 49644 9268 49700
rect 4464 49364 4520 49420
rect 4568 49364 4624 49420
rect 4672 49364 4728 49420
rect 24464 49364 24520 49420
rect 24568 49364 24624 49420
rect 24672 49364 24728 49420
rect 16268 49196 16324 49252
rect 6300 48972 6356 49028
rect 14812 48860 14868 48916
rect 3804 48580 3860 48636
rect 3908 48580 3964 48636
rect 4012 48580 4068 48636
rect 23804 48580 23860 48636
rect 23908 48580 23964 48636
rect 24012 48580 24068 48636
rect 16716 48076 16772 48132
rect 4464 47796 4520 47852
rect 4568 47796 4624 47852
rect 4672 47796 4728 47852
rect 24464 47796 24520 47852
rect 24568 47796 24624 47852
rect 24672 47796 24728 47852
rect 19292 47404 19348 47460
rect 3804 47012 3860 47068
rect 3908 47012 3964 47068
rect 4012 47012 4068 47068
rect 23804 47012 23860 47068
rect 23908 47012 23964 47068
rect 24012 47012 24068 47068
rect 1484 46284 1540 46340
rect 4464 46228 4520 46284
rect 4568 46228 4624 46284
rect 4672 46228 4728 46284
rect 24464 46228 24520 46284
rect 24568 46228 24624 46284
rect 24672 46228 24728 46284
rect 3804 45444 3860 45500
rect 3908 45444 3964 45500
rect 4012 45444 4068 45500
rect 23804 45444 23860 45500
rect 23908 45444 23964 45500
rect 24012 45444 24068 45500
rect 4464 44660 4520 44716
rect 4568 44660 4624 44716
rect 4672 44660 4728 44716
rect 24464 44660 24520 44716
rect 24568 44660 24624 44716
rect 24672 44660 24728 44716
rect 1596 44380 1652 44436
rect 3804 43876 3860 43932
rect 3908 43876 3964 43932
rect 4012 43876 4068 43932
rect 23804 43876 23860 43932
rect 23908 43876 23964 43932
rect 24012 43876 24068 43932
rect 1708 43708 1764 43764
rect 4464 43092 4520 43148
rect 4568 43092 4624 43148
rect 4672 43092 4728 43148
rect 24464 43092 24520 43148
rect 24568 43092 24624 43148
rect 24672 43092 24728 43148
rect 3804 42308 3860 42364
rect 3908 42308 3964 42364
rect 4012 42308 4068 42364
rect 23804 42308 23860 42364
rect 23908 42308 23964 42364
rect 24012 42308 24068 42364
rect 11228 41804 11284 41860
rect 1708 41580 1764 41636
rect 4464 41524 4520 41580
rect 4568 41524 4624 41580
rect 4672 41524 4728 41580
rect 24464 41524 24520 41580
rect 24568 41524 24624 41580
rect 24672 41524 24728 41580
rect 5516 41468 5572 41524
rect 1596 41244 1652 41300
rect 3804 40740 3860 40796
rect 3908 40740 3964 40796
rect 4012 40740 4068 40796
rect 23804 40740 23860 40796
rect 23908 40740 23964 40796
rect 24012 40740 24068 40796
rect 4464 39956 4520 40012
rect 4568 39956 4624 40012
rect 4672 39956 4728 40012
rect 24464 39956 24520 40012
rect 24568 39956 24624 40012
rect 24672 39956 24728 40012
rect 7308 39788 7364 39844
rect 26908 39676 26964 39732
rect 8428 39564 8484 39620
rect 3804 39172 3860 39228
rect 3908 39172 3964 39228
rect 4012 39172 4068 39228
rect 23804 39172 23860 39228
rect 23908 39172 23964 39228
rect 24012 39172 24068 39228
rect 4464 38388 4520 38444
rect 4568 38388 4624 38444
rect 4672 38388 4728 38444
rect 24464 38388 24520 38444
rect 24568 38388 24624 38444
rect 24672 38388 24728 38444
rect 3804 37604 3860 37660
rect 3908 37604 3964 37660
rect 4012 37604 4068 37660
rect 23804 37604 23860 37660
rect 23908 37604 23964 37660
rect 24012 37604 24068 37660
rect 1484 36876 1540 36932
rect 4464 36820 4520 36876
rect 4568 36820 4624 36876
rect 4672 36820 4728 36876
rect 24464 36820 24520 36876
rect 24568 36820 24624 36876
rect 24672 36820 24728 36876
rect 3804 36036 3860 36092
rect 3908 36036 3964 36092
rect 4012 36036 4068 36092
rect 23804 36036 23860 36092
rect 23908 36036 23964 36092
rect 24012 36036 24068 36092
rect 1260 35644 1316 35700
rect 1596 35644 1652 35700
rect 9884 35308 9940 35364
rect 4464 35252 4520 35308
rect 4568 35252 4624 35308
rect 4672 35252 4728 35308
rect 24464 35252 24520 35308
rect 24568 35252 24624 35308
rect 24672 35252 24728 35308
rect 2940 35196 2996 35252
rect 10444 35196 10500 35252
rect 1372 35084 1428 35140
rect 10892 34860 10948 34916
rect 3804 34468 3860 34524
rect 3908 34468 3964 34524
rect 4012 34468 4068 34524
rect 23804 34468 23860 34524
rect 23908 34468 23964 34524
rect 24012 34468 24068 34524
rect 1596 34412 1652 34468
rect 8876 34412 8932 34468
rect 14028 34412 14084 34468
rect 1372 34076 1428 34132
rect 9660 33964 9716 34020
rect 4464 33684 4520 33740
rect 4568 33684 4624 33740
rect 4672 33684 4728 33740
rect 24464 33684 24520 33740
rect 24568 33684 24624 33740
rect 24672 33684 24728 33740
rect 3052 33628 3108 33684
rect 4284 33404 4340 33460
rect 6748 33404 6804 33460
rect 11676 32956 11732 33012
rect 3804 32900 3860 32956
rect 3908 32900 3964 32956
rect 4012 32900 4068 32956
rect 23804 32900 23860 32956
rect 23908 32900 23964 32956
rect 24012 32900 24068 32956
rect 10220 32844 10276 32900
rect 4956 32732 5012 32788
rect 13244 32508 13300 32564
rect 1260 32396 1316 32452
rect 4284 32396 4340 32452
rect 4464 32116 4520 32172
rect 4568 32116 4624 32172
rect 4672 32116 4728 32172
rect 24464 32116 24520 32172
rect 24568 32116 24624 32172
rect 24672 32116 24728 32172
rect 13468 32060 13524 32116
rect 9660 31836 9716 31892
rect 13132 31836 13188 31892
rect 1260 31724 1316 31780
rect 7420 31612 7476 31668
rect 10668 31612 10724 31668
rect 26348 31388 26404 31444
rect 3804 31332 3860 31388
rect 3908 31332 3964 31388
rect 4012 31332 4068 31388
rect 23804 31332 23860 31388
rect 23908 31332 23964 31388
rect 24012 31332 24068 31388
rect 13244 31276 13300 31332
rect 13692 30716 13748 30772
rect 4464 30548 4520 30604
rect 4568 30548 4624 30604
rect 4672 30548 4728 30604
rect 24464 30548 24520 30604
rect 24568 30548 24624 30604
rect 24672 30548 24728 30604
rect 11004 30380 11060 30436
rect 23548 30044 23604 30100
rect 2940 29820 2996 29876
rect 3804 29764 3860 29820
rect 3908 29764 3964 29820
rect 4012 29764 4068 29820
rect 23804 29764 23860 29820
rect 23908 29764 23964 29820
rect 24012 29764 24068 29820
rect 4956 29372 5012 29428
rect 11004 29372 11060 29428
rect 7420 29260 7476 29316
rect 8764 29260 8820 29316
rect 26348 29260 26404 29316
rect 11004 29148 11060 29204
rect 4464 28980 4520 29036
rect 4568 28980 4624 29036
rect 4672 28980 4728 29036
rect 24464 28980 24520 29036
rect 24568 28980 24624 29036
rect 24672 28980 24728 29036
rect 2380 28700 2436 28756
rect 8876 28700 8932 28756
rect 11676 28476 11732 28532
rect 16044 28364 16100 28420
rect 7980 28252 8036 28308
rect 3804 28196 3860 28252
rect 3908 28196 3964 28252
rect 4012 28196 4068 28252
rect 23804 28196 23860 28252
rect 23908 28196 23964 28252
rect 24012 28196 24068 28252
rect 10668 28028 10724 28084
rect 26236 27692 26292 27748
rect 4464 27412 4520 27468
rect 4568 27412 4624 27468
rect 4672 27412 4728 27468
rect 24464 27412 24520 27468
rect 24568 27412 24624 27468
rect 24672 27412 24728 27468
rect 10108 27244 10164 27300
rect 11228 27244 11284 27300
rect 13468 27132 13524 27188
rect 1260 27020 1316 27076
rect 5292 27020 5348 27076
rect 5404 26908 5460 26964
rect 7980 26908 8036 26964
rect 15932 26796 15988 26852
rect 13132 26684 13188 26740
rect 14028 26684 14084 26740
rect 3804 26628 3860 26684
rect 3908 26628 3964 26684
rect 4012 26628 4068 26684
rect 23804 26628 23860 26684
rect 23908 26628 23964 26684
rect 24012 26628 24068 26684
rect 6188 26348 6244 26404
rect 6188 26124 6244 26180
rect 25228 26124 25284 26180
rect 6748 26012 6804 26068
rect 10108 26012 10164 26068
rect 15932 25900 15988 25956
rect 4464 25844 4520 25900
rect 4568 25844 4624 25900
rect 4672 25844 4728 25900
rect 24464 25844 24520 25900
rect 24568 25844 24624 25900
rect 24672 25844 24728 25900
rect 10220 25452 10276 25508
rect 3804 25060 3860 25116
rect 3908 25060 3964 25116
rect 4012 25060 4068 25116
rect 23804 25060 23860 25116
rect 23908 25060 23964 25116
rect 24012 25060 24068 25116
rect 5404 25004 5460 25060
rect 9660 25004 9716 25060
rect 13692 24892 13748 24948
rect 26236 24780 26292 24836
rect 2380 24556 2436 24612
rect 7980 24444 8036 24500
rect 4464 24276 4520 24332
rect 4568 24276 4624 24332
rect 4672 24276 4728 24332
rect 24464 24276 24520 24332
rect 24568 24276 24624 24332
rect 24672 24276 24728 24332
rect 10220 23996 10276 24052
rect 20636 23884 20692 23940
rect 11004 23772 11060 23828
rect 4172 23660 4228 23716
rect 5292 23548 5348 23604
rect 16268 23548 16324 23604
rect 3804 23492 3860 23548
rect 3908 23492 3964 23548
rect 4012 23492 4068 23548
rect 23804 23492 23860 23548
rect 23908 23492 23964 23548
rect 24012 23492 24068 23548
rect 20076 23100 20132 23156
rect 14140 22988 14196 23044
rect 18620 22988 18676 23044
rect 20636 22876 20692 22932
rect 4464 22708 4520 22764
rect 4568 22708 4624 22764
rect 4672 22708 4728 22764
rect 24464 22708 24520 22764
rect 24568 22708 24624 22764
rect 24672 22708 24728 22764
rect 19516 22092 19572 22148
rect 19964 22092 20020 22148
rect 3804 21924 3860 21980
rect 3908 21924 3964 21980
rect 4012 21924 4068 21980
rect 12012 21868 12068 21924
rect 23804 21924 23860 21980
rect 23908 21924 23964 21980
rect 24012 21924 24068 21980
rect 2380 21532 2436 21588
rect 23548 21532 23604 21588
rect 27132 21420 27188 21476
rect 9996 21196 10052 21252
rect 4464 21140 4520 21196
rect 4568 21140 4624 21196
rect 4672 21140 4728 21196
rect 24464 21140 24520 21196
rect 24568 21140 24624 21196
rect 24672 21140 24728 21196
rect 8540 21084 8596 21140
rect 19964 21084 20020 21140
rect 25900 20748 25956 20804
rect 25228 20636 25284 20692
rect 3804 20356 3860 20412
rect 3908 20356 3964 20412
rect 4012 20356 4068 20412
rect 23804 20356 23860 20412
rect 23908 20356 23964 20412
rect 24012 20356 24068 20412
rect 13468 20300 13524 20356
rect 13132 19964 13188 20020
rect 18732 19964 18788 20020
rect 20076 19964 20132 20020
rect 13356 19628 13412 19684
rect 4464 19572 4520 19628
rect 4568 19572 4624 19628
rect 4672 19572 4728 19628
rect 24464 19572 24520 19628
rect 24568 19572 24624 19628
rect 24672 19572 24728 19628
rect 9884 19292 9940 19348
rect 26908 19292 26964 19348
rect 12908 18956 12964 19012
rect 3804 18788 3860 18844
rect 3908 18788 3964 18844
rect 4012 18788 4068 18844
rect 23804 18788 23860 18844
rect 23908 18788 23964 18844
rect 24012 18788 24068 18844
rect 3612 18732 3668 18788
rect 13132 18732 13188 18788
rect 6300 18620 6356 18676
rect 18620 18508 18676 18564
rect 10220 18284 10276 18340
rect 12908 18284 12964 18340
rect 13356 18284 13412 18340
rect 18844 18172 18900 18228
rect 19068 18060 19124 18116
rect 4464 18004 4520 18060
rect 4568 18004 4624 18060
rect 4672 18004 4728 18060
rect 24464 18004 24520 18060
rect 24568 18004 24624 18060
rect 24672 18004 24728 18060
rect 19516 17612 19572 17668
rect 19404 17388 19460 17444
rect 14924 17276 14980 17332
rect 3804 17220 3860 17276
rect 3908 17220 3964 17276
rect 4012 17220 4068 17276
rect 23804 17220 23860 17276
rect 23908 17220 23964 17276
rect 24012 17220 24068 17276
rect 19628 17164 19684 17220
rect 26012 17052 26068 17108
rect 4172 16940 4228 16996
rect 14924 16940 14980 16996
rect 4284 16828 4340 16884
rect 9996 16828 10052 16884
rect 3612 16716 3668 16772
rect 13804 16716 13860 16772
rect 26908 16716 26964 16772
rect 4956 16492 5012 16548
rect 19068 16492 19124 16548
rect 4464 16436 4520 16492
rect 4568 16436 4624 16492
rect 4672 16436 4728 16492
rect 24464 16436 24520 16492
rect 24568 16436 24624 16492
rect 24672 16436 24728 16492
rect 18956 16380 19012 16436
rect 19404 16380 19460 16436
rect 19628 16380 19684 16436
rect 13804 16268 13860 16324
rect 10444 16156 10500 16212
rect 18732 16044 18788 16100
rect 18956 16044 19012 16100
rect 13468 15820 13524 15876
rect 19628 15820 19684 15876
rect 3804 15652 3860 15708
rect 3908 15652 3964 15708
rect 4012 15652 4068 15708
rect 23804 15652 23860 15708
rect 23908 15652 23964 15708
rect 24012 15652 24068 15708
rect 19628 15372 19684 15428
rect 19852 15372 19908 15428
rect 4464 14868 4520 14924
rect 4568 14868 4624 14924
rect 4672 14868 4728 14924
rect 24464 14868 24520 14924
rect 24568 14868 24624 14924
rect 24672 14868 24728 14924
rect 15372 14812 15428 14868
rect 19852 14812 19908 14868
rect 8540 14700 8596 14756
rect 19852 14588 19908 14644
rect 8316 14364 8372 14420
rect 9212 14140 9268 14196
rect 15372 14140 15428 14196
rect 15596 14140 15652 14196
rect 3804 14084 3860 14140
rect 3908 14084 3964 14140
rect 4012 14084 4068 14140
rect 23804 14084 23860 14140
rect 23908 14084 23964 14140
rect 24012 14084 24068 14140
rect 27132 13804 27188 13860
rect 21756 13580 21812 13636
rect 6412 13468 6468 13524
rect 8540 13468 8596 13524
rect 12572 13468 12628 13524
rect 12796 13468 12852 13524
rect 11676 13356 11732 13412
rect 13356 13356 13412 13412
rect 4464 13300 4520 13356
rect 4568 13300 4624 13356
rect 4672 13300 4728 13356
rect 24464 13300 24520 13356
rect 24568 13300 24624 13356
rect 24672 13300 24728 13356
rect 8316 13132 8372 13188
rect 9996 13020 10052 13076
rect 17836 13020 17892 13076
rect 19180 13020 19236 13076
rect 15596 12908 15652 12964
rect 18060 12796 18116 12852
rect 17164 12684 17220 12740
rect 17948 12684 18004 12740
rect 3804 12516 3860 12572
rect 3908 12516 3964 12572
rect 4012 12516 4068 12572
rect 23804 12516 23860 12572
rect 23908 12516 23964 12572
rect 24012 12516 24068 12572
rect 4956 12460 5012 12516
rect 12012 12460 12068 12516
rect 12796 12460 12852 12516
rect 17948 12348 18004 12404
rect 12460 12236 12516 12292
rect 9100 12124 9156 12180
rect 26012 12124 26068 12180
rect 12460 11900 12516 11956
rect 19516 11900 19572 11956
rect 25900 11900 25956 11956
rect 4464 11732 4520 11788
rect 4568 11732 4624 11788
rect 4672 11732 4728 11788
rect 17836 11788 17892 11844
rect 18060 11788 18116 11844
rect 19180 11788 19236 11844
rect 24464 11732 24520 11788
rect 24568 11732 24624 11788
rect 24672 11732 24728 11788
rect 26908 11452 26964 11508
rect 17164 11228 17220 11284
rect 10780 11116 10836 11172
rect 11676 11116 11732 11172
rect 9100 11004 9156 11060
rect 12012 11004 12068 11060
rect 17948 11004 18004 11060
rect 3804 10948 3860 11004
rect 3908 10948 3964 11004
rect 4012 10948 4068 11004
rect 23804 10948 23860 11004
rect 23908 10948 23964 11004
rect 24012 10948 24068 11004
rect 8764 10668 8820 10724
rect 12012 10444 12068 10500
rect 4464 10164 4520 10220
rect 4568 10164 4624 10220
rect 4672 10164 4728 10220
rect 24464 10164 24520 10220
rect 24568 10164 24624 10220
rect 24672 10164 24728 10220
rect 3804 9380 3860 9436
rect 3908 9380 3964 9436
rect 4012 9380 4068 9436
rect 23804 9380 23860 9436
rect 23908 9380 23964 9436
rect 24012 9380 24068 9436
rect 5516 9100 5572 9156
rect 6412 9100 6468 9156
rect 4464 8596 4520 8652
rect 4568 8596 4624 8652
rect 4672 8596 4728 8652
rect 24464 8596 24520 8652
rect 24568 8596 24624 8652
rect 24672 8596 24728 8652
rect 26124 7980 26180 8036
rect 27468 7868 27524 7924
rect 3804 7812 3860 7868
rect 3908 7812 3964 7868
rect 4012 7812 4068 7868
rect 23804 7812 23860 7868
rect 23908 7812 23964 7868
rect 24012 7812 24068 7868
rect 7308 7644 7364 7700
rect 27468 7308 27524 7364
rect 14812 7084 14868 7140
rect 4464 7028 4520 7084
rect 4568 7028 4624 7084
rect 4672 7028 4728 7084
rect 24464 7028 24520 7084
rect 24568 7028 24624 7084
rect 24672 7028 24728 7084
rect 19292 6636 19348 6692
rect 21308 6636 21364 6692
rect 22428 6524 22484 6580
rect 22764 6412 22820 6468
rect 3804 6244 3860 6300
rect 3908 6244 3964 6300
rect 4012 6244 4068 6300
rect 23804 6244 23860 6300
rect 23908 6244 23964 6300
rect 24012 6244 24068 6300
rect 4464 5460 4520 5516
rect 4568 5460 4624 5516
rect 4672 5460 4728 5516
rect 24464 5460 24520 5516
rect 24568 5460 24624 5516
rect 24672 5460 24728 5516
rect 3804 4676 3860 4732
rect 3908 4676 3964 4732
rect 4012 4676 4068 4732
rect 23804 4676 23860 4732
rect 23908 4676 23964 4732
rect 24012 4676 24068 4732
rect 18844 4172 18900 4228
rect 4464 3892 4520 3948
rect 4568 3892 4624 3948
rect 4672 3892 4728 3948
rect 24464 3892 24520 3948
rect 24568 3892 24624 3948
rect 24672 3892 24728 3948
rect 3804 3108 3860 3164
rect 3908 3108 3964 3164
rect 4012 3108 4068 3164
rect 23804 3108 23860 3164
rect 23908 3108 23964 3164
rect 24012 3108 24068 3164
rect 4464 2324 4520 2380
rect 4568 2324 4624 2380
rect 4672 2324 4728 2380
rect 24464 2324 24520 2380
rect 24568 2324 24624 2380
rect 24672 2324 24728 2380
rect 16716 1596 16772 1652
rect 20860 1596 20916 1652
rect 3804 1540 3860 1596
rect 3908 1540 3964 1596
rect 4012 1540 4068 1596
rect 23804 1540 23860 1596
rect 23908 1540 23964 1596
rect 24012 1540 24068 1596
rect 16044 1260 16100 1316
rect 27020 1036 27076 1092
rect 4464 756 4520 812
rect 4568 756 4624 812
rect 4672 756 4728 812
rect 24464 756 24520 812
rect 24568 756 24624 812
rect 24672 756 24728 812
rect 10892 588 10948 644
rect 8428 364 8484 420
rect 18396 364 18452 420
<< metal4 >>
rect 3776 56476 4096 57456
rect 3776 56420 3804 56476
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 4068 56420 4096 56476
rect 3052 55972 3108 55982
rect 1484 46340 1540 46350
rect 1484 36932 1540 46284
rect 1596 44436 1652 44446
rect 1596 41300 1652 44380
rect 1708 43764 1764 43774
rect 1708 41636 1764 43708
rect 1708 41570 1764 41580
rect 1596 41234 1652 41244
rect 1484 36866 1540 36876
rect 1260 35700 1316 35710
rect 1260 32452 1316 35644
rect 1596 35700 1652 35710
rect 1372 35140 1428 35150
rect 1372 34132 1428 35084
rect 1596 34468 1652 35644
rect 1596 34402 1652 34412
rect 2940 35252 2996 35262
rect 1372 34066 1428 34076
rect 1260 32386 1316 32396
rect 1260 31780 1316 31790
rect 1260 27076 1316 31724
rect 2940 29876 2996 35196
rect 3052 33684 3108 55916
rect 3052 33618 3108 33628
rect 3776 54908 4096 56420
rect 3776 54852 3804 54908
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 4068 54852 4096 54908
rect 3776 53340 4096 54852
rect 3776 53284 3804 53340
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 4068 53284 4096 53340
rect 3776 51772 4096 53284
rect 3776 51716 3804 51772
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 4068 51716 4096 51772
rect 3776 50204 4096 51716
rect 3776 50148 3804 50204
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 4068 50148 4096 50204
rect 3776 48636 4096 50148
rect 3776 48580 3804 48636
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 4068 48580 4096 48636
rect 3776 47068 4096 48580
rect 3776 47012 3804 47068
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 4068 47012 4096 47068
rect 3776 45500 4096 47012
rect 3776 45444 3804 45500
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 4068 45444 4096 45500
rect 3776 43932 4096 45444
rect 3776 43876 3804 43932
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 4068 43876 4096 43932
rect 3776 42364 4096 43876
rect 3776 42308 3804 42364
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 4068 42308 4096 42364
rect 3776 40796 4096 42308
rect 3776 40740 3804 40796
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 4068 40740 4096 40796
rect 3776 39228 4096 40740
rect 3776 39172 3804 39228
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 4068 39172 4096 39228
rect 3776 37660 4096 39172
rect 3776 37604 3804 37660
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 4068 37604 4096 37660
rect 3776 36092 4096 37604
rect 3776 36036 3804 36092
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 4068 36036 4096 36092
rect 3776 34524 4096 36036
rect 3776 34468 3804 34524
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 4068 34468 4096 34524
rect 2940 29810 2996 29820
rect 3776 32956 4096 34468
rect 4436 55692 4756 57456
rect 23776 56476 24096 57456
rect 23776 56420 23804 56476
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 24068 56420 24096 56476
rect 4436 55636 4464 55692
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4728 55636 4756 55692
rect 4436 54124 4756 55636
rect 4436 54068 4464 54124
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4728 54068 4756 54124
rect 4436 52556 4756 54068
rect 21308 55972 21364 55982
rect 4436 52500 4464 52556
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4728 52500 4756 52556
rect 4436 50988 4756 52500
rect 4436 50932 4464 50988
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4728 50932 4756 50988
rect 4436 49420 4756 50932
rect 12572 53956 12628 53966
rect 10780 50708 10836 50718
rect 4436 49364 4464 49420
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4728 49364 4756 49420
rect 4436 47852 4756 49364
rect 9212 49700 9268 49710
rect 4436 47796 4464 47852
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4728 47796 4756 47852
rect 4436 46284 4756 47796
rect 4436 46228 4464 46284
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4728 46228 4756 46284
rect 4436 44716 4756 46228
rect 4436 44660 4464 44716
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4728 44660 4756 44716
rect 4436 43148 4756 44660
rect 4436 43092 4464 43148
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4728 43092 4756 43148
rect 4436 41580 4756 43092
rect 4436 41524 4464 41580
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4728 41524 4756 41580
rect 6300 49028 6356 49038
rect 4436 40012 4756 41524
rect 4436 39956 4464 40012
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4728 39956 4756 40012
rect 4436 38444 4756 39956
rect 4436 38388 4464 38444
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4728 38388 4756 38444
rect 4436 36876 4756 38388
rect 4436 36820 4464 36876
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4728 36820 4756 36876
rect 4436 35308 4756 36820
rect 4436 35252 4464 35308
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4728 35252 4756 35308
rect 4436 33740 4756 35252
rect 4436 33684 4464 33740
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4728 33684 4756 33740
rect 3776 32900 3804 32956
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 4068 32900 4096 32956
rect 3776 31388 4096 32900
rect 3776 31332 3804 31388
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 4068 31332 4096 31388
rect 3776 29820 4096 31332
rect 3776 29764 3804 29820
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 4068 29764 4096 29820
rect 1260 27010 1316 27020
rect 2380 28756 2436 28766
rect 2380 24612 2436 28700
rect 2380 21588 2436 24556
rect 2380 21522 2436 21532
rect 3776 28252 4096 29764
rect 3776 28196 3804 28252
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 4068 28196 4096 28252
rect 3776 26684 4096 28196
rect 3776 26628 3804 26684
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 4068 26628 4096 26684
rect 3776 25116 4096 26628
rect 3776 25060 3804 25116
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 4068 25060 4096 25116
rect 3776 23548 4096 25060
rect 4284 33460 4340 33470
rect 4284 32452 4340 33404
rect 3776 23492 3804 23548
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 4068 23492 4096 23548
rect 3776 21980 4096 23492
rect 3776 21924 3804 21980
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 4068 21924 4096 21980
rect 3776 20412 4096 21924
rect 3776 20356 3804 20412
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 4068 20356 4096 20412
rect 3776 18844 4096 20356
rect 3612 18788 3668 18798
rect 3612 16772 3668 18732
rect 3612 16706 3668 16716
rect 3776 18788 3804 18844
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 4068 18788 4096 18844
rect 3776 17276 4096 18788
rect 3776 17220 3804 17276
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 4068 17220 4096 17276
rect 3776 15708 4096 17220
rect 4172 23716 4228 23726
rect 4172 16996 4228 23660
rect 4172 16930 4228 16940
rect 4284 16884 4340 32396
rect 4284 16818 4340 16828
rect 4436 32172 4756 33684
rect 5516 41524 5572 41534
rect 4436 32116 4464 32172
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4728 32116 4756 32172
rect 4436 30604 4756 32116
rect 4436 30548 4464 30604
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4728 30548 4756 30604
rect 4436 29036 4756 30548
rect 4956 32788 5012 32798
rect 4956 29428 5012 32732
rect 4956 29362 5012 29372
rect 4436 28980 4464 29036
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4728 28980 4756 29036
rect 4436 27468 4756 28980
rect 4436 27412 4464 27468
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4728 27412 4756 27468
rect 4436 25900 4756 27412
rect 4436 25844 4464 25900
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4728 25844 4756 25900
rect 4436 24332 4756 25844
rect 4436 24276 4464 24332
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4728 24276 4756 24332
rect 4436 22764 4756 24276
rect 5292 27076 5348 27086
rect 5292 23604 5348 27020
rect 5404 26964 5460 26974
rect 5404 25060 5460 26908
rect 5404 24994 5460 25004
rect 5292 23538 5348 23548
rect 4436 22708 4464 22764
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4728 22708 4756 22764
rect 4436 21196 4756 22708
rect 4436 21140 4464 21196
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4728 21140 4756 21196
rect 4436 19628 4756 21140
rect 4436 19572 4464 19628
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4728 19572 4756 19628
rect 4436 18060 4756 19572
rect 4436 18004 4464 18060
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4728 18004 4756 18060
rect 3776 15652 3804 15708
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 4068 15652 4096 15708
rect 3776 14140 4096 15652
rect 3776 14084 3804 14140
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 4068 14084 4096 14140
rect 3776 12572 4096 14084
rect 3776 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4096 12572
rect 3776 11004 4096 12516
rect 3776 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4096 11004
rect 3776 9436 4096 10948
rect 3776 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4096 9436
rect 3776 7868 4096 9380
rect 3776 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4096 7868
rect 3776 6300 4096 7812
rect 3776 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4096 6300
rect 3776 4732 4096 6244
rect 3776 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4096 4732
rect 3776 3164 4096 4676
rect 3776 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4096 3164
rect 3776 1596 4096 3108
rect 3776 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4096 1596
rect 3776 0 4096 1540
rect 4436 16492 4756 18004
rect 4436 16436 4464 16492
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4728 16436 4756 16492
rect 4436 14924 4756 16436
rect 4436 14868 4464 14924
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4728 14868 4756 14924
rect 4436 13356 4756 14868
rect 4436 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4756 13356
rect 4436 11788 4756 13300
rect 4956 16548 5012 16558
rect 4956 12516 5012 16492
rect 4956 12450 5012 12460
rect 4436 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4756 11788
rect 4436 10220 4756 11732
rect 4436 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4756 10220
rect 4436 8652 4756 10164
rect 5516 9156 5572 41468
rect 6188 26404 6244 26414
rect 6188 26180 6244 26348
rect 6188 26114 6244 26124
rect 6300 18676 6356 48972
rect 7308 39844 7364 39854
rect 6748 33460 6804 33470
rect 6748 26068 6804 33404
rect 6748 26002 6804 26012
rect 6300 18610 6356 18620
rect 5516 9090 5572 9100
rect 6412 13524 6468 13534
rect 6412 9156 6468 13468
rect 6412 9090 6468 9100
rect 4436 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4756 8652
rect 4436 7084 4756 8596
rect 7308 7700 7364 39788
rect 8428 39620 8484 39630
rect 7420 31668 7476 31678
rect 7420 29316 7476 31612
rect 7420 29250 7476 29260
rect 7980 28308 8036 28318
rect 7980 26964 8036 28252
rect 7980 24500 8036 26908
rect 7980 24434 8036 24444
rect 8316 14420 8372 14430
rect 8316 13188 8372 14364
rect 8316 13122 8372 13132
rect 7308 7634 7364 7644
rect 4436 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4756 7084
rect 4436 5516 4756 7028
rect 4436 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4756 5516
rect 4436 3948 4756 5460
rect 4436 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4756 3948
rect 4436 2380 4756 3892
rect 4436 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4756 2380
rect 4436 812 4756 2324
rect 4436 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4756 812
rect 4436 0 4756 756
rect 8428 420 8484 39564
rect 8876 34468 8932 34478
rect 8764 29316 8820 29326
rect 8540 21140 8596 21150
rect 8540 14756 8596 21084
rect 8540 13524 8596 14700
rect 8540 13458 8596 13468
rect 8764 10724 8820 29260
rect 8876 28756 8932 34412
rect 8876 28690 8932 28700
rect 9212 14196 9268 49644
rect 9884 35364 9940 35374
rect 9660 34020 9716 34030
rect 9660 31892 9716 33964
rect 9660 25060 9716 31836
rect 9660 24994 9716 25004
rect 9884 19348 9940 35308
rect 10444 35252 10500 35262
rect 10220 32900 10276 32910
rect 10108 27300 10164 27310
rect 10108 26068 10164 27244
rect 10108 26002 10164 26012
rect 10220 25508 10276 32844
rect 10220 25442 10276 25452
rect 10220 24052 10276 24062
rect 9884 19282 9940 19292
rect 9996 21252 10052 21262
rect 9212 14130 9268 14140
rect 9996 16884 10052 21196
rect 10220 18340 10276 23996
rect 10220 18274 10276 18284
rect 9996 13076 10052 16828
rect 10444 16212 10500 35196
rect 10668 31668 10724 31678
rect 10668 28084 10724 31612
rect 10668 28018 10724 28028
rect 10444 16146 10500 16156
rect 9996 13010 10052 13020
rect 9100 12180 9156 12190
rect 9100 11060 9156 12124
rect 10780 11172 10836 50652
rect 11228 41860 11284 41870
rect 10780 11106 10836 11116
rect 10892 34916 10948 34926
rect 9100 10994 9156 11004
rect 8764 10658 8820 10668
rect 10892 644 10948 34860
rect 11004 30436 11060 30446
rect 11004 29428 11060 30380
rect 11004 29362 11060 29372
rect 11004 29204 11060 29214
rect 11004 23828 11060 29148
rect 11228 27300 11284 41804
rect 11676 33012 11732 33022
rect 11676 28532 11732 32956
rect 11676 28466 11732 28476
rect 11228 27234 11284 27244
rect 11004 23762 11060 23772
rect 12012 21924 12068 21934
rect 11676 13412 11732 13422
rect 11676 11172 11732 13356
rect 12012 12516 12068 21868
rect 12572 13524 12628 53900
rect 20860 52164 20916 52174
rect 14140 51156 14196 51166
rect 14028 34468 14084 34478
rect 13244 32564 13300 32574
rect 13132 31892 13188 31902
rect 13132 26740 13188 31836
rect 13244 31332 13300 32508
rect 13244 31266 13300 31276
rect 13468 32116 13524 32126
rect 13468 27188 13524 32060
rect 13468 27122 13524 27132
rect 13692 30772 13748 30782
rect 13132 26674 13188 26684
rect 13692 24948 13748 30716
rect 14028 26740 14084 34412
rect 14028 26674 14084 26684
rect 13692 24882 13748 24892
rect 14140 23044 14196 51100
rect 18396 50596 18452 50606
rect 16268 49252 16324 49262
rect 14140 22978 14196 22988
rect 14812 48916 14868 48926
rect 13468 20356 13524 20366
rect 13132 20020 13188 20030
rect 12908 19012 12964 19022
rect 12908 18340 12964 18956
rect 13132 18788 13188 19964
rect 13132 18722 13188 18732
rect 13356 19684 13412 19694
rect 12908 18274 12964 18284
rect 13356 18340 13412 19628
rect 12572 13458 12628 13468
rect 12796 13524 12852 13534
rect 12012 12450 12068 12460
rect 12796 12516 12852 13468
rect 13356 13412 13412 18284
rect 13468 15876 13524 20300
rect 13804 16772 13860 16782
rect 13804 16324 13860 16716
rect 13804 16258 13860 16268
rect 13468 15810 13524 15820
rect 13356 13346 13412 13356
rect 12796 12450 12852 12460
rect 12460 12292 12516 12302
rect 12460 11956 12516 12236
rect 12460 11890 12516 11900
rect 11676 11106 11732 11116
rect 12012 11060 12068 11070
rect 12012 10500 12068 11004
rect 12012 10434 12068 10444
rect 14812 7140 14868 48860
rect 16044 28420 16100 28430
rect 15932 26852 15988 26862
rect 15932 25956 15988 26796
rect 15932 25890 15988 25900
rect 14924 17332 14980 17342
rect 14924 16996 14980 17276
rect 14924 16930 14980 16940
rect 15372 14868 15428 14878
rect 15372 14196 15428 14812
rect 15372 14130 15428 14140
rect 15596 14196 15652 14206
rect 15596 12964 15652 14140
rect 15596 12898 15652 12908
rect 14812 7074 14868 7084
rect 16044 1316 16100 28364
rect 16268 23604 16324 49196
rect 16268 23538 16324 23548
rect 16716 48132 16772 48142
rect 16716 1652 16772 48076
rect 17836 13076 17892 13086
rect 17164 12740 17220 12750
rect 17164 11284 17220 12684
rect 17836 11844 17892 13020
rect 18060 12852 18116 12862
rect 17836 11778 17892 11788
rect 17948 12740 18004 12750
rect 17948 12404 18004 12684
rect 17164 11218 17220 11228
rect 17948 11060 18004 12348
rect 18060 11844 18116 12796
rect 18060 11778 18116 11788
rect 17948 10994 18004 11004
rect 16716 1586 16772 1596
rect 16044 1250 16100 1260
rect 10892 578 10948 588
rect 8428 354 8484 364
rect 18396 420 18452 50540
rect 19292 47460 19348 47470
rect 18620 23044 18676 23054
rect 18620 18564 18676 22988
rect 18620 18498 18676 18508
rect 18732 20020 18788 20030
rect 18732 16100 18788 19964
rect 18732 16034 18788 16044
rect 18844 18228 18900 18238
rect 18844 4228 18900 18172
rect 19068 18116 19124 18126
rect 19068 16548 19124 18060
rect 19068 16482 19124 16492
rect 18956 16436 19012 16446
rect 18956 16100 19012 16380
rect 18956 16034 19012 16044
rect 19180 13076 19236 13086
rect 19180 11844 19236 13020
rect 19180 11778 19236 11788
rect 19292 6692 19348 47404
rect 20636 23940 20692 23950
rect 20076 23156 20132 23166
rect 19516 22148 19572 22158
rect 19516 17668 19572 22092
rect 19964 22148 20020 22158
rect 19964 21140 20020 22092
rect 19964 21074 20020 21084
rect 20076 20020 20132 23100
rect 20636 22932 20692 23884
rect 20636 22866 20692 22876
rect 20076 19954 20132 19964
rect 19404 17444 19460 17454
rect 19404 16436 19460 17388
rect 19404 16370 19460 16380
rect 19516 11956 19572 17612
rect 19628 17220 19684 17230
rect 19628 16436 19684 17164
rect 19628 16370 19684 16380
rect 19628 15876 19684 15886
rect 19628 15428 19684 15820
rect 19628 15362 19684 15372
rect 19852 15428 19908 15438
rect 19852 14868 19908 15372
rect 19852 14644 19908 14812
rect 19852 14578 19908 14588
rect 19516 11890 19572 11900
rect 19292 6626 19348 6636
rect 18844 4162 18900 4172
rect 20860 1652 20916 52108
rect 21308 6692 21364 55916
rect 22428 55300 22484 55310
rect 21756 54516 21812 54526
rect 21756 13636 21812 54460
rect 21756 13570 21812 13580
rect 21308 6626 21364 6636
rect 22428 6580 22484 55244
rect 23776 54908 24096 56420
rect 23776 54852 23804 54908
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 24068 54852 24096 54908
rect 23776 53340 24096 54852
rect 23776 53284 23804 53340
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 24068 53284 24096 53340
rect 22428 6514 22484 6524
rect 22764 52164 22820 52174
rect 22764 6468 22820 52108
rect 23776 51772 24096 53284
rect 23776 51716 23804 51772
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 24068 51716 24096 51772
rect 23776 50204 24096 51716
rect 23776 50148 23804 50204
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 24068 50148 24096 50204
rect 23776 48636 24096 50148
rect 23776 48580 23804 48636
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 24068 48580 24096 48636
rect 23776 47068 24096 48580
rect 23776 47012 23804 47068
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 24068 47012 24096 47068
rect 23776 45500 24096 47012
rect 23776 45444 23804 45500
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 24068 45444 24096 45500
rect 23776 43932 24096 45444
rect 23776 43876 23804 43932
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 24068 43876 24096 43932
rect 23776 42364 24096 43876
rect 23776 42308 23804 42364
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 24068 42308 24096 42364
rect 23776 40796 24096 42308
rect 23776 40740 23804 40796
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 24068 40740 24096 40796
rect 23776 39228 24096 40740
rect 23776 39172 23804 39228
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 24068 39172 24096 39228
rect 23776 37660 24096 39172
rect 23776 37604 23804 37660
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 24068 37604 24096 37660
rect 23776 36092 24096 37604
rect 23776 36036 23804 36092
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 24068 36036 24096 36092
rect 23776 34524 24096 36036
rect 23776 34468 23804 34524
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 24068 34468 24096 34524
rect 23776 32956 24096 34468
rect 23776 32900 23804 32956
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 24068 32900 24096 32956
rect 23776 31388 24096 32900
rect 23776 31332 23804 31388
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 24068 31332 24096 31388
rect 23548 30100 23604 30110
rect 23548 21588 23604 30044
rect 23548 21522 23604 21532
rect 23776 29820 24096 31332
rect 23776 29764 23804 29820
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 24068 29764 24096 29820
rect 23776 28252 24096 29764
rect 23776 28196 23804 28252
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 24068 28196 24096 28252
rect 23776 26684 24096 28196
rect 23776 26628 23804 26684
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 24068 26628 24096 26684
rect 23776 25116 24096 26628
rect 23776 25060 23804 25116
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 24068 25060 24096 25116
rect 23776 23548 24096 25060
rect 23776 23492 23804 23548
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 24068 23492 24096 23548
rect 23776 21980 24096 23492
rect 23776 21924 23804 21980
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 24068 21924 24096 21980
rect 22764 6402 22820 6412
rect 23776 20412 24096 21924
rect 23776 20356 23804 20412
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 24068 20356 24096 20412
rect 23776 18844 24096 20356
rect 23776 18788 23804 18844
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 24068 18788 24096 18844
rect 23776 17276 24096 18788
rect 23776 17220 23804 17276
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 24068 17220 24096 17276
rect 23776 15708 24096 17220
rect 23776 15652 23804 15708
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 24068 15652 24096 15708
rect 23776 14140 24096 15652
rect 23776 14084 23804 14140
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 24068 14084 24096 14140
rect 23776 12572 24096 14084
rect 23776 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24096 12572
rect 23776 11004 24096 12516
rect 23776 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24096 11004
rect 23776 9436 24096 10948
rect 23776 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24096 9436
rect 23776 7868 24096 9380
rect 23776 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24096 7868
rect 20860 1586 20916 1596
rect 23776 6300 24096 7812
rect 23776 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24096 6300
rect 23776 4732 24096 6244
rect 23776 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24096 4732
rect 23776 3164 24096 4676
rect 23776 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24096 3164
rect 23776 1596 24096 3108
rect 18396 354 18452 364
rect 23776 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24096 1596
rect 23776 0 24096 1540
rect 24436 55692 24756 57456
rect 24436 55636 24464 55692
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24728 55636 24756 55692
rect 24436 54124 24756 55636
rect 24436 54068 24464 54124
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24728 54068 24756 54124
rect 24436 52556 24756 54068
rect 24436 52500 24464 52556
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24728 52500 24756 52556
rect 24436 50988 24756 52500
rect 24436 50932 24464 50988
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24728 50932 24756 50988
rect 24436 49420 24756 50932
rect 24436 49364 24464 49420
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24728 49364 24756 49420
rect 24436 47852 24756 49364
rect 24436 47796 24464 47852
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24728 47796 24756 47852
rect 24436 46284 24756 47796
rect 24436 46228 24464 46284
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24728 46228 24756 46284
rect 24436 44716 24756 46228
rect 24436 44660 24464 44716
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24728 44660 24756 44716
rect 24436 43148 24756 44660
rect 24436 43092 24464 43148
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24728 43092 24756 43148
rect 24436 41580 24756 43092
rect 24436 41524 24464 41580
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24728 41524 24756 41580
rect 24436 40012 24756 41524
rect 24436 39956 24464 40012
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24728 39956 24756 40012
rect 24436 38444 24756 39956
rect 24436 38388 24464 38444
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24728 38388 24756 38444
rect 24436 36876 24756 38388
rect 24436 36820 24464 36876
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24728 36820 24756 36876
rect 24436 35308 24756 36820
rect 24436 35252 24464 35308
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24728 35252 24756 35308
rect 24436 33740 24756 35252
rect 24436 33684 24464 33740
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24728 33684 24756 33740
rect 24436 32172 24756 33684
rect 24436 32116 24464 32172
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24728 32116 24756 32172
rect 24436 30604 24756 32116
rect 24436 30548 24464 30604
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24728 30548 24756 30604
rect 24436 29036 24756 30548
rect 24436 28980 24464 29036
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24728 28980 24756 29036
rect 24436 27468 24756 28980
rect 24436 27412 24464 27468
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24728 27412 24756 27468
rect 24436 25900 24756 27412
rect 26124 55300 26180 55310
rect 24436 25844 24464 25900
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24728 25844 24756 25900
rect 24436 24332 24756 25844
rect 24436 24276 24464 24332
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24728 24276 24756 24332
rect 24436 22764 24756 24276
rect 24436 22708 24464 22764
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24728 22708 24756 22764
rect 24436 21196 24756 22708
rect 24436 21140 24464 21196
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24728 21140 24756 21196
rect 24436 19628 24756 21140
rect 25228 26180 25284 26190
rect 25228 20692 25284 26124
rect 25228 20626 25284 20636
rect 25900 20804 25956 20814
rect 24436 19572 24464 19628
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24728 19572 24756 19628
rect 24436 18060 24756 19572
rect 24436 18004 24464 18060
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24728 18004 24756 18060
rect 24436 16492 24756 18004
rect 24436 16436 24464 16492
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24728 16436 24756 16492
rect 24436 14924 24756 16436
rect 24436 14868 24464 14924
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24728 14868 24756 14924
rect 24436 13356 24756 14868
rect 24436 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24756 13356
rect 24436 11788 24756 13300
rect 25900 11956 25956 20748
rect 26012 17108 26068 17118
rect 26012 12180 26068 17052
rect 26012 12114 26068 12124
rect 25900 11890 25956 11900
rect 24436 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24756 11788
rect 24436 10220 24756 11732
rect 24436 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24756 10220
rect 24436 8652 24756 10164
rect 24436 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24756 8652
rect 24436 7084 24756 8596
rect 26124 8036 26180 55244
rect 27020 50820 27076 50830
rect 26908 39732 26964 39742
rect 26348 31444 26404 31454
rect 26348 29316 26404 31388
rect 26348 29250 26404 29260
rect 26236 27748 26292 27758
rect 26236 24836 26292 27692
rect 26236 24770 26292 24780
rect 26908 19348 26964 39676
rect 26908 19282 26964 19292
rect 26908 16772 26964 16782
rect 26908 11508 26964 16716
rect 26908 11442 26964 11452
rect 26124 7970 26180 7980
rect 24436 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24756 7084
rect 24436 5516 24756 7028
rect 24436 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24756 5516
rect 24436 3948 24756 5460
rect 24436 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24756 3948
rect 24436 2380 24756 3892
rect 24436 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24756 2380
rect 24436 812 24756 2324
rect 27020 1092 27076 50764
rect 27132 21476 27188 21486
rect 27132 13860 27188 21420
rect 27132 13794 27188 13804
rect 27468 7924 27524 7934
rect 27468 7364 27524 7868
rect 27468 7298 27524 7308
rect 27020 1026 27076 1036
rect 24436 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24756 812
rect 24436 0 24756 756
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _078_
timestamp 1486834041
transform 1 0 15904 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _079_
timestamp 1486834041
transform -1 0 10080 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _080_
timestamp 1486834041
transform -1 0 17584 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _081_
timestamp 1486834041
transform -1 0 16352 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _082_
timestamp 1486834041
transform 1 0 14784 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _083_
timestamp 1486834041
transform 1 0 3360 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _084_
timestamp 1486834041
transform 1 0 11984 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _085_
timestamp 1486834041
transform 1 0 8064 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _086_
timestamp 1486834041
transform -1 0 21840 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _087_
timestamp 1486834041
transform 1 0 16576 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _088_
timestamp 1486834041
transform 1 0 15904 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _089_
timestamp 1486834041
transform -1 0 20272 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _090_
timestamp 1486834041
transform 1 0 6832 0 1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _091_
timestamp 1486834041
transform 1 0 4928 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _092_
timestamp 1486834041
transform 1 0 4928 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _093_
timestamp 1486834041
transform 1 0 13440 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _094_
timestamp 1486834041
transform 1 0 11088 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _095_
timestamp 1486834041
transform 1 0 18144 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _096_
timestamp 1486834041
transform 1 0 11312 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _097_
timestamp 1486834041
transform 1 0 15232 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _098_
timestamp 1486834041
transform 1 0 14784 0 -1 10192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _099_
timestamp 1486834041
transform 1 0 15232 0 -1 8624
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _100_
timestamp 1486834041
transform 1 0 16016 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _101_
timestamp 1486834041
transform -1 0 17472 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _102_
timestamp 1486834041
transform 1 0 15456 0 1 7056
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _103_
timestamp 1486834041
transform 1 0 16576 0 1 10192
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _104_
timestamp 1486834041
transform 1 0 16576 0 -1 8624
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _105_
timestamp 1486834041
transform 1 0 8736 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _106_
timestamp 1486834041
transform 1 0 6944 0 -1 11760
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _107_
timestamp 1486834041
transform 1 0 3808 0 -1 14896
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _108_
timestamp 1486834041
transform 1 0 7616 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _109_
timestamp 1486834041
transform -1 0 7952 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _110_
timestamp 1486834041
transform 1 0 5712 0 -1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _111_
timestamp 1486834041
transform -1 0 9520 0 -1 14896
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _112_
timestamp 1486834041
transform 1 0 7168 0 -1 14896
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _113_
timestamp 1486834041
transform -1 0 13328 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _114_
timestamp 1486834041
transform 1 0 11312 0 1 10192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _115_
timestamp 1486834041
transform -1 0 13664 0 -1 10192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _116_
timestamp 1486834041
transform 1 0 13664 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _117_
timestamp 1486834041
transform 1 0 11312 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _118_
timestamp 1486834041
transform -1 0 11312 0 -1 11760
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _119_
timestamp 1486834041
transform 1 0 10528 0 1 10192
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _120_
timestamp 1486834041
transform 1 0 12656 0 1 10192
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _121_
timestamp 1486834041
transform -1 0 9408 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _122_
timestamp 1486834041
transform 1 0 6944 0 -1 10192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _123_
timestamp 1486834041
transform -1 0 9072 0 1 11760
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _124_
timestamp 1486834041
transform 1 0 8736 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _125_
timestamp 1486834041
transform -1 0 7728 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _126_
timestamp 1486834041
transform 1 0 7952 0 -1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _127_
timestamp 1486834041
transform -1 0 10304 0 1 10192
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _128_
timestamp 1486834041
transform 1 0 7056 0 1 10192
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _129_
timestamp 1486834041
transform 1 0 19376 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _130_
timestamp 1486834041
transform 1 0 20496 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _131_
timestamp 1486834041
transform 1 0 19040 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _132_
timestamp 1486834041
transform 1 0 20496 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _133_
timestamp 1486834041
transform 1 0 20496 0 1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _134_
timestamp 1486834041
transform -1 0 20272 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _135_
timestamp 1486834041
transform 1 0 17136 0 1 13328
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _136_
timestamp 1486834041
transform -1 0 21168 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _137_
timestamp 1486834041
transform 1 0 17696 0 -1 16464
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _138_
timestamp 1486834041
transform 1 0 16576 0 -1 16464
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _139_
timestamp 1486834041
transform 1 0 18928 0 1 13328
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _140_
timestamp 1486834041
transform 1 0 20496 0 1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _141_
timestamp 1486834041
transform -1 0 20160 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _142_
timestamp 1486834041
transform 1 0 18816 0 -1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _143_
timestamp 1486834041
transform -1 0 19936 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _144_
timestamp 1486834041
transform -1 0 19040 0 1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _145_
timestamp 1486834041
transform 1 0 18480 0 1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _146_
timestamp 1486834041
transform 1 0 17696 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _147_
timestamp 1486834041
transform -1 0 17696 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _148_
timestamp 1486834041
transform 1 0 18144 0 1 16464
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _149_
timestamp 1486834041
transform 1 0 17808 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _150_
timestamp 1486834041
transform -1 0 18032 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _151_
timestamp 1486834041
transform 1 0 17584 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _152_
timestamp 1486834041
transform 1 0 19264 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _153_
timestamp 1486834041
transform 1 0 17584 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _154_
timestamp 1486834041
transform -1 0 18928 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _155_
timestamp 1486834041
transform 1 0 16576 0 -1 13328
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _156_
timestamp 1486834041
transform 1 0 16576 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _157_
timestamp 1486834041
transform -1 0 19376 0 1 14896
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _158_
timestamp 1486834041
transform 1 0 16800 0 1 11760
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _159_
timestamp 1486834041
transform 1 0 17920 0 1 11760
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _160_
timestamp 1486834041
transform 1 0 19152 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _161_
timestamp 1486834041
transform 1 0 20496 0 1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _162_
timestamp 1486834041
transform 1 0 18592 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _163_
timestamp 1486834041
transform -1 0 20272 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _164_
timestamp 1486834041
transform -1 0 21504 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _165_
timestamp 1486834041
transform -1 0 20272 0 1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _166_
timestamp 1486834041
transform -1 0 18256 0 -1 21168
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _167_
timestamp 1486834041
transform -1 0 18704 0 1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _168_
timestamp 1486834041
transform 1 0 16800 0 -1 19600
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _169_
timestamp 1486834041
transform 1 0 18704 0 1 21168
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _170_
timestamp 1486834041
transform 1 0 20496 0 1 21168
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _171_
timestamp 1486834041
transform 1 0 15008 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _172_
timestamp 1486834041
transform 1 0 8624 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _173_
timestamp 1486834041
transform 1 0 12432 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _174_
timestamp 1486834041
transform 1 0 2016 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _175_
timestamp 1486834041
transform 1 0 14448 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _176_
timestamp 1486834041
transform 1 0 8848 0 1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _177_
timestamp 1486834041
transform 1 0 19264 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _178_
timestamp 1486834041
transform -1 0 12432 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _179_
timestamp 1486834041
transform 1 0 20496 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _180_
timestamp 1486834041
transform 1 0 2240 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _181_
timestamp 1486834041
transform 1 0 15344 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _182_
timestamp 1486834041
transform 1 0 3360 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _183_
timestamp 1486834041
transform 1 0 12320 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _184_
timestamp 1486834041
transform 1 0 14560 0 1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _185_
timestamp 1486834041
transform 1 0 20496 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _186_
timestamp 1486834041
transform 1 0 7840 0 1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _187_
timestamp 1486834041
transform 1 0 2688 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _188_
timestamp 1486834041
transform 1 0 6832 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _189_
timestamp 1486834041
transform 1 0 4928 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _190_
timestamp 1486834041
transform 1 0 2128 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _191_
timestamp 1486834041
transform 1 0 12656 0 1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _192_
timestamp 1486834041
transform 1 0 14560 0 1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _193_
timestamp 1486834041
transform 1 0 10192 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _194_
timestamp 1486834041
transform 1 0 8848 0 1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _195_
timestamp 1486834041
transform 1 0 20048 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _196_
timestamp 1486834041
transform 1 0 5936 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _197_
timestamp 1486834041
transform 1 0 1008 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _198_
timestamp 1486834041
transform 1 0 2464 0 -1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _199_
timestamp 1486834041
transform 1 0 13664 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _200_
timestamp 1486834041
transform 1 0 8960 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _201_
timestamp 1486834041
transform 1 0 17248 0 -1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _202_
timestamp 1486834041
transform 1 0 12656 0 1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _203_
timestamp 1486834041
transform 1 0 14224 0 1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _204_
timestamp 1486834041
transform -1 0 8736 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _205_
timestamp 1486834041
transform -1 0 4928 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _206_
timestamp 1486834041
transform 1 0 3136 0 -1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _207_
timestamp 1486834041
transform 1 0 13552 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _208_
timestamp 1486834041
transform 1 0 8848 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _209_
timestamp 1486834041
transform 1 0 16576 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _210_
timestamp 1486834041
transform 1 0 11424 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _211_
timestamp 1486834041
transform 1 0 14336 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _212_
timestamp 1486834041
transform -1 0 8848 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _213_
timestamp 1486834041
transform -1 0 7056 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _214_
timestamp 1486834041
transform -1 0 25648 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _215_
timestamp 1486834041
transform -1 0 19040 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _216_
timestamp 1486834041
transform -1 0 9744 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _217_
timestamp 1486834041
transform -1 0 24528 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _218_
timestamp 1486834041
transform 1 0 24416 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _219_
timestamp 1486834041
transform -1 0 24192 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _220_
timestamp 1486834041
transform 1 0 1456 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _221_
timestamp 1486834041
transform 1 0 1680 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _222_
timestamp 1486834041
transform -1 0 3584 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _223_
timestamp 1486834041
transform 1 0 1680 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _224_
timestamp 1486834041
transform -1 0 8512 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _225_
timestamp 1486834041
transform -1 0 8624 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _226_
timestamp 1486834041
transform 1 0 1904 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _227_
timestamp 1486834041
transform -1 0 7280 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _228_
timestamp 1486834041
transform 1 0 10080 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _229_
timestamp 1486834041
transform 1 0 9520 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _230_
timestamp 1486834041
transform 1 0 17024 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _231_
timestamp 1486834041
transform 1 0 17472 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _232_
timestamp 1486834041
transform 1 0 5712 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _233_
timestamp 1486834041
transform 1 0 10976 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _234_
timestamp 1486834041
transform 1 0 11200 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _235_
timestamp 1486834041
transform 1 0 13440 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _236_
timestamp 1486834041
transform 1 0 2688 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _237_
timestamp 1486834041
transform -1 0 7840 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _238_
timestamp 1486834041
transform 1 0 3248 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _239_
timestamp 1486834041
transform 1 0 2352 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _240_
timestamp 1486834041
transform 1 0 2352 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _241_
timestamp 1486834041
transform 1 0 5264 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _242_
timestamp 1486834041
transform 1 0 10192 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _243_
timestamp 1486834041
transform -1 0 18816 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _244_
timestamp 1486834041
transform 1 0 9184 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _245_
timestamp 1486834041
transform 1 0 10192 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _246_
timestamp 1486834041
transform 1 0 14336 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _247_
timestamp 1486834041
transform 1 0 11424 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _248_
timestamp 1486834041
transform 1 0 6608 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _249_
timestamp 1486834041
transform 1 0 9072 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _250_
timestamp 1486834041
transform 1 0 12208 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _251_
timestamp 1486834041
transform 1 0 11872 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _252_
timestamp 1486834041
transform 1 0 2016 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _253_
timestamp 1486834041
transform 1 0 1680 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _254_
timestamp 1486834041
transform 1 0 1344 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _255_
timestamp 1486834041
transform 1 0 1008 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _256_
timestamp 1486834041
transform 1 0 5824 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _257_
timestamp 1486834041
transform -1 0 9744 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _258_
timestamp 1486834041
transform 1 0 12768 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _259_
timestamp 1486834041
transform 1 0 13888 0 1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _260_
timestamp 1486834041
transform 1 0 6272 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _261_
timestamp 1486834041
transform 1 0 10192 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _262_
timestamp 1486834041
transform 1 0 16688 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _263_
timestamp 1486834041
transform 1 0 17024 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _264_
timestamp 1486834041
transform 1 0 7728 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _265_
timestamp 1486834041
transform 1 0 8960 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _266_
timestamp 1486834041
transform 1 0 12544 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _267_
timestamp 1486834041
transform 1 0 12992 0 -1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _268_
timestamp 1486834041
transform 1 0 896 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _269_
timestamp 1486834041
transform 1 0 1568 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _270_
timestamp 1486834041
transform -1 0 3136 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _271_
timestamp 1486834041
transform 1 0 1008 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _272_
timestamp 1486834041
transform 1 0 4032 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _273_
timestamp 1486834041
transform 1 0 5040 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _274_
timestamp 1486834041
transform 1 0 18928 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _275_
timestamp 1486834041
transform 1 0 21168 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _276_
timestamp 1486834041
transform -1 0 10976 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _277_
timestamp 1486834041
transform 1 0 8736 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _278_
timestamp 1486834041
transform 1 0 9184 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _279_
timestamp 1486834041
transform 1 0 10080 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _280_
timestamp 1486834041
transform 1 0 10528 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _281_
timestamp 1486834041
transform 1 0 13104 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _282_
timestamp 1486834041
transform 1 0 12656 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _283_
timestamp 1486834041
transform 1 0 10192 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _284_
timestamp 1486834041
transform 1 0 896 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _285_
timestamp 1486834041
transform 1 0 1344 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _286_
timestamp 1486834041
transform 1 0 5264 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _287_
timestamp 1486834041
transform 1 0 2352 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _288_
timestamp 1486834041
transform 1 0 6048 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _289_
timestamp 1486834041
transform 1 0 6272 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _290_
timestamp 1486834041
transform -1 0 5040 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _291_
timestamp 1486834041
transform 1 0 2352 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _292_
timestamp 1486834041
transform 1 0 6160 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _293_
timestamp 1486834041
transform -1 0 10976 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _294_
timestamp 1486834041
transform 1 0 18032 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _295_
timestamp 1486834041
transform 1 0 17808 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _296_
timestamp 1486834041
transform 1 0 10864 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _297_
timestamp 1486834041
transform 1 0 9632 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _298_
timestamp 1486834041
transform 1 0 11872 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _299_
timestamp 1486834041
transform 1 0 10080 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _300_
timestamp 1486834041
transform 1 0 2352 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _301_
timestamp 1486834041
transform 1 0 1680 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _302_
timestamp 1486834041
transform 1 0 13104 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _303_
timestamp 1486834041
transform 1 0 6944 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _304_
timestamp 1486834041
transform 1 0 896 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _305_
timestamp 1486834041
transform 1 0 1904 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _306_
timestamp 1486834041
transform 1 0 20160 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _307_
timestamp 1486834041
transform 1 0 20496 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _308_
timestamp 1486834041
transform 1 0 8176 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _309_
timestamp 1486834041
transform 1 0 7840 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _310_
timestamp 1486834041
transform 1 0 19376 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _311_
timestamp 1486834041
transform 1 0 18032 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _312_
timestamp 1486834041
transform 1 0 7952 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _313_
timestamp 1486834041
transform 1 0 6272 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _314_
timestamp 1486834041
transform 1 0 14112 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _315_
timestamp 1486834041
transform 1 0 12880 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _316_
timestamp 1486834041
transform 1 0 896 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _317_
timestamp 1486834041
transform 1 0 1344 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _318_
timestamp 1486834041
transform 1 0 6608 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _319_
timestamp 1486834041
transform 1 0 10192 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _320_
timestamp 1486834041
transform 1 0 6160 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _321_
timestamp 1486834041
transform 1 0 6272 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _322_
timestamp 1486834041
transform 1 0 14112 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _323_
timestamp 1486834041
transform 1 0 13552 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _324_
timestamp 1486834041
transform 1 0 14112 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _325_
timestamp 1486834041
transform 1 0 14112 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _326_
timestamp 1486834041
transform 1 0 17808 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _327_
timestamp 1486834041
transform 1 0 17808 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _328_
timestamp 1486834041
transform 1 0 14560 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _329_
timestamp 1486834041
transform 1 0 11984 0 -1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _330_
timestamp 1486834041
transform 1 0 12656 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _331_
timestamp 1486834041
transform 1 0 14336 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _332_
timestamp 1486834041
transform 1 0 12768 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _333_
timestamp 1486834041
transform 1 0 14112 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _334_
timestamp 1486834041
transform 1 0 14560 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _335_
timestamp 1486834041
transform 1 0 4928 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _336_
timestamp 1486834041
transform -1 0 4592 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _337_
timestamp 1486834041
transform 1 0 4816 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _338_
timestamp 1486834041
transform 1 0 16240 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _339_
timestamp 1486834041
transform -1 0 23520 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _340_
timestamp 1486834041
transform 1 0 7952 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _341_
timestamp 1486834041
transform 1 0 10192 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _342_
timestamp 1486834041
transform 1 0 9632 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _343_
timestamp 1486834041
transform 1 0 10192 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _344_
timestamp 1486834041
transform 1 0 10304 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _345_
timestamp 1486834041
transform -1 0 23408 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _346_
timestamp 1486834041
transform -1 0 20272 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _347_
timestamp 1486834041
transform -1 0 23408 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _348_
timestamp 1486834041
transform 1 0 3808 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _349_
timestamp 1486834041
transform 1 0 4816 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _350_
timestamp 1486834041
transform 1 0 4704 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _351_
timestamp 1486834041
transform 1 0 4592 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _352_
timestamp 1486834041
transform 1 0 12320 0 -1 33712
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _353_
timestamp 1486834041
transform 1 0 8400 0 1 36848
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _354_
timestamp 1486834041
transform 1 0 12656 0 1 33712
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _355_
timestamp 1486834041
transform 1 0 8400 0 1 35280
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _356_
timestamp 1486834041
transform -1 0 11312 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _357_
timestamp 1486834041
transform 1 0 19376 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _358_
timestamp 1486834041
transform 1 0 12656 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _359_
timestamp 1486834041
transform 1 0 15120 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _360_
timestamp 1486834041
transform -1 0 5712 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _361_
timestamp 1486834041
transform 1 0 8736 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _362_
timestamp 1486834041
transform 1 0 8736 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _363_
timestamp 1486834041
transform 1 0 15344 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _364_
timestamp 1486834041
transform -1 0 12432 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _365_
timestamp 1486834041
transform 1 0 18032 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _366_
timestamp 1486834041
transform 1 0 9632 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _367_
timestamp 1486834041
transform 1 0 15008 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _368_
timestamp 1486834041
transform 1 0 4816 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _369_
timestamp 1486834041
transform 1 0 3136 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _370_
timestamp 1486834041
transform -1 0 5936 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _371_
timestamp 1486834041
transform 1 0 15344 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _372_
timestamp 1486834041
transform -1 0 13552 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _373_
timestamp 1486834041
transform 1 0 18480 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _374_
timestamp 1486834041
transform -1 0 10416 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _375_
timestamp 1486834041
transform 1 0 15232 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _376_
timestamp 1486834041
transform 1 0 4816 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _377_
timestamp 1486834041
transform 1 0 16576 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _378_
timestamp 1486834041
transform -1 0 1904 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _379_
timestamp 1486834041
transform 1 0 21616 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _380_
timestamp 1486834041
transform -1 0 10416 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _381_
timestamp 1486834041
transform 1 0 20496 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _382_
timestamp 1486834041
transform 1 0 9744 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _383_
timestamp 1486834041
transform 1 0 16576 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _384_
timestamp 1486834041
transform -1 0 2016 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _385_
timestamp 1486834041
transform 1 0 13328 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _386_
timestamp 1486834041
transform 1 0 9408 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _387_
timestamp 1486834041
transform 1 0 16576 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _388_
timestamp 1486834041
transform 1 0 4816 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _389_
timestamp 1486834041
transform -1 0 2352 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _390_
timestamp 1486834041
transform -1 0 7168 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _391_
timestamp 1486834041
transform 1 0 21392 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _392_
timestamp 1486834041
transform 1 0 10416 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _393_
timestamp 1486834041
transform -1 0 11088 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _394_
timestamp 1486834041
transform 1 0 15344 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _395_
timestamp 1486834041
transform -1 0 14000 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _396_
timestamp 1486834041
transform 1 0 3136 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _397_
timestamp 1486834041
transform 1 0 5712 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _398_
timestamp 1486834041
transform 1 0 7616 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _399_
timestamp 1486834041
transform -1 0 2800 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _400_
timestamp 1486834041
transform 1 0 8848 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _401_
timestamp 1486834041
transform -1 0 21392 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _402_
timestamp 1486834041
transform -1 0 15904 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _403_
timestamp 1486834041
transform 1 0 13328 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _404_
timestamp 1486834041
transform 1 0 8736 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _405_
timestamp 1486834041
transform -1 0 6160 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _406_
timestamp 1486834041
transform 1 0 3696 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _407_
timestamp 1486834041
transform 1 0 11536 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _408_
timestamp 1486834041
transform 1 0 16240 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _409_
timestamp 1486834041
transform 1 0 15008 0 -1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _410_
timestamp 1486834041
transform 1 0 19040 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _411_
timestamp 1486834041
transform 1 0 17248 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _412_
timestamp 1486834041
transform 1 0 7056 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _413_
timestamp 1486834041
transform 1 0 10864 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _414_
timestamp 1486834041
transform 1 0 12096 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _415_
timestamp 1486834041
transform 1 0 11424 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _416_
timestamp 1486834041
transform 1 0 1456 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _417_
timestamp 1486834041
transform 1 0 3584 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _418_
timestamp 1486834041
transform 1 0 3696 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _419_
timestamp 1486834041
transform 1 0 1456 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _420_
timestamp 1486834041
transform 1 0 1792 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _421_
timestamp 1486834041
transform 1 0 2352 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _422_
timestamp 1486834041
transform 1 0 22400 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _423_
timestamp 1486834041
transform 1 0 22736 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _424_
timestamp 1486834041
transform 1 0 9184 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _425_
timestamp 1486834041
transform 1 0 6608 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _426_
timestamp 1486834041
transform 1 0 23296 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _427_
timestamp 1486834041
transform 1 0 17136 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _428_
timestamp 1486834041
transform 1 0 7616 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _429_
timestamp 1486834041
transform 1 0 23072 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _430_
timestamp 1486834041
transform -1 0 25312 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _431_
timestamp 1486834041
transform 1 0 11312 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _432_
timestamp 1486834041
transform 1 0 4816 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _433_
timestamp 1486834041
transform 1 0 2464 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _434_
timestamp 1486834041
transform 1 0 5712 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _435_
timestamp 1486834041
transform 1 0 2464 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _436_
timestamp 1486834041
transform -1 0 8064 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _437_
timestamp 1486834041
transform 1 0 2464 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _438_
timestamp 1486834041
transform -1 0 20608 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _439_
timestamp 1486834041
transform 1 0 1456 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _440_
timestamp 1486834041
transform -1 0 25312 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _441_
timestamp 1486834041
transform 1 0 25760 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _442_
timestamp 1486834041
transform 1 0 20496 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _443_
timestamp 1486834041
transform 1 0 25200 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _444_
timestamp 1486834041
transform 1 0 18928 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _445_
timestamp 1486834041
transform 1 0 25760 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _446_
timestamp 1486834041
transform 1 0 26656 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _447_
timestamp 1486834041
transform 1 0 19824 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _448_
timestamp 1486834041
transform 1 0 25872 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _449_
timestamp 1486834041
transform 1 0 26768 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _450_
timestamp 1486834041
transform 1 0 21280 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _451_
timestamp 1486834041
transform -1 0 14000 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _452_
timestamp 1486834041
transform -1 0 22624 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _453_
timestamp 1486834041
transform -1 0 24192 0 -1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _454_
timestamp 1486834041
transform -1 0 12208 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _455_
timestamp 1486834041
transform -1 0 4256 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _456_
timestamp 1486834041
transform -1 0 10752 0 -1 36848
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_UserCLK_regs
timestamp 1486834041
transform 1 0 12656 0 1 35280
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_UserCLK
timestamp 1486834041
transform 1 0 10752 0 -1 35280
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_UserCLK
timestamp 1486834041
transform -1 0 15344 0 -1 39984
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_UserCLK_regs
timestamp 1486834041
transform 1 0 13440 0 1 32144
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_UserCLK_regs
timestamp 1486834041
transform -1 0 14896 0 -1 38416
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_regs_0_UserCLK
timestamp 1486834041
transform 1 0 10752 0 -1 36848
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout38
timestamp 1486834041
transform 1 0 6384 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout39
timestamp 1486834041
transform 1 0 10416 0 1 19600
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout40
timestamp 1486834041
transform 1 0 6272 0 1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout41
timestamp 1486834041
transform 1 0 6944 0 -1 29008
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout42
timestamp 1486834041
transform 1 0 8736 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout43
timestamp 1486834041
transform 1 0 5936 0 1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout44
timestamp 1486834041
transform 1 0 4816 0 1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout45
timestamp 1486834041
transform 1 0 4816 0 1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout46
timestamp 1486834041
transform -1 0 4144 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout47
timestamp 1486834041
transform -1 0 2464 0 -1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout48
timestamp 1486834041
transform 1 0 6944 0 -1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout49
timestamp 1486834041
transform 1 0 3920 0 -1 29008
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout50
timestamp 1486834041
transform -1 0 1792 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout51
timestamp 1486834041
transform -1 0 14224 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout52
timestamp 1486834041
transform 1 0 12656 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout53
timestamp 1486834041
transform 1 0 8624 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout54
timestamp 1486834041
transform -1 0 8176 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout55
timestamp 1486834041
transform 1 0 11536 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2
timestamp 1486834041
transform 1 0 896 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36
timestamp 1486834041
transform 1 0 4704 0 1 784
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52
timestamp 1486834041
transform 1 0 6496 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70
timestamp 1486834041
transform 1 0 8512 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104
timestamp 1486834041
transform 1 0 12320 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 16128 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_172
timestamp 1486834041
transform 1 0 19936 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_206
timestamp 1486834041
transform 1 0 23744 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_240
timestamp 1486834041
transform 1 0 27552 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_10
timestamp 1486834041
transform 1 0 1792 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_42
timestamp 1486834041
transform 1 0 5376 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_58
timestamp 1486834041
transform 1 0 7168 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1486834041
transform 1 0 8064 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_72
timestamp 1486834041
transform 1 0 8736 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_88
timestamp 1486834041
transform 1 0 10528 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_92
timestamp 1486834041
transform 1 0 10976 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_94
timestamp 1486834041
transform 1 0 11200 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_103
timestamp 1486834041
transform 1 0 12208 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_119
timestamp 1486834041
transform 1 0 14000 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_135
timestamp 1486834041
transform 1 0 15792 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_139
timestamp 1486834041
transform 1 0 16240 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_142
timestamp 1486834041
transform 1 0 16576 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_206
timestamp 1486834041
transform 1 0 23744 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_212
timestamp 1486834041
transform 1 0 24416 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_216
timestamp 1486834041
transform 1 0 24864 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_10
timestamp 1486834041
transform 1 0 1792 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_26
timestamp 1486834041
transform 1 0 3584 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1486834041
transform 1 0 4480 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1486834041
transform 1 0 4816 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1486834041
transform 1 0 11984 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_107
timestamp 1486834041
transform 1 0 12656 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 19824 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_177
timestamp 1486834041
transform 1 0 20496 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_209
timestamp 1486834041
transform 1 0 24080 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_16
timestamp 1486834041
transform 1 0 2464 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_48
timestamp 1486834041
transform 1 0 6048 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_64
timestamp 1486834041
transform 1 0 7840 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_68
timestamp 1486834041
transform 1 0 8288 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_72
timestamp 1486834041
transform 1 0 8736 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_136
timestamp 1486834041
transform 1 0 15904 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_142
timestamp 1486834041
transform 1 0 16576 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_206
timestamp 1486834041
transform 1 0 23744 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_212
timestamp 1486834041
transform 1 0 24416 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_220
timestamp 1486834041
transform 1 0 25312 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_224
timestamp 1486834041
transform 1 0 25760 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_16
timestamp 1486834041
transform 1 0 2464 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_32
timestamp 1486834041
transform 1 0 4256 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 4480 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1486834041
transform 1 0 4816 0 1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1486834041
transform 1 0 11984 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_107
timestamp 1486834041
transform 1 0 12656 0 1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_171
timestamp 1486834041
transform 1 0 19824 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_177
timestamp 1486834041
transform 1 0 20496 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_209
timestamp 1486834041
transform 1 0 24080 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_225
timestamp 1486834041
transform 1 0 25872 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_32
timestamp 1486834041
transform 1 0 4256 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_48
timestamp 1486834041
transform 1 0 6048 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_56
timestamp 1486834041
transform 1 0 6944 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_60
timestamp 1486834041
transform 1 0 7392 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_72
timestamp 1486834041
transform 1 0 8736 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_88
timestamp 1486834041
transform 1 0 10528 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_96
timestamp 1486834041
transform 1 0 11424 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_100
timestamp 1486834041
transform 1 0 11872 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_138
timestamp 1486834041
transform 1 0 16128 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_142
timestamp 1486834041
transform 1 0 16576 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_206
timestamp 1486834041
transform 1 0 23744 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_212
timestamp 1486834041
transform 1 0 24416 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_220
timestamp 1486834041
transform 1 0 25312 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_224
timestamp 1486834041
transform 1 0 25760 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_226
timestamp 1486834041
transform 1 0 25984 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_24
timestamp 1486834041
transform 1 0 3360 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_32
timestamp 1486834041
transform 1 0 4256 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 4480 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_37
timestamp 1486834041
transform 1 0 4816 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_53
timestamp 1486834041
transform 1 0 6608 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_81
timestamp 1486834041
transform 1 0 9744 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_89
timestamp 1486834041
transform 1 0 10640 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_93
timestamp 1486834041
transform 1 0 11088 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_95
timestamp 1486834041
transform 1 0 11312 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_104
timestamp 1486834041
transform 1 0 12320 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_107
timestamp 1486834041
transform 1 0 12656 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_115
timestamp 1486834041
transform 1 0 13552 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_148
timestamp 1486834041
transform 1 0 17248 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_164
timestamp 1486834041
transform 1 0 19040 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_172
timestamp 1486834041
transform 1 0 19936 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_174
timestamp 1486834041
transform 1 0 20160 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_177
timestamp 1486834041
transform 1 0 20496 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_209
timestamp 1486834041
transform 1 0 24080 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_217
timestamp 1486834041
transform 1 0 24976 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_30
timestamp 1486834041
transform 1 0 4032 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_62
timestamp 1486834041
transform 1 0 7616 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_72
timestamp 1486834041
transform 1 0 8736 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_76
timestamp 1486834041
transform 1 0 9184 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_78
timestamp 1486834041
transform 1 0 9408 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_87
timestamp 1486834041
transform 1 0 10416 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_99
timestamp 1486834041
transform 1 0 11760 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_121
timestamp 1486834041
transform 1 0 14224 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_137
timestamp 1486834041
transform 1 0 16016 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_139
timestamp 1486834041
transform 1 0 16240 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_142
timestamp 1486834041
transform 1 0 16576 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_206
timestamp 1486834041
transform 1 0 23744 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_212
timestamp 1486834041
transform 1 0 24416 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_220
timestamp 1486834041
transform 1 0 25312 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_224
timestamp 1486834041
transform 1 0 25760 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_30
timestamp 1486834041
transform 1 0 4032 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 4480 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_45
timestamp 1486834041
transform 1 0 5712 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_61
timestamp 1486834041
transform 1 0 7504 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_69
timestamp 1486834041
transform 1 0 8400 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_73
timestamp 1486834041
transform 1 0 8848 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_94
timestamp 1486834041
transform 1 0 11200 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_98
timestamp 1486834041
transform 1 0 11648 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_100
timestamp 1486834041
transform 1 0 11872 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_127
timestamp 1486834041
transform 1 0 14896 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_131
timestamp 1486834041
transform 1 0 15344 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_151
timestamp 1486834041
transform 1 0 17584 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_167
timestamp 1486834041
transform 1 0 19376 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_177
timestamp 1486834041
transform 1 0 20496 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_209
timestamp 1486834041
transform 1 0 24080 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_30
timestamp 1486834041
transform 1 0 4032 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_34
timestamp 1486834041
transform 1 0 4480 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_36
timestamp 1486834041
transform 1 0 4704 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_72
timestamp 1486834041
transform 1 0 8736 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_80
timestamp 1486834041
transform 1 0 9632 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_84
timestamp 1486834041
transform 1 0 10080 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_154
timestamp 1486834041
transform 1 0 17920 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_162
timestamp 1486834041
transform 1 0 18816 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_166
timestamp 1486834041
transform 1 0 19264 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_199
timestamp 1486834041
transform 1 0 22960 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_207
timestamp 1486834041
transform 1 0 23856 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_209
timestamp 1486834041
transform 1 0 24080 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_212
timestamp 1486834041
transform 1 0 24416 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_220
timestamp 1486834041
transform 1 0 25312 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_224
timestamp 1486834041
transform 1 0 25760 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_226
timestamp 1486834041
transform 1 0 25984 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_30
timestamp 1486834041
transform 1 0 4032 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1486834041
transform 1 0 4480 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_53
timestamp 1486834041
transform 1 0 6608 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_83
timestamp 1486834041
transform 1 0 9968 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_121
timestamp 1486834041
transform 1 0 14224 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_123
timestamp 1486834041
transform 1 0 14448 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_164
timestamp 1486834041
transform 1 0 19040 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_172
timestamp 1486834041
transform 1 0 19936 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_174
timestamp 1486834041
transform 1 0 20160 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_177
timestamp 1486834041
transform 1 0 20496 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_209
timestamp 1486834041
transform 1 0 24080 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_217
timestamp 1486834041
transform 1 0 24976 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_30
timestamp 1486834041
transform 1 0 4032 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_34
timestamp 1486834041
transform 1 0 4480 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_55
timestamp 1486834041
transform 1 0 6832 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1486834041
transform 1 0 8064 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_72
timestamp 1486834041
transform 1 0 8736 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_124
timestamp 1486834041
transform 1 0 14560 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_150
timestamp 1486834041
transform 1 0 17472 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_152
timestamp 1486834041
transform 1 0 17696 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_185
timestamp 1486834041
transform 1 0 21392 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_201
timestamp 1486834041
transform 1 0 23184 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_209
timestamp 1486834041
transform 1 0 24080 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_212
timestamp 1486834041
transform 1 0 24416 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_216
timestamp 1486834041
transform 1 0 24864 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_2
timestamp 1486834041
transform 1 0 896 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_6
timestamp 1486834041
transform 1 0 1344 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_8
timestamp 1486834041
transform 1 0 1568 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_29
timestamp 1486834041
transform 1 0 3920 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_33
timestamp 1486834041
transform 1 0 4368 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_69
timestamp 1486834041
transform 1 0 8400 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_86
timestamp 1486834041
transform 1 0 10304 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_119
timestamp 1486834041
transform 1 0 14000 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_121
timestamp 1486834041
transform 1 0 14224 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_177
timestamp 1486834041
transform 1 0 20496 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_209
timestamp 1486834041
transform 1 0 24080 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_2
timestamp 1486834041
transform 1 0 896 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_34
timestamp 1486834041
transform 1 0 4480 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_84
timestamp 1486834041
transform 1 0 10080 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_88
timestamp 1486834041
transform 1 0 10528 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_123
timestamp 1486834041
transform 1 0 14448 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_127
timestamp 1486834041
transform 1 0 14896 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_129
timestamp 1486834041
transform 1 0 15120 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_136
timestamp 1486834041
transform 1 0 15904 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_148
timestamp 1486834041
transform 1 0 17248 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_150
timestamp 1486834041
transform 1 0 17472 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_183
timestamp 1486834041
transform 1 0 21168 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_199
timestamp 1486834041
transform 1 0 22960 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_208
timestamp 1486834041
transform 1 0 23968 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_212
timestamp 1486834041
transform 1 0 24416 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_220
timestamp 1486834041
transform 1 0 25312 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_224
timestamp 1486834041
transform 1 0 25760 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_2
timestamp 1486834041
transform 1 0 896 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_6
timestamp 1486834041
transform 1 0 1344 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_8
timestamp 1486834041
transform 1 0 1568 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_29
timestamp 1486834041
transform 1 0 3920 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_33
timestamp 1486834041
transform 1 0 4368 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_103
timestamp 1486834041
transform 1 0 12208 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_121
timestamp 1486834041
transform 1 0 14224 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_123
timestamp 1486834041
transform 1 0 14448 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_174
timestamp 1486834041
transform 1 0 20160 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_189
timestamp 1486834041
transform 1 0 21840 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_213
timestamp 1486834041
transform 1 0 24528 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_221
timestamp 1486834041
transform 1 0 25424 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_78
timestamp 1486834041
transform 1 0 9408 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_163
timestamp 1486834041
transform 1 0 18928 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_196
timestamp 1486834041
transform 1 0 22624 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_204
timestamp 1486834041
transform 1 0 23520 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_208
timestamp 1486834041
transform 1 0 23968 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_220
timestamp 1486834041
transform 1 0 25312 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_224
timestamp 1486834041
transform 1 0 25760 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_2
timestamp 1486834041
transform 1 0 896 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_6
timestamp 1486834041
transform 1 0 1344 0 1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_51
timestamp 1486834041
transform 1 0 6384 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_113
timestamp 1486834041
transform 1 0 13328 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_162
timestamp 1486834041
transform 1 0 18816 0 1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_223
timestamp 1486834041
transform 1 0 25648 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_2
timestamp 1486834041
transform 1 0 896 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_26
timestamp 1486834041
transform 1 0 3584 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_79
timestamp 1486834041
transform 1 0 9520 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_148
timestamp 1486834041
transform 1 0 17248 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_150
timestamp 1486834041
transform 1 0 17472 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_203
timestamp 1486834041
transform 1 0 23408 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_207
timestamp 1486834041
transform 1 0 23856 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_209
timestamp 1486834041
transform 1 0 24080 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_232
timestamp 1486834041
transform 1 0 26656 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_2
timestamp 1486834041
transform 1 0 896 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_6
timestamp 1486834041
transform 1 0 1344 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_107
timestamp 1486834041
transform 1 0 12656 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_115
timestamp 1486834041
transform 1 0 13552 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_117
timestamp 1486834041
transform 1 0 13776 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_156
timestamp 1486834041
transform 1 0 18144 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_167
timestamp 1486834041
transform 1 0 19376 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_209
timestamp 1486834041
transform 1 0 24080 0 1 14896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_2
timestamp 1486834041
transform 1 0 896 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_43
timestamp 1486834041
transform 1 0 5488 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_78
timestamp 1486834041
transform 1 0 9408 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_80
timestamp 1486834041
transform 1 0 9632 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_89
timestamp 1486834041
transform 1 0 10640 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_139
timestamp 1486834041
transform 1 0 16240 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_194
timestamp 1486834041
transform 1 0 22400 0 -1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_212
timestamp 1486834041
transform 1 0 24416 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_220
timestamp 1486834041
transform 1 0 25312 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_224
timestamp 1486834041
transform 1 0 25760 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_30
timestamp 1486834041
transform 1 0 4032 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1486834041
transform 1 0 4480 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_51
timestamp 1486834041
transform 1 0 6384 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_107
timestamp 1486834041
transform 1 0 12656 0 1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_123
timestamp 1486834041
transform 1 0 14448 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_174
timestamp 1486834041
transform 1 0 20160 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_183
timestamp 1486834041
transform 1 0 21168 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_187
timestamp 1486834041
transform 1 0 21616 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_189
timestamp 1486834041
transform 1 0 21840 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_210
timestamp 1486834041
transform 1 0 24192 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_218
timestamp 1486834041
transform 1 0 25088 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_222
timestamp 1486834041
transform 1 0 25536 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_224
timestamp 1486834041
transform 1 0 25760 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_2
timestamp 1486834041
transform 1 0 896 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_120
timestamp 1486834041
transform 1 0 14112 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_136
timestamp 1486834041
transform 1 0 15904 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_204
timestamp 1486834041
transform 1 0 23520 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_208
timestamp 1486834041
transform 1 0 23968 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_220
timestamp 1486834041
transform 1 0 25312 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_224
timestamp 1486834041
transform 1 0 25760 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_2
timestamp 1486834041
transform 1 0 896 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_6
timestamp 1486834041
transform 1 0 1344 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_127
timestamp 1486834041
transform 1 0 14896 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_131
timestamp 1486834041
transform 1 0 15344 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_172
timestamp 1486834041
transform 1 0 19936 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_174
timestamp 1486834041
transform 1 0 20160 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_209
timestamp 1486834041
transform 1 0 24080 0 1 18032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_16
timestamp 1486834041
transform 1 0 2464 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_72
timestamp 1486834041
transform 1 0 8736 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_142
timestamp 1486834041
transform 1 0 16576 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_186
timestamp 1486834041
transform 1 0 21504 0 -1 19600
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_202
timestamp 1486834041
transform 1 0 23296 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_212
timestamp 1486834041
transform 1 0 24416 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_220
timestamp 1486834041
transform 1 0 25312 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_232
timestamp 1486834041
transform 1 0 26656 0 -1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_2
timestamp 1486834041
transform 1 0 896 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_26
timestamp 1486834041
transform 1 0 3584 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1486834041
transform 1 0 4480 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_51
timestamp 1486834041
transform 1 0 6384 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1486834041
transform 1 0 11984 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_165
timestamp 1486834041
transform 1 0 19152 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_183
timestamp 1486834041
transform 1 0 21168 0 1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_215
timestamp 1486834041
transform 1 0 24752 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_223
timestamp 1486834041
transform 1 0 25648 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_2
timestamp 1486834041
transform 1 0 896 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_64
timestamp 1486834041
transform 1 0 7840 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_68
timestamp 1486834041
transform 1 0 8288 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_80
timestamp 1486834041
transform 1 0 9632 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_84
timestamp 1486834041
transform 1 0 10080 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_117
timestamp 1486834041
transform 1 0 13776 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_119
timestamp 1486834041
transform 1 0 14000 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_157
timestamp 1486834041
transform 1 0 18256 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_159
timestamp 1486834041
transform 1 0 18480 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_192
timestamp 1486834041
transform 1 0 22176 0 -1 21168
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_208
timestamp 1486834041
transform 1 0 23968 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_212
timestamp 1486834041
transform 1 0 24416 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_240
timestamp 1486834041
transform 1 0 27552 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_2
timestamp 1486834041
transform 1 0 896 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_10
timestamp 1486834041
transform 1 0 1792 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_14
timestamp 1486834041
transform 1 0 2240 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_37
timestamp 1486834041
transform 1 0 4816 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_39
timestamp 1486834041
transform 1 0 5040 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_72
timestamp 1486834041
transform 1 0 8736 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_80
timestamp 1486834041
transform 1 0 9632 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_84
timestamp 1486834041
transform 1 0 10080 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_107
timestamp 1486834041
transform 1 0 12656 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_111
timestamp 1486834041
transform 1 0 13104 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_121
timestamp 1486834041
transform 1 0 14224 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_154
timestamp 1486834041
transform 1 0 17920 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_200
timestamp 1486834041
transform 1 0 23072 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_210
timestamp 1486834041
transform 1 0 24192 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_218
timestamp 1486834041
transform 1 0 25088 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_36
timestamp 1486834041
transform 1 0 4704 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_40
timestamp 1486834041
transform 1 0 5152 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_61
timestamp 1486834041
transform 1 0 7504 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_69
timestamp 1486834041
transform 1 0 8400 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_72
timestamp 1486834041
transform 1 0 8736 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_116
timestamp 1486834041
transform 1 0 13664 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_162
timestamp 1486834041
transform 1 0 18816 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_164
timestamp 1486834041
transform 1 0 19040 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_205
timestamp 1486834041
transform 1 0 23632 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_209
timestamp 1486834041
transform 1 0 24080 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1486834041
transform 1 0 24416 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_2
timestamp 1486834041
transform 1 0 896 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_31
timestamp 1486834041
transform 1 0 4144 0 1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_37
timestamp 1486834041
transform 1 0 4816 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_81
timestamp 1486834041
transform 1 0 9744 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_83
timestamp 1486834041
transform 1 0 9968 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_104
timestamp 1486834041
transform 1 0 12320 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_107
timestamp 1486834041
transform 1 0 12656 0 1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_119
timestamp 1486834041
transform 1 0 14000 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_121
timestamp 1486834041
transform 1 0 14224 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_142
timestamp 1486834041
transform 1 0 16576 0 1 22736
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_158
timestamp 1486834041
transform 1 0 18368 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_166
timestamp 1486834041
transform 1 0 19264 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_177
timestamp 1486834041
transform 1 0 20496 0 1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_209
timestamp 1486834041
transform 1 0 24080 0 1 22736
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_225
timestamp 1486834041
transform 1 0 25872 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_10
timestamp 1486834041
transform 1 0 1792 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1486834041
transform 1 0 8064 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_72
timestamp 1486834041
transform 1 0 8736 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_80
timestamp 1486834041
transform 1 0 9632 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_84
timestamp 1486834041
transform 1 0 10080 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_125
timestamp 1486834041
transform 1 0 14672 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_129
timestamp 1486834041
transform 1 0 15120 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_139
timestamp 1486834041
transform 1 0 16240 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_202
timestamp 1486834041
transform 1 0 23296 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1486834041
transform 1 0 24416 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_2
timestamp 1486834041
transform 1 0 896 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_6
timestamp 1486834041
transform 1 0 1344 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_28
timestamp 1486834041
transform 1 0 3808 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_32
timestamp 1486834041
transform 1 0 4256 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1486834041
transform 1 0 4480 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_51
timestamp 1486834041
transform 1 0 6384 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_95
timestamp 1486834041
transform 1 0 11312 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_103
timestamp 1486834041
transform 1 0 12208 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_115
timestamp 1486834041
transform 1 0 13552 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_163
timestamp 1486834041
transform 1 0 18928 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_171
timestamp 1486834041
transform 1 0 19824 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_209
timestamp 1486834041
transform 1 0 24080 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_48
timestamp 1486834041
transform 1 0 6048 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_112
timestamp 1486834041
transform 1 0 13216 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_150
timestamp 1486834041
transform 1 0 17472 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_158
timestamp 1486834041
transform 1 0 18368 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_195
timestamp 1486834041
transform 1 0 22512 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_203
timestamp 1486834041
transform 1 0 23408 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_207
timestamp 1486834041
transform 1 0 23856 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_209
timestamp 1486834041
transform 1 0 24080 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1486834041
transform 1 0 24416 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_2
timestamp 1486834041
transform 1 0 896 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_6
timestamp 1486834041
transform 1 0 1344 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_8
timestamp 1486834041
transform 1 0 1568 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_29
timestamp 1486834041
transform 1 0 3920 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_33
timestamp 1486834041
transform 1 0 4368 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_45
timestamp 1486834041
transform 1 0 5712 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_47
timestamp 1486834041
transform 1 0 5936 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_68
timestamp 1486834041
transform 1 0 8288 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_72
timestamp 1486834041
transform 1 0 8736 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_107
timestamp 1486834041
transform 1 0 12656 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_137
timestamp 1486834041
transform 1 0 16016 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_145
timestamp 1486834041
transform 1 0 16912 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_197
timestamp 1486834041
transform 1 0 22736 0 1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_213
timestamp 1486834041
transform 1 0 24528 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_221
timestamp 1486834041
transform 1 0 25424 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_225
timestamp 1486834041
transform 1 0 25872 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_54
timestamp 1486834041
transform 1 0 6720 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_92
timestamp 1486834041
transform 1 0 10976 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_134
timestamp 1486834041
transform 1 0 15680 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_138
timestamp 1486834041
transform 1 0 16128 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_142
timestamp 1486834041
transform 1 0 16576 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_146
timestamp 1486834041
transform 1 0 17024 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_180
timestamp 1486834041
transform 1 0 20832 0 -1 27440
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_196
timestamp 1486834041
transform 1 0 22624 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_204
timestamp 1486834041
transform 1 0 23520 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_208
timestamp 1486834041
transform 1 0 23968 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1486834041
transform 1 0 24416 0 -1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_10
timestamp 1486834041
transform 1 0 1792 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_32
timestamp 1486834041
transform 1 0 4256 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1486834041
transform 1 0 4480 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_45
timestamp 1486834041
transform 1 0 5712 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_49
timestamp 1486834041
transform 1 0 6160 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_84
timestamp 1486834041
transform 1 0 10080 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_107
timestamp 1486834041
transform 1 0 12656 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_111
timestamp 1486834041
transform 1 0 13104 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_113
timestamp 1486834041
transform 1 0 13328 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_146
timestamp 1486834041
transform 1 0 17024 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_150
timestamp 1486834041
transform 1 0 17472 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_152
timestamp 1486834041
transform 1 0 17696 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_173
timestamp 1486834041
transform 1 0 20048 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_185
timestamp 1486834041
transform 1 0 21392 0 1 27440
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_201
timestamp 1486834041
transform 1 0 23184 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_209
timestamp 1486834041
transform 1 0 24080 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_2
timestamp 1486834041
transform 1 0 896 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_6
timestamp 1486834041
transform 1 0 1344 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_8
timestamp 1486834041
transform 1 0 1568 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_51
timestamp 1486834041
transform 1 0 6384 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_55
timestamp 1486834041
transform 1 0 6832 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_72
timestamp 1486834041
transform 1 0 8736 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_128
timestamp 1486834041
transform 1 0 15008 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_130
timestamp 1486834041
transform 1 0 15232 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_139
timestamp 1486834041
transform 1 0 16240 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_142
timestamp 1486834041
transform 1 0 16576 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_198
timestamp 1486834041
transform 1 0 22848 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_206
timestamp 1486834041
transform 1 0 23744 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_212
timestamp 1486834041
transform 1 0 24416 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_220
timestamp 1486834041
transform 1 0 25312 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_224
timestamp 1486834041
transform 1 0 25760 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_226
timestamp 1486834041
transform 1 0 25984 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_10
timestamp 1486834041
transform 1 0 1792 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_14
timestamp 1486834041
transform 1 0 2240 0 1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_37
timestamp 1486834041
transform 1 0 4816 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_61
timestamp 1486834041
transform 1 0 7504 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_65
timestamp 1486834041
transform 1 0 7952 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_87
timestamp 1486834041
transform 1 0 10416 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_95
timestamp 1486834041
transform 1 0 11312 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_107
timestamp 1486834041
transform 1 0 12656 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_111
timestamp 1486834041
transform 1 0 13104 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_173
timestamp 1486834041
transform 1 0 20048 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_177
timestamp 1486834041
transform 1 0 20496 0 1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_209
timestamp 1486834041
transform 1 0 24080 0 1 29008
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_225
timestamp 1486834041
transform 1 0 25872 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_80
timestamp 1486834041
transform 1 0 9632 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_84
timestamp 1486834041
transform 1 0 10080 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_137
timestamp 1486834041
transform 1 0 16016 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_139
timestamp 1486834041
transform 1 0 16240 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_142
timestamp 1486834041
transform 1 0 16576 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_203
timestamp 1486834041
transform 1 0 23408 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_207
timestamp 1486834041
transform 1 0 23856 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_209
timestamp 1486834041
transform 1 0 24080 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_212
timestamp 1486834041
transform 1 0 24416 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_220
timestamp 1486834041
transform 1 0 25312 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_224
timestamp 1486834041
transform 1 0 25760 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_226
timestamp 1486834041
transform 1 0 25984 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_10
timestamp 1486834041
transform 1 0 1792 0 1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_14
timestamp 1486834041
transform 1 0 2240 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_107
timestamp 1486834041
transform 1 0 12656 0 1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_163
timestamp 1486834041
transform 1 0 18928 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_171
timestamp 1486834041
transform 1 0 19824 0 1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_209
timestamp 1486834041
transform 1 0 24080 0 1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_2
timestamp 1486834041
transform 1 0 896 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_26
timestamp 1486834041
transform 1 0 3584 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_34
timestamp 1486834041
transform 1 0 4480 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_72
timestamp 1486834041
transform 1 0 8736 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_76
timestamp 1486834041
transform 1 0 9184 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_78
timestamp 1486834041
transform 1 0 9408 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_127
timestamp 1486834041
transform 1 0 14896 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_135
timestamp 1486834041
transform 1 0 15792 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_139
timestamp 1486834041
transform 1 0 16240 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_150
timestamp 1486834041
transform 1 0 17472 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_152
timestamp 1486834041
transform 1 0 17696 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_205
timestamp 1486834041
transform 1 0 23632 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_209
timestamp 1486834041
transform 1 0 24080 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1486834041
transform 1 0 24416 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_30
timestamp 1486834041
transform 1 0 4032 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1486834041
transform 1 0 4480 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_51
timestamp 1486834041
transform 1 0 6384 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_55
timestamp 1486834041
transform 1 0 6832 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_76
timestamp 1486834041
transform 1 0 9184 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_78
timestamp 1486834041
transform 1 0 9408 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_99
timestamp 1486834041
transform 1 0 11760 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_103
timestamp 1486834041
transform 1 0 12208 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_107
timestamp 1486834041
transform 1 0 12656 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_111
timestamp 1486834041
transform 1 0 13104 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_113
timestamp 1486834041
transform 1 0 13328 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_172
timestamp 1486834041
transform 1 0 19936 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_174
timestamp 1486834041
transform 1 0 20160 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_193
timestamp 1486834041
transform 1 0 22288 0 1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_225
timestamp 1486834041
transform 1 0 25872 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_10
timestamp 1486834041
transform 1 0 1792 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_12
timestamp 1486834041
transform 1 0 2016 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_45
timestamp 1486834041
transform 1 0 5712 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_49
timestamp 1486834041
transform 1 0 6160 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_80
timestamp 1486834041
transform 1 0 9632 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_142
timestamp 1486834041
transform 1 0 16576 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_150
timestamp 1486834041
transform 1 0 17472 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_154
timestamp 1486834041
transform 1 0 17920 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_175
timestamp 1486834041
transform 1 0 20272 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_207
timestamp 1486834041
transform 1 0 23856 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_209
timestamp 1486834041
transform 1 0 24080 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1486834041
transform 1 0 24416 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_2
timestamp 1486834041
transform 1 0 896 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_103
timestamp 1486834041
transform 1 0 12208 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_143
timestamp 1486834041
transform 1 0 16688 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_145
timestamp 1486834041
transform 1 0 16912 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_166
timestamp 1486834041
transform 1 0 19264 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_177
timestamp 1486834041
transform 1 0 20496 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_209
timestamp 1486834041
transform 1 0 24080 0 1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_72
timestamp 1486834041
transform 1 0 8736 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_76
timestamp 1486834041
transform 1 0 9184 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_86
timestamp 1486834041
transform 1 0 10304 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_142
timestamp 1486834041
transform 1 0 16576 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_146
timestamp 1486834041
transform 1 0 17024 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_188
timestamp 1486834041
transform 1 0 21728 0 -1 35280
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_204
timestamp 1486834041
transform 1 0 23520 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_208
timestamp 1486834041
transform 1 0 23968 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1486834041
transform 1 0 24416 0 -1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_22
timestamp 1486834041
transform 1 0 3136 0 1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_26
timestamp 1486834041
transform 1 0 3584 0 1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_37
timestamp 1486834041
transform 1 0 4816 0 1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_157
timestamp 1486834041
transform 1 0 18256 0 1 35280
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_173
timestamp 1486834041
transform 1 0 20048 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_177
timestamp 1486834041
transform 1 0 20496 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_209
timestamp 1486834041
transform 1 0 24080 0 1 35280
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_225
timestamp 1486834041
transform 1 0 25872 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_2
timestamp 1486834041
transform 1 0 896 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_10
timestamp 1486834041
transform 1 0 1792 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_67
timestamp 1486834041
transform 1 0 8176 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_69
timestamp 1486834041
transform 1 0 8400 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_72
timestamp 1486834041
transform 1 0 8736 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_80
timestamp 1486834041
transform 1 0 9632 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_178
timestamp 1486834041
transform 1 0 20608 0 -1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1486834041
transform 1 0 24416 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_2
timestamp 1486834041
transform 1 0 896 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_6
timestamp 1486834041
transform 1 0 1344 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_37
timestamp 1486834041
transform 1 0 4816 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_45
timestamp 1486834041
transform 1 0 5712 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_107
timestamp 1486834041
transform 1 0 12656 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_160
timestamp 1486834041
transform 1 0 18592 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_168
timestamp 1486834041
transform 1 0 19488 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_172
timestamp 1486834041
transform 1 0 19936 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_174
timestamp 1486834041
transform 1 0 20160 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_177
timestamp 1486834041
transform 1 0 20496 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_209
timestamp 1486834041
transform 1 0 24080 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_2
timestamp 1486834041
transform 1 0 896 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_23
timestamp 1486834041
transform 1 0 3248 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_27
timestamp 1486834041
transform 1 0 3696 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_29
timestamp 1486834041
transform 1 0 3920 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_72
timestamp 1486834041
transform 1 0 8736 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_76
timestamp 1486834041
transform 1 0 9184 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_127
timestamp 1486834041
transform 1 0 14896 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_136
timestamp 1486834041
transform 1 0 15904 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_142
timestamp 1486834041
transform 1 0 16576 0 -1 38416
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_206
timestamp 1486834041
transform 1 0 23744 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1486834041
transform 1 0 24416 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_10
timestamp 1486834041
transform 1 0 1792 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_31
timestamp 1486834041
transform 1 0 4144 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_37
timestamp 1486834041
transform 1 0 4816 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_59
timestamp 1486834041
transform 1 0 7280 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_63
timestamp 1486834041
transform 1 0 7728 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_96
timestamp 1486834041
transform 1 0 11424 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_147
timestamp 1486834041
transform 1 0 17136 0 1 38416
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_163
timestamp 1486834041
transform 1 0 18928 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_171
timestamp 1486834041
transform 1 0 19824 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_177
timestamp 1486834041
transform 1 0 20496 0 1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_209
timestamp 1486834041
transform 1 0 24080 0 1 38416
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_225
timestamp 1486834041
transform 1 0 25872 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_2
timestamp 1486834041
transform 1 0 896 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_6
timestamp 1486834041
transform 1 0 1344 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_31
timestamp 1486834041
transform 1 0 4144 0 -1 39984
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_47
timestamp 1486834041
transform 1 0 5936 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_49
timestamp 1486834041
transform 1 0 6160 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_66
timestamp 1486834041
transform 1 0 8064 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_72
timestamp 1486834041
transform 1 0 8736 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_131
timestamp 1486834041
transform 1 0 15344 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_139
timestamp 1486834041
transform 1 0 16240 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_142
timestamp 1486834041
transform 1 0 16576 0 -1 39984
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_206
timestamp 1486834041
transform 1 0 23744 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1486834041
transform 1 0 24416 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_26
timestamp 1486834041
transform 1 0 3584 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1486834041
transform 1 0 4480 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_37
timestamp 1486834041
transform 1 0 4816 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_45
timestamp 1486834041
transform 1 0 5712 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_79
timestamp 1486834041
transform 1 0 9520 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_83
timestamp 1486834041
transform 1 0 9968 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_115
timestamp 1486834041
transform 1 0 13552 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_119
timestamp 1486834041
transform 1 0 14000 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_140
timestamp 1486834041
transform 1 0 16352 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_172
timestamp 1486834041
transform 1 0 19936 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_174
timestamp 1486834041
transform 1 0 20160 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_177
timestamp 1486834041
transform 1 0 20496 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_209
timestamp 1486834041
transform 1 0 24080 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_18
timestamp 1486834041
transform 1 0 2688 0 -1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_50
timestamp 1486834041
transform 1 0 6272 0 -1 41552
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_66
timestamp 1486834041
transform 1 0 8064 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_92
timestamp 1486834041
transform 1 0 10976 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_96
timestamp 1486834041
transform 1 0 11424 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_105
timestamp 1486834041
transform 1 0 12432 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_113
timestamp 1486834041
transform 1 0 13328 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_135
timestamp 1486834041
transform 1 0 15792 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_139
timestamp 1486834041
transform 1 0 16240 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_142
timestamp 1486834041
transform 1 0 16576 0 -1 41552
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_206
timestamp 1486834041
transform 1 0 23744 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1486834041
transform 1 0 24416 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_18
timestamp 1486834041
transform 1 0 2688 0 1 41552
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1486834041
transform 1 0 4480 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1486834041
transform 1 0 4816 0 1 41552
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1486834041
transform 1 0 11984 0 1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_107
timestamp 1486834041
transform 1 0 12656 0 1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_115
timestamp 1486834041
transform 1 0 13552 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_117
timestamp 1486834041
transform 1 0 13776 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_138
timestamp 1486834041
transform 1 0 16128 0 1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_170
timestamp 1486834041
transform 1 0 19712 0 1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_174
timestamp 1486834041
transform 1 0 20160 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_177
timestamp 1486834041
transform 1 0 20496 0 1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_209
timestamp 1486834041
transform 1 0 24080 0 1 41552
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_225
timestamp 1486834041
transform 1 0 25872 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_18
timestamp 1486834041
transform 1 0 2688 0 -1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_50
timestamp 1486834041
transform 1 0 6272 0 -1 43120
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_66
timestamp 1486834041
transform 1 0 8064 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_72
timestamp 1486834041
transform 1 0 8736 0 -1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_136
timestamp 1486834041
transform 1 0 15904 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_142
timestamp 1486834041
transform 1 0 16576 0 -1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_206
timestamp 1486834041
transform 1 0 23744 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1486834041
transform 1 0 24416 0 -1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_10
timestamp 1486834041
transform 1 0 1792 0 1 43120
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_26
timestamp 1486834041
transform 1 0 3584 0 1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1486834041
transform 1 0 4480 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_37
timestamp 1486834041
transform 1 0 4816 0 1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_101
timestamp 1486834041
transform 1 0 11984 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_107
timestamp 1486834041
transform 1 0 12656 0 1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_171
timestamp 1486834041
transform 1 0 19824 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_177
timestamp 1486834041
transform 1 0 20496 0 1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_209
timestamp 1486834041
transform 1 0 24080 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_10
timestamp 1486834041
transform 1 0 1792 0 -1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_42
timestamp 1486834041
transform 1 0 5376 0 -1 44688
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_58
timestamp 1486834041
transform 1 0 7168 0 -1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_66
timestamp 1486834041
transform 1 0 8064 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_72
timestamp 1486834041
transform 1 0 8736 0 -1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_136
timestamp 1486834041
transform 1 0 15904 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_142
timestamp 1486834041
transform 1 0 16576 0 -1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_206
timestamp 1486834041
transform 1 0 23744 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1486834041
transform 1 0 24416 0 -1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_10
timestamp 1486834041
transform 1 0 1792 0 1 44688
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_26
timestamp 1486834041
transform 1 0 3584 0 1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1486834041
transform 1 0 4480 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_37
timestamp 1486834041
transform 1 0 4816 0 1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_101
timestamp 1486834041
transform 1 0 11984 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_107
timestamp 1486834041
transform 1 0 12656 0 1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_171
timestamp 1486834041
transform 1 0 19824 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_177
timestamp 1486834041
transform 1 0 20496 0 1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_209
timestamp 1486834041
transform 1 0 24080 0 1 44688
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_225
timestamp 1486834041
transform 1 0 25872 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_10
timestamp 1486834041
transform 1 0 1792 0 -1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_42
timestamp 1486834041
transform 1 0 5376 0 -1 46256
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_58
timestamp 1486834041
transform 1 0 7168 0 -1 46256
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_66
timestamp 1486834041
transform 1 0 8064 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_72
timestamp 1486834041
transform 1 0 8736 0 -1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_136
timestamp 1486834041
transform 1 0 15904 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_142
timestamp 1486834041
transform 1 0 16576 0 -1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_206
timestamp 1486834041
transform 1 0 23744 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1486834041
transform 1 0 24416 0 -1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_18
timestamp 1486834041
transform 1 0 2688 0 1 46256
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1486834041
transform 1 0 4480 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_37
timestamp 1486834041
transform 1 0 4816 0 1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_101
timestamp 1486834041
transform 1 0 11984 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_107
timestamp 1486834041
transform 1 0 12656 0 1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_171
timestamp 1486834041
transform 1 0 19824 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_177
timestamp 1486834041
transform 1 0 20496 0 1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_209
timestamp 1486834041
transform 1 0 24080 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_16
timestamp 1486834041
transform 1 0 2464 0 -1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_48
timestamp 1486834041
transform 1 0 6048 0 -1 47824
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_64
timestamp 1486834041
transform 1 0 7840 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_68
timestamp 1486834041
transform 1 0 8288 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_72
timestamp 1486834041
transform 1 0 8736 0 -1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_136
timestamp 1486834041
transform 1 0 15904 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_142
timestamp 1486834041
transform 1 0 16576 0 -1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_206
timestamp 1486834041
transform 1 0 23744 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1486834041
transform 1 0 24416 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_10
timestamp 1486834041
transform 1 0 1792 0 1 47824
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_26
timestamp 1486834041
transform 1 0 3584 0 1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1486834041
transform 1 0 4480 0 1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_37
timestamp 1486834041
transform 1 0 4816 0 1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_101
timestamp 1486834041
transform 1 0 11984 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_107
timestamp 1486834041
transform 1 0 12656 0 1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_171
timestamp 1486834041
transform 1 0 19824 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_177
timestamp 1486834041
transform 1 0 20496 0 1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_209
timestamp 1486834041
transform 1 0 24080 0 1 47824
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_225
timestamp 1486834041
transform 1 0 25872 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_10
timestamp 1486834041
transform 1 0 1792 0 -1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_42
timestamp 1486834041
transform 1 0 5376 0 -1 49392
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_58
timestamp 1486834041
transform 1 0 7168 0 -1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_66
timestamp 1486834041
transform 1 0 8064 0 -1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_72
timestamp 1486834041
transform 1 0 8736 0 -1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_136
timestamp 1486834041
transform 1 0 15904 0 -1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_142
timestamp 1486834041
transform 1 0 16576 0 -1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_206
timestamp 1486834041
transform 1 0 23744 0 -1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1486834041
transform 1 0 24416 0 -1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_2
timestamp 1486834041
transform 1 0 896 0 1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1486834041
transform 1 0 4480 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_37
timestamp 1486834041
transform 1 0 4816 0 1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_101
timestamp 1486834041
transform 1 0 11984 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_107
timestamp 1486834041
transform 1 0 12656 0 1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_171
timestamp 1486834041
transform 1 0 19824 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_177
timestamp 1486834041
transform 1 0 20496 0 1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_209
timestamp 1486834041
transform 1 0 24080 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_10
timestamp 1486834041
transform 1 0 1792 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_42
timestamp 1486834041
transform 1 0 5376 0 -1 50960
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_58
timestamp 1486834041
transform 1 0 7168 0 -1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_66
timestamp 1486834041
transform 1 0 8064 0 -1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_72
timestamp 1486834041
transform 1 0 8736 0 -1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_136
timestamp 1486834041
transform 1 0 15904 0 -1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_142
timestamp 1486834041
transform 1 0 16576 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_174
timestamp 1486834041
transform 1 0 20160 0 -1 50960
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_190
timestamp 1486834041
transform 1 0 21952 0 -1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_198
timestamp 1486834041
transform 1 0 22848 0 -1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1486834041
transform 1 0 24416 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_10
timestamp 1486834041
transform 1 0 1792 0 1 50960
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_26
timestamp 1486834041
transform 1 0 3584 0 1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1486834041
transform 1 0 4480 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1486834041
transform 1 0 4816 0 1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_101
timestamp 1486834041
transform 1 0 11984 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_107
timestamp 1486834041
transform 1 0 12656 0 1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_171
timestamp 1486834041
transform 1 0 19824 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_177
timestamp 1486834041
transform 1 0 20496 0 1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_209
timestamp 1486834041
transform 1 0 24080 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_10
timestamp 1486834041
transform 1 0 1792 0 -1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_42
timestamp 1486834041
transform 1 0 5376 0 -1 52528
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_58
timestamp 1486834041
transform 1 0 7168 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_66
timestamp 1486834041
transform 1 0 8064 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_72
timestamp 1486834041
transform 1 0 8736 0 -1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_136
timestamp 1486834041
transform 1 0 15904 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_142
timestamp 1486834041
transform 1 0 16576 0 -1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_174
timestamp 1486834041
transform 1 0 20160 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_182
timestamp 1486834041
transform 1 0 21056 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_192
timestamp 1486834041
transform 1 0 22176 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1486834041
transform 1 0 24416 0 -1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_10
timestamp 1486834041
transform 1 0 1792 0 1 52528
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_26
timestamp 1486834041
transform 1 0 3584 0 1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_34
timestamp 1486834041
transform 1 0 4480 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_37
timestamp 1486834041
transform 1 0 4816 0 1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_101
timestamp 1486834041
transform 1 0 11984 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_107
timestamp 1486834041
transform 1 0 12656 0 1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_171
timestamp 1486834041
transform 1 0 19824 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_177
timestamp 1486834041
transform 1 0 20496 0 1 52528
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_193
timestamp 1486834041
transform 1 0 22288 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_197
timestamp 1486834041
transform 1 0 22736 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_10
timestamp 1486834041
transform 1 0 1792 0 -1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_42
timestamp 1486834041
transform 1 0 5376 0 -1 54096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_58
timestamp 1486834041
transform 1 0 7168 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_66
timestamp 1486834041
transform 1 0 8064 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_72
timestamp 1486834041
transform 1 0 8736 0 -1 54096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_136
timestamp 1486834041
transform 1 0 15904 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_142
timestamp 1486834041
transform 1 0 16576 0 -1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_174
timestamp 1486834041
transform 1 0 20160 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_182
timestamp 1486834041
transform 1 0 21056 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_186
timestamp 1486834041
transform 1 0 21504 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1486834041
transform 1 0 24416 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_10
timestamp 1486834041
transform 1 0 1792 0 1 54096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_26
timestamp 1486834041
transform 1 0 3584 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_34
timestamp 1486834041
transform 1 0 4480 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_37
timestamp 1486834041
transform 1 0 4816 0 1 54096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_101
timestamp 1486834041
transform 1 0 11984 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_107
timestamp 1486834041
transform 1 0 12656 0 1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_139
timestamp 1486834041
transform 1 0 16240 0 1 54096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_155
timestamp 1486834041
transform 1 0 18032 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_171
timestamp 1486834041
transform 1 0 19824 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_10
timestamp 1486834041
transform 1 0 1792 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_12
timestamp 1486834041
transform 1 0 2016 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_27
timestamp 1486834041
transform 1 0 3696 0 -1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_43
timestamp 1486834041
transform 1 0 5488 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_47
timestamp 1486834041
transform 1 0 5936 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_63
timestamp 1486834041
transform 1 0 7728 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_67
timestamp 1486834041
transform 1 0 8176 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_69
timestamp 1486834041
transform 1 0 8400 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_72
timestamp 1486834041
transform 1 0 8736 0 -1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_88
timestamp 1486834041
transform 1 0 10528 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_96
timestamp 1486834041
transform 1 0 11424 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_111
timestamp 1486834041
transform 1 0 13104 0 -1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_127
timestamp 1486834041
transform 1 0 14896 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_135
timestamp 1486834041
transform 1 0 15792 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_139
timestamp 1486834041
transform 1 0 16240 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_142
timestamp 1486834041
transform 1 0 16576 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_144
timestamp 1486834041
transform 1 0 16800 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_159
timestamp 1486834041
transform 1 0 18480 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_167
timestamp 1486834041
transform 1 0 19376 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_207
timestamp 1486834041
transform 1 0 23856 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_209
timestamp 1486834041
transform 1 0 24080 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_212
timestamp 1486834041
transform 1 0 24416 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_8
timestamp 1486834041
transform 1 0 1568 0 1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_16
timestamp 1486834041
transform 1 0 2464 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_36
timestamp 1486834041
transform 1 0 4704 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_51
timestamp 1486834041
transform 1 0 6384 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_53
timestamp 1486834041
transform 1 0 6608 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_70
timestamp 1486834041
transform 1 0 8512 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_99
timestamp 1486834041
transform 1 0 11760 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_101
timestamp 1486834041
transform 1 0 11984 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_104
timestamp 1486834041
transform 1 0 12320 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_106
timestamp 1486834041
transform 1 0 12544 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_135
timestamp 1486834041
transform 1 0 15792 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_152
timestamp 1486834041
transform 1 0 17696 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_200
timestamp 1486834041
transform 1 0 23072 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_234
timestamp 1486834041
transform 1 0 26880 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_240
timestamp 1486834041
transform 1 0 27552 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input1
timestamp 1486834041
transform 1 0 896 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input2
timestamp 1486834041
transform 1 0 896 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input3
timestamp 1486834041
transform 1 0 2464 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input4
timestamp 1486834041
transform 1 0 4816 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input5
timestamp 1486834041
transform 1 0 896 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input6
timestamp 1486834041
transform 1 0 896 0 1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input7
timestamp 1486834041
transform 1 0 896 0 -1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input8
timestamp 1486834041
transform 1 0 2688 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input9
timestamp 1486834041
transform 1 0 896 0 1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input10
timestamp 1486834041
transform 1 0 1792 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input11
timestamp 1486834041
transform 1 0 1792 0 -1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input12
timestamp 1486834041
transform 1 0 1792 0 1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input13
timestamp 1486834041
transform 1 0 896 0 -1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input14
timestamp 1486834041
transform 1 0 896 0 1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input15
timestamp 1486834041
transform 1 0 896 0 -1 46256
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input16
timestamp 1486834041
transform 1 0 5488 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input17
timestamp 1486834041
transform 1 0 896 0 1 46256
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input18
timestamp 1486834041
transform 1 0 1792 0 1 46256
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input19
timestamp 1486834041
transform 1 0 896 0 -1 47824
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input20
timestamp 1486834041
transform 1 0 896 0 1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input21
timestamp 1486834041
transform 1 0 896 0 -1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input22
timestamp 1486834041
transform 1 0 896 0 -1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input23
timestamp 1486834041
transform 1 0 896 0 1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input24
timestamp 1486834041
transform 1 0 896 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input25
timestamp 1486834041
transform 1 0 896 0 1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input26
timestamp 1486834041
transform 1 0 896 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input27
timestamp 1486834041
transform 1 0 896 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input28
timestamp 1486834041
transform 1 0 896 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input29
timestamp 1486834041
transform 1 0 896 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input30
timestamp 1486834041
transform 1 0 896 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input31
timestamp 1486834041
transform 1 0 896 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input32
timestamp 1486834041
transform 1 0 896 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input33
timestamp 1486834041
transform 1 0 1792 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input34
timestamp 1486834041
transform 1 0 896 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input35
timestamp 1486834041
transform 1 0 896 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input36
timestamp 1486834041
transform 1 0 896 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input37
timestamp 1486834041
transform 1 0 7392 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input38
timestamp 1486834041
transform -1 0 26432 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input39
timestamp 1486834041
transform -1 0 25536 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input40
timestamp 1486834041
transform -1 0 25872 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input41
timestamp 1486834041
transform -1 0 27328 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input42
timestamp 1486834041
transform -1 0 26096 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input43
timestamp 1486834041
transform -1 0 26768 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input44
timestamp 1486834041
transform -1 0 26768 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input45
timestamp 1486834041
transform -1 0 27664 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input46
timestamp 1486834041
transform -1 0 27664 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input47
timestamp 1486834041
transform -1 0 27664 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input48
timestamp 1486834041
transform -1 0 27664 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input49
timestamp 1486834041
transform -1 0 26096 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input50
timestamp 1486834041
transform -1 0 25872 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input51
timestamp 1486834041
transform -1 0 26768 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input52
timestamp 1486834041
transform -1 0 26768 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input53
timestamp 1486834041
transform -1 0 27664 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input54
timestamp 1486834041
transform -1 0 27664 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input55
timestamp 1486834041
transform -1 0 27664 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input56
timestamp 1486834041
transform -1 0 27664 0 -1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input57
timestamp 1486834041
transform -1 0 27664 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input58
timestamp 1486834041
transform -1 0 27664 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input59
timestamp 1486834041
transform -1 0 27664 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input60
timestamp 1486834041
transform -1 0 27664 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input61
timestamp 1486834041
transform -1 0 26768 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input62
timestamp 1486834041
transform -1 0 27664 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input63
timestamp 1486834041
transform -1 0 26768 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input64
timestamp 1486834041
transform -1 0 27664 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input65
timestamp 1486834041
transform -1 0 26768 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input66
timestamp 1486834041
transform -1 0 27664 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input67
timestamp 1486834041
transform -1 0 27664 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input68
timestamp 1486834041
transform -1 0 25760 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input69
timestamp 1486834041
transform -1 0 26768 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input70
timestamp 1486834041
transform -1 0 25872 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input71
timestamp 1486834041
transform -1 0 26768 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input72
timestamp 1486834041
transform -1 0 27664 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input73
timestamp 1486834041
transform -1 0 27664 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input74
timestamp 1486834041
transform -1 0 26768 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input75
timestamp 1486834041
transform -1 0 27664 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input76
timestamp 1486834041
transform -1 0 26768 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input77
timestamp 1486834041
transform -1 0 26768 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input78
timestamp 1486834041
transform -1 0 26768 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input79
timestamp 1486834041
transform -1 0 27664 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input80
timestamp 1486834041
transform -1 0 26768 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input81
timestamp 1486834041
transform -1 0 27664 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input82
timestamp 1486834041
transform -1 0 26768 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input83
timestamp 1486834041
transform -1 0 27664 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input84
timestamp 1486834041
transform -1 0 26768 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input85
timestamp 1486834041
transform -1 0 27664 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform -1 0 2464 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform -1 0 2464 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform -1 0 4032 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform -1 0 2464 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform -1 0 7616 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform -1 0 4032 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform -1 0 4032 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform -1 0 2464 0 -1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform -1 0 6384 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform -1 0 2464 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform -1 0 2464 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform -1 0 2464 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform -1 0 2464 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform -1 0 4032 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform 1 0 4816 0 1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform 1 0 4816 0 1 16464
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform -1 0 2464 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform 1 0 4816 0 1 19600
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform -1 0 4032 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output105
timestamp 1486834041
transform -1 0 2464 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output106
timestamp 1486834041
transform -1 0 2464 0 -1 19600
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output107
timestamp 1486834041
transform -1 0 4704 0 -1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output108
timestamp 1486834041
transform 1 0 4816 0 1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output109
timestamp 1486834041
transform -1 0 2464 0 -1 25872
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output110
timestamp 1486834041
transform 1 0 24528 0 -1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output111
timestamp 1486834041
transform 1 0 26096 0 1 21168
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output112
timestamp 1486834041
transform 1 0 26096 0 -1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output113
timestamp 1486834041
transform 1 0 24528 0 -1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output114
timestamp 1486834041
transform 1 0 26096 0 1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output115
timestamp 1486834041
transform 1 0 24528 0 1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output116
timestamp 1486834041
transform 1 0 26096 0 -1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output117
timestamp 1486834041
transform 1 0 24528 0 -1 25872
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output118
timestamp 1486834041
transform 1 0 26096 0 1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output119
timestamp 1486834041
transform 1 0 26096 0 -1 25872
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output120
timestamp 1486834041
transform 1 0 24528 0 -1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output121
timestamp 1486834041
transform 1 0 26096 0 1 25872
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output122
timestamp 1486834041
transform 1 0 24528 0 1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output123
timestamp 1486834041
transform 1 0 26096 0 -1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output124
timestamp 1486834041
transform 1 0 26096 0 1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output125
timestamp 1486834041
transform 1 0 26096 0 -1 29008
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output126
timestamp 1486834041
transform 1 0 26096 0 1 29008
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output127
timestamp 1486834041
transform 1 0 26096 0 -1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output128
timestamp 1486834041
transform 1 0 26096 0 1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output129
timestamp 1486834041
transform 1 0 26096 0 -1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output130
timestamp 1486834041
transform 1 0 24528 0 -1 38416
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output131
timestamp 1486834041
transform 1 0 24528 0 -1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output132
timestamp 1486834041
transform 1 0 26096 0 -1 44688
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output133
timestamp 1486834041
transform 1 0 26096 0 -1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output134
timestamp 1486834041
transform 1 0 26096 0 1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output135
timestamp 1486834041
transform 1 0 24528 0 -1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output136
timestamp 1486834041
transform 1 0 26096 0 -1 41552
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output137
timestamp 1486834041
transform 1 0 24528 0 1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output138
timestamp 1486834041
transform 1 0 26096 0 1 41552
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output139
timestamp 1486834041
transform 1 0 24528 0 -1 41552
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output140
timestamp 1486834041
transform 1 0 26096 0 -1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output141
timestamp 1486834041
transform 1 0 26096 0 1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output142
timestamp 1486834041
transform 1 0 24528 0 1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output143
timestamp 1486834041
transform 1 0 26096 0 -1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output144
timestamp 1486834041
transform 1 0 26096 0 1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output145
timestamp 1486834041
transform 1 0 24528 0 -1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output146
timestamp 1486834041
transform 1 0 26096 0 -1 38416
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output147
timestamp 1486834041
transform 1 0 24528 0 1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output148
timestamp 1486834041
transform 1 0 26096 0 1 38416
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output149
timestamp 1486834041
transform 1 0 26096 0 1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output150
timestamp 1486834041
transform 1 0 24528 0 -1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output151
timestamp 1486834041
transform 1 0 26096 0 -1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output152
timestamp 1486834041
transform 1 0 26096 0 1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output153
timestamp 1486834041
transform 1 0 24528 0 -1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output154
timestamp 1486834041
transform 1 0 26096 0 -1 35280
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output155
timestamp 1486834041
transform 1 0 24528 0 1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output156
timestamp 1486834041
transform 1 0 26096 0 1 35280
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output157
timestamp 1486834041
transform 1 0 24528 0 -1 35280
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output158
timestamp 1486834041
transform 1 0 24528 0 1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output159
timestamp 1486834041
transform 1 0 26096 0 -1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output160
timestamp 1486834041
transform 1 0 26096 0 1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output161
timestamp 1486834041
transform 1 0 24528 0 -1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output162
timestamp 1486834041
transform 1 0 26096 0 -1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output163
timestamp 1486834041
transform 1 0 24528 0 1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output164
timestamp 1486834041
transform 1 0 26096 0 1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output165
timestamp 1486834041
transform 1 0 24528 0 -1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output166
timestamp 1486834041
transform 1 0 26096 0 -1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output167
timestamp 1486834041
transform 1 0 26096 0 1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output168
timestamp 1486834041
transform 1 0 24528 0 -1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output169
timestamp 1486834041
transform 1 0 26096 0 1 44688
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output170
timestamp 1486834041
transform 1 0 26096 0 -1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output171
timestamp 1486834041
transform 1 0 24528 0 1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output172
timestamp 1486834041
transform 1 0 26096 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output173
timestamp 1486834041
transform 1 0 24528 0 -1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output174
timestamp 1486834041
transform 1 0 26096 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output175
timestamp 1486834041
transform 1 0 24528 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output176
timestamp 1486834041
transform -1 0 24528 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output177
timestamp 1486834041
transform 1 0 22624 0 -1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output178
timestamp 1486834041
transform 1 0 20720 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output179
timestamp 1486834041
transform 1 0 21392 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output180
timestamp 1486834041
transform 1 0 24528 0 -1 44688
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output181
timestamp 1486834041
transform 1 0 24528 0 1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output182
timestamp 1486834041
transform 1 0 22960 0 1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output183
timestamp 1486834041
transform 1 0 26096 0 -1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output184
timestamp 1486834041
transform 1 0 26096 0 1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output185
timestamp 1486834041
transform 1 0 24528 0 -1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output186
timestamp 1486834041
transform 1 0 26096 0 -1 47824
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output187
timestamp 1486834041
transform 1 0 24528 0 1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output188
timestamp 1486834041
transform 1 0 26096 0 1 47824
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output189
timestamp 1486834041
transform 1 0 24528 0 -1 47824
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output190
timestamp 1486834041
transform -1 0 3696 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output191
timestamp 1486834041
transform -1 0 17696 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output192
timestamp 1486834041
transform -1 0 18480 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output193
timestamp 1486834041
transform -1 0 19712 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output194
timestamp 1486834041
transform -1 0 21504 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output195
timestamp 1486834041
transform 1 0 21504 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output196
timestamp 1486834041
transform 1 0 22288 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output197
timestamp 1486834041
transform 1 0 23744 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output198
timestamp 1486834041
transform 1 0 25312 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output199
timestamp 1486834041
transform 1 0 24528 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output200
timestamp 1486834041
transform 1 0 22624 0 -1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output201
timestamp 1486834041
transform 1 0 2912 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output202
timestamp 1486834041
transform -1 0 6384 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output203
timestamp 1486834041
transform 1 0 6160 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output204
timestamp 1486834041
transform -1 0 8288 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output205
timestamp 1486834041
transform -1 0 10192 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output206
timestamp 1486834041
transform -1 0 11760 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output207
timestamp 1486834041
transform -1 0 13104 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output208
timestamp 1486834041
transform -1 0 14224 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output209
timestamp 1486834041
transform -1 0 15792 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output210
timestamp 1486834041
transform -1 0 1568 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_71
timestamp 1486834041
transform 1 0 672 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 27888 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_72
timestamp 1486834041
transform 1 0 672 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 27888 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_73
timestamp 1486834041
transform 1 0 672 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 27888 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_74
timestamp 1486834041
transform 1 0 672 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 27888 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_75
timestamp 1486834041
transform 1 0 672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 27888 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_76
timestamp 1486834041
transform 1 0 672 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 27888 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_77
timestamp 1486834041
transform 1 0 672 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 27888 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_78
timestamp 1486834041
transform 1 0 672 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 27888 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_79
timestamp 1486834041
transform 1 0 672 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 27888 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_80
timestamp 1486834041
transform 1 0 672 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 27888 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_81
timestamp 1486834041
transform 1 0 672 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 27888 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_82
timestamp 1486834041
transform 1 0 672 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 27888 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_83
timestamp 1486834041
transform 1 0 672 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 27888 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_84
timestamp 1486834041
transform 1 0 672 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 27888 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_85
timestamp 1486834041
transform 1 0 672 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 27888 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_86
timestamp 1486834041
transform 1 0 672 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 27888 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_87
timestamp 1486834041
transform 1 0 672 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1486834041
transform -1 0 27888 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_88
timestamp 1486834041
transform 1 0 672 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1486834041
transform -1 0 27888 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_89
timestamp 1486834041
transform 1 0 672 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1486834041
transform -1 0 27888 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_90
timestamp 1486834041
transform 1 0 672 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1486834041
transform -1 0 27888 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_91
timestamp 1486834041
transform 1 0 672 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1486834041
transform -1 0 27888 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_92
timestamp 1486834041
transform 1 0 672 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1486834041
transform -1 0 27888 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_93
timestamp 1486834041
transform 1 0 672 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1486834041
transform -1 0 27888 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_94
timestamp 1486834041
transform 1 0 672 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1486834041
transform -1 0 27888 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_95
timestamp 1486834041
transform 1 0 672 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1486834041
transform -1 0 27888 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_96
timestamp 1486834041
transform 1 0 672 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1486834041
transform -1 0 27888 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_97
timestamp 1486834041
transform 1 0 672 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1486834041
transform -1 0 27888 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_98
timestamp 1486834041
transform 1 0 672 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1486834041
transform -1 0 27888 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_99
timestamp 1486834041
transform 1 0 672 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1486834041
transform -1 0 27888 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_100
timestamp 1486834041
transform 1 0 672 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1486834041
transform -1 0 27888 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_101
timestamp 1486834041
transform 1 0 672 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1486834041
transform -1 0 27888 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_102
timestamp 1486834041
transform 1 0 672 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1486834041
transform -1 0 27888 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_103
timestamp 1486834041
transform 1 0 672 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1486834041
transform -1 0 27888 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_104
timestamp 1486834041
transform 1 0 672 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1486834041
transform -1 0 27888 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_105
timestamp 1486834041
transform 1 0 672 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1486834041
transform -1 0 27888 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_106
timestamp 1486834041
transform 1 0 672 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1486834041
transform -1 0 27888 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_107
timestamp 1486834041
transform 1 0 672 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1486834041
transform -1 0 27888 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_108
timestamp 1486834041
transform 1 0 672 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1486834041
transform -1 0 27888 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_109
timestamp 1486834041
transform 1 0 672 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1486834041
transform -1 0 27888 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_110
timestamp 1486834041
transform 1 0 672 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1486834041
transform -1 0 27888 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_111
timestamp 1486834041
transform 1 0 672 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1486834041
transform -1 0 27888 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_112
timestamp 1486834041
transform 1 0 672 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1486834041
transform -1 0 27888 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_113
timestamp 1486834041
transform 1 0 672 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1486834041
transform -1 0 27888 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_114
timestamp 1486834041
transform 1 0 672 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1486834041
transform -1 0 27888 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_115
timestamp 1486834041
transform 1 0 672 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1486834041
transform -1 0 27888 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_116
timestamp 1486834041
transform 1 0 672 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1486834041
transform -1 0 27888 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_117
timestamp 1486834041
transform 1 0 672 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1486834041
transform -1 0 27888 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_118
timestamp 1486834041
transform 1 0 672 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1486834041
transform -1 0 27888 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_119
timestamp 1486834041
transform 1 0 672 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1486834041
transform -1 0 27888 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_120
timestamp 1486834041
transform 1 0 672 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1486834041
transform -1 0 27888 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_121
timestamp 1486834041
transform 1 0 672 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1486834041
transform -1 0 27888 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_122
timestamp 1486834041
transform 1 0 672 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1486834041
transform -1 0 27888 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_123
timestamp 1486834041
transform 1 0 672 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1486834041
transform -1 0 27888 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_124
timestamp 1486834041
transform 1 0 672 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1486834041
transform -1 0 27888 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_125
timestamp 1486834041
transform 1 0 672 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1486834041
transform -1 0 27888 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_126
timestamp 1486834041
transform 1 0 672 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1486834041
transform -1 0 27888 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_127
timestamp 1486834041
transform 1 0 672 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1486834041
transform -1 0 27888 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_128
timestamp 1486834041
transform 1 0 672 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1486834041
transform -1 0 27888 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_129
timestamp 1486834041
transform 1 0 672 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1486834041
transform -1 0 27888 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_130
timestamp 1486834041
transform 1 0 672 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1486834041
transform -1 0 27888 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_131
timestamp 1486834041
transform 1 0 672 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1486834041
transform -1 0 27888 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_132
timestamp 1486834041
transform 1 0 672 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1486834041
transform -1 0 27888 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_133
timestamp 1486834041
transform 1 0 672 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1486834041
transform -1 0 27888 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_134
timestamp 1486834041
transform 1 0 672 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1486834041
transform -1 0 27888 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_135
timestamp 1486834041
transform 1 0 672 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1486834041
transform -1 0 27888 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_136
timestamp 1486834041
transform 1 0 672 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1486834041
transform -1 0 27888 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_137
timestamp 1486834041
transform 1 0 672 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1486834041
transform -1 0 27888 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_138
timestamp 1486834041
transform 1 0 672 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1486834041
transform -1 0 27888 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_139
timestamp 1486834041
transform 1 0 672 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1486834041
transform -1 0 27888 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_140
timestamp 1486834041
transform 1 0 672 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1486834041
transform -1 0 27888 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_141
timestamp 1486834041
transform 1 0 672 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1486834041
transform -1 0 27888 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1486834041
transform 1 0 4480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1486834041
transform 1 0 8288 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1486834041
transform 1 0 12096 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1486834041
transform 1 0 15904 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1486834041
transform 1 0 19712 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1486834041
transform 1 0 23520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1486834041
transform 1 0 27328 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_149
timestamp 1486834041
transform 1 0 8512 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_150
timestamp 1486834041
transform 1 0 16352 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_151
timestamp 1486834041
transform 1 0 24192 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_152
timestamp 1486834041
transform 1 0 4592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_153
timestamp 1486834041
transform 1 0 12432 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_154
timestamp 1486834041
transform 1 0 20272 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_155
timestamp 1486834041
transform 1 0 8512 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_156
timestamp 1486834041
transform 1 0 16352 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_157
timestamp 1486834041
transform 1 0 24192 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_158
timestamp 1486834041
transform 1 0 4592 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_159
timestamp 1486834041
transform 1 0 12432 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_160
timestamp 1486834041
transform 1 0 20272 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_161
timestamp 1486834041
transform 1 0 8512 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_162
timestamp 1486834041
transform 1 0 16352 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_163
timestamp 1486834041
transform 1 0 24192 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_164
timestamp 1486834041
transform 1 0 4592 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_165
timestamp 1486834041
transform 1 0 12432 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_166
timestamp 1486834041
transform 1 0 20272 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_167
timestamp 1486834041
transform 1 0 8512 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_168
timestamp 1486834041
transform 1 0 16352 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_169
timestamp 1486834041
transform 1 0 24192 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_170
timestamp 1486834041
transform 1 0 4592 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_171
timestamp 1486834041
transform 1 0 12432 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_172
timestamp 1486834041
transform 1 0 20272 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_173
timestamp 1486834041
transform 1 0 8512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_174
timestamp 1486834041
transform 1 0 16352 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_175
timestamp 1486834041
transform 1 0 24192 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_176
timestamp 1486834041
transform 1 0 4592 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_177
timestamp 1486834041
transform 1 0 12432 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_178
timestamp 1486834041
transform 1 0 20272 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_179
timestamp 1486834041
transform 1 0 8512 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_180
timestamp 1486834041
transform 1 0 16352 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_181
timestamp 1486834041
transform 1 0 24192 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_182
timestamp 1486834041
transform 1 0 4592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_183
timestamp 1486834041
transform 1 0 12432 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_184
timestamp 1486834041
transform 1 0 20272 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_185
timestamp 1486834041
transform 1 0 8512 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_186
timestamp 1486834041
transform 1 0 16352 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_187
timestamp 1486834041
transform 1 0 24192 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_188
timestamp 1486834041
transform 1 0 4592 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_189
timestamp 1486834041
transform 1 0 12432 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_190
timestamp 1486834041
transform 1 0 20272 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_191
timestamp 1486834041
transform 1 0 8512 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_192
timestamp 1486834041
transform 1 0 16352 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_193
timestamp 1486834041
transform 1 0 24192 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_194
timestamp 1486834041
transform 1 0 4592 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_195
timestamp 1486834041
transform 1 0 12432 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_196
timestamp 1486834041
transform 1 0 20272 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_197
timestamp 1486834041
transform 1 0 8512 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_198
timestamp 1486834041
transform 1 0 16352 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_199
timestamp 1486834041
transform 1 0 24192 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_200
timestamp 1486834041
transform 1 0 4592 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_201
timestamp 1486834041
transform 1 0 12432 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_202
timestamp 1486834041
transform 1 0 20272 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_203
timestamp 1486834041
transform 1 0 8512 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_204
timestamp 1486834041
transform 1 0 16352 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_205
timestamp 1486834041
transform 1 0 24192 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_206
timestamp 1486834041
transform 1 0 4592 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_207
timestamp 1486834041
transform 1 0 12432 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_208
timestamp 1486834041
transform 1 0 20272 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_209
timestamp 1486834041
transform 1 0 8512 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_210
timestamp 1486834041
transform 1 0 16352 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_211
timestamp 1486834041
transform 1 0 24192 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_212
timestamp 1486834041
transform 1 0 4592 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_213
timestamp 1486834041
transform 1 0 12432 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_214
timestamp 1486834041
transform 1 0 20272 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_215
timestamp 1486834041
transform 1 0 8512 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_216
timestamp 1486834041
transform 1 0 16352 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_217
timestamp 1486834041
transform 1 0 24192 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_218
timestamp 1486834041
transform 1 0 4592 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_219
timestamp 1486834041
transform 1 0 12432 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_220
timestamp 1486834041
transform 1 0 20272 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_221
timestamp 1486834041
transform 1 0 8512 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_222
timestamp 1486834041
transform 1 0 16352 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_223
timestamp 1486834041
transform 1 0 24192 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_224
timestamp 1486834041
transform 1 0 4592 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_225
timestamp 1486834041
transform 1 0 12432 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_226
timestamp 1486834041
transform 1 0 20272 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_227
timestamp 1486834041
transform 1 0 8512 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_228
timestamp 1486834041
transform 1 0 16352 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_229
timestamp 1486834041
transform 1 0 24192 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_230
timestamp 1486834041
transform 1 0 4592 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_231
timestamp 1486834041
transform 1 0 12432 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_232
timestamp 1486834041
transform 1 0 20272 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_233
timestamp 1486834041
transform 1 0 8512 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_234
timestamp 1486834041
transform 1 0 16352 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_235
timestamp 1486834041
transform 1 0 24192 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_236
timestamp 1486834041
transform 1 0 4592 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_237
timestamp 1486834041
transform 1 0 12432 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_238
timestamp 1486834041
transform 1 0 20272 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_239
timestamp 1486834041
transform 1 0 8512 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_240
timestamp 1486834041
transform 1 0 16352 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_241
timestamp 1486834041
transform 1 0 24192 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1486834041
transform 1 0 4592 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1486834041
transform 1 0 12432 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_244
timestamp 1486834041
transform 1 0 20272 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1486834041
transform 1 0 8512 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1486834041
transform 1 0 16352 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1486834041
transform 1 0 24192 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1486834041
transform 1 0 4592 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1486834041
transform 1 0 12432 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1486834041
transform 1 0 20272 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_251
timestamp 1486834041
transform 1 0 8512 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_252
timestamp 1486834041
transform 1 0 16352 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1486834041
transform 1 0 24192 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_254
timestamp 1486834041
transform 1 0 4592 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_255
timestamp 1486834041
transform 1 0 12432 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_256
timestamp 1486834041
transform 1 0 20272 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_257
timestamp 1486834041
transform 1 0 8512 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_258
timestamp 1486834041
transform 1 0 16352 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_259
timestamp 1486834041
transform 1 0 24192 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_260
timestamp 1486834041
transform 1 0 4592 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_261
timestamp 1486834041
transform 1 0 12432 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_262
timestamp 1486834041
transform 1 0 20272 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_263
timestamp 1486834041
transform 1 0 8512 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_264
timestamp 1486834041
transform 1 0 16352 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_265
timestamp 1486834041
transform 1 0 24192 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_266
timestamp 1486834041
transform 1 0 4592 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_267
timestamp 1486834041
transform 1 0 12432 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_268
timestamp 1486834041
transform 1 0 20272 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_269
timestamp 1486834041
transform 1 0 8512 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_270
timestamp 1486834041
transform 1 0 16352 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_271
timestamp 1486834041
transform 1 0 24192 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_272
timestamp 1486834041
transform 1 0 4592 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_273
timestamp 1486834041
transform 1 0 12432 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_274
timestamp 1486834041
transform 1 0 20272 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_275
timestamp 1486834041
transform 1 0 8512 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_276
timestamp 1486834041
transform 1 0 16352 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_277
timestamp 1486834041
transform 1 0 24192 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_278
timestamp 1486834041
transform 1 0 4592 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_279
timestamp 1486834041
transform 1 0 12432 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_280
timestamp 1486834041
transform 1 0 20272 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_281
timestamp 1486834041
transform 1 0 8512 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_282
timestamp 1486834041
transform 1 0 16352 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_283
timestamp 1486834041
transform 1 0 24192 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_284
timestamp 1486834041
transform 1 0 4592 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_285
timestamp 1486834041
transform 1 0 12432 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_286
timestamp 1486834041
transform 1 0 20272 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_287
timestamp 1486834041
transform 1 0 8512 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_288
timestamp 1486834041
transform 1 0 16352 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_289
timestamp 1486834041
transform 1 0 24192 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_290
timestamp 1486834041
transform 1 0 4592 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_291
timestamp 1486834041
transform 1 0 12432 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_292
timestamp 1486834041
transform 1 0 20272 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_293
timestamp 1486834041
transform 1 0 8512 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_294
timestamp 1486834041
transform 1 0 16352 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_295
timestamp 1486834041
transform 1 0 24192 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_296
timestamp 1486834041
transform 1 0 4592 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_297
timestamp 1486834041
transform 1 0 12432 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_298
timestamp 1486834041
transform 1 0 20272 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_299
timestamp 1486834041
transform 1 0 8512 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_300
timestamp 1486834041
transform 1 0 16352 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_301
timestamp 1486834041
transform 1 0 24192 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_302
timestamp 1486834041
transform 1 0 4592 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_303
timestamp 1486834041
transform 1 0 12432 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_304
timestamp 1486834041
transform 1 0 20272 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_305
timestamp 1486834041
transform 1 0 8512 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_306
timestamp 1486834041
transform 1 0 16352 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_307
timestamp 1486834041
transform 1 0 24192 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_308
timestamp 1486834041
transform 1 0 4592 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_309
timestamp 1486834041
transform 1 0 12432 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_310
timestamp 1486834041
transform 1 0 20272 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_311
timestamp 1486834041
transform 1 0 8512 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_312
timestamp 1486834041
transform 1 0 16352 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_313
timestamp 1486834041
transform 1 0 24192 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_314
timestamp 1486834041
transform 1 0 4592 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_315
timestamp 1486834041
transform 1 0 12432 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_316
timestamp 1486834041
transform 1 0 20272 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_317
timestamp 1486834041
transform 1 0 8512 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_318
timestamp 1486834041
transform 1 0 16352 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_319
timestamp 1486834041
transform 1 0 24192 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_320
timestamp 1486834041
transform 1 0 4592 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_321
timestamp 1486834041
transform 1 0 12432 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_322
timestamp 1486834041
transform 1 0 20272 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_323
timestamp 1486834041
transform 1 0 8512 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_324
timestamp 1486834041
transform 1 0 16352 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_325
timestamp 1486834041
transform 1 0 24192 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_326
timestamp 1486834041
transform 1 0 4592 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_327
timestamp 1486834041
transform 1 0 12432 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_328
timestamp 1486834041
transform 1 0 20272 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_329
timestamp 1486834041
transform 1 0 8512 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_330
timestamp 1486834041
transform 1 0 16352 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_331
timestamp 1486834041
transform 1 0 24192 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_332
timestamp 1486834041
transform 1 0 4592 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_333
timestamp 1486834041
transform 1 0 12432 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_334
timestamp 1486834041
transform 1 0 20272 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_335
timestamp 1486834041
transform 1 0 8512 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_336
timestamp 1486834041
transform 1 0 16352 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_337
timestamp 1486834041
transform 1 0 24192 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_338
timestamp 1486834041
transform 1 0 4592 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_339
timestamp 1486834041
transform 1 0 12432 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_340
timestamp 1486834041
transform 1 0 20272 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_341
timestamp 1486834041
transform 1 0 8512 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_342
timestamp 1486834041
transform 1 0 16352 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_343
timestamp 1486834041
transform 1 0 24192 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_344
timestamp 1486834041
transform 1 0 4592 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_345
timestamp 1486834041
transform 1 0 12432 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_346
timestamp 1486834041
transform 1 0 20272 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_347
timestamp 1486834041
transform 1 0 8512 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_348
timestamp 1486834041
transform 1 0 16352 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_349
timestamp 1486834041
transform 1 0 24192 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_350
timestamp 1486834041
transform 1 0 4592 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_351
timestamp 1486834041
transform 1 0 12432 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_352
timestamp 1486834041
transform 1 0 20272 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_353
timestamp 1486834041
transform 1 0 8512 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_354
timestamp 1486834041
transform 1 0 16352 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_355
timestamp 1486834041
transform 1 0 24192 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_356
timestamp 1486834041
transform 1 0 4480 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_357
timestamp 1486834041
transform 1 0 8288 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_358
timestamp 1486834041
transform 1 0 12096 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_359
timestamp 1486834041
transform 1 0 15904 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_360
timestamp 1486834041
transform 1 0 19712 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_361
timestamp 1486834041
transform 1 0 23520 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_362
timestamp 1486834041
transform 1 0 27328 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  wire211
timestamp 1486834041
transform -1 0 17248 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  wire212
timestamp 1486834041
transform -1 0 14560 0 1 14896
box -86 -86 758 870
<< labels >>
flabel metal3 s 0 3136 112 3248 0 FreeSans 448 0 0 0 A_I_top
port 0 nsew signal output
flabel metal3 s 0 2240 112 2352 0 FreeSans 448 0 0 0 A_O_top
port 1 nsew signal input
flabel metal3 s 0 4032 112 4144 0 FreeSans 448 0 0 0 A_T_top
port 2 nsew signal output
flabel metal3 s 0 12992 112 13104 0 FreeSans 448 0 0 0 A_config_C_bit0
port 3 nsew signal output
flabel metal3 s 0 13888 112 14000 0 FreeSans 448 0 0 0 A_config_C_bit1
port 4 nsew signal output
flabel metal3 s 0 14784 112 14896 0 FreeSans 448 0 0 0 A_config_C_bit2
port 5 nsew signal output
flabel metal3 s 0 15680 112 15792 0 FreeSans 448 0 0 0 A_config_C_bit3
port 6 nsew signal output
flabel metal3 s 0 5824 112 5936 0 FreeSans 448 0 0 0 B_I_top
port 7 nsew signal output
flabel metal3 s 0 4928 112 5040 0 FreeSans 448 0 0 0 B_O_top
port 8 nsew signal input
flabel metal3 s 0 6720 112 6832 0 FreeSans 448 0 0 0 B_T_top
port 9 nsew signal output
flabel metal3 s 0 16576 112 16688 0 FreeSans 448 0 0 0 B_config_C_bit0
port 10 nsew signal output
flabel metal3 s 0 17472 112 17584 0 FreeSans 448 0 0 0 B_config_C_bit1
port 11 nsew signal output
flabel metal3 s 0 18368 112 18480 0 FreeSans 448 0 0 0 B_config_C_bit2
port 12 nsew signal output
flabel metal3 s 0 19264 112 19376 0 FreeSans 448 0 0 0 B_config_C_bit3
port 13 nsew signal output
flabel metal3 s 0 8512 112 8624 0 FreeSans 448 0 0 0 C_I_top
port 14 nsew signal output
flabel metal3 s 0 7616 112 7728 0 FreeSans 448 0 0 0 C_O_top
port 15 nsew signal input
flabel metal3 s 0 9408 112 9520 0 FreeSans 448 0 0 0 C_T_top
port 16 nsew signal output
flabel metal3 s 0 20160 112 20272 0 FreeSans 448 0 0 0 C_config_C_bit0
port 17 nsew signal output
flabel metal3 s 0 21056 112 21168 0 FreeSans 448 0 0 0 C_config_C_bit1
port 18 nsew signal output
flabel metal3 s 0 21952 112 22064 0 FreeSans 448 0 0 0 C_config_C_bit2
port 19 nsew signal output
flabel metal3 s 0 22848 112 22960 0 FreeSans 448 0 0 0 C_config_C_bit3
port 20 nsew signal output
flabel metal3 s 0 11200 112 11312 0 FreeSans 448 0 0 0 D_I_top
port 21 nsew signal output
flabel metal3 s 0 10304 112 10416 0 FreeSans 448 0 0 0 D_O_top
port 22 nsew signal input
flabel metal3 s 0 12096 112 12208 0 FreeSans 448 0 0 0 D_T_top
port 23 nsew signal output
flabel metal3 s 0 23744 112 23856 0 FreeSans 448 0 0 0 D_config_C_bit0
port 24 nsew signal output
flabel metal3 s 0 24640 112 24752 0 FreeSans 448 0 0 0 D_config_C_bit1
port 25 nsew signal output
flabel metal3 s 0 25536 112 25648 0 FreeSans 448 0 0 0 D_config_C_bit2
port 26 nsew signal output
flabel metal3 s 0 26432 112 26544 0 FreeSans 448 0 0 0 D_config_C_bit3
port 27 nsew signal output
flabel metal3 s 28448 21728 28560 21840 0 FreeSans 448 0 0 0 E1BEG[0]
port 28 nsew signal output
flabel metal3 s 28448 22176 28560 22288 0 FreeSans 448 0 0 0 E1BEG[1]
port 29 nsew signal output
flabel metal3 s 28448 22624 28560 22736 0 FreeSans 448 0 0 0 E1BEG[2]
port 30 nsew signal output
flabel metal3 s 28448 23072 28560 23184 0 FreeSans 448 0 0 0 E1BEG[3]
port 31 nsew signal output
flabel metal3 s 28448 23520 28560 23632 0 FreeSans 448 0 0 0 E2BEG[0]
port 32 nsew signal output
flabel metal3 s 28448 23968 28560 24080 0 FreeSans 448 0 0 0 E2BEG[1]
port 33 nsew signal output
flabel metal3 s 28448 24416 28560 24528 0 FreeSans 448 0 0 0 E2BEG[2]
port 34 nsew signal output
flabel metal3 s 28448 24864 28560 24976 0 FreeSans 448 0 0 0 E2BEG[3]
port 35 nsew signal output
flabel metal3 s 28448 25312 28560 25424 0 FreeSans 448 0 0 0 E2BEG[4]
port 36 nsew signal output
flabel metal3 s 28448 25760 28560 25872 0 FreeSans 448 0 0 0 E2BEG[5]
port 37 nsew signal output
flabel metal3 s 28448 26208 28560 26320 0 FreeSans 448 0 0 0 E2BEG[6]
port 38 nsew signal output
flabel metal3 s 28448 26656 28560 26768 0 FreeSans 448 0 0 0 E2BEG[7]
port 39 nsew signal output
flabel metal3 s 28448 27104 28560 27216 0 FreeSans 448 0 0 0 E2BEGb[0]
port 40 nsew signal output
flabel metal3 s 28448 27552 28560 27664 0 FreeSans 448 0 0 0 E2BEGb[1]
port 41 nsew signal output
flabel metal3 s 28448 28000 28560 28112 0 FreeSans 448 0 0 0 E2BEGb[2]
port 42 nsew signal output
flabel metal3 s 28448 28448 28560 28560 0 FreeSans 448 0 0 0 E2BEGb[3]
port 43 nsew signal output
flabel metal3 s 28448 28896 28560 29008 0 FreeSans 448 0 0 0 E2BEGb[4]
port 44 nsew signal output
flabel metal3 s 28448 29344 28560 29456 0 FreeSans 448 0 0 0 E2BEGb[5]
port 45 nsew signal output
flabel metal3 s 28448 29792 28560 29904 0 FreeSans 448 0 0 0 E2BEGb[6]
port 46 nsew signal output
flabel metal3 s 28448 30240 28560 30352 0 FreeSans 448 0 0 0 E2BEGb[7]
port 47 nsew signal output
flabel metal3 s 28448 37856 28560 37968 0 FreeSans 448 0 0 0 E6BEG[0]
port 48 nsew signal output
flabel metal3 s 28448 42336 28560 42448 0 FreeSans 448 0 0 0 E6BEG[10]
port 49 nsew signal output
flabel metal3 s 28448 42784 28560 42896 0 FreeSans 448 0 0 0 E6BEG[11]
port 50 nsew signal output
flabel metal3 s 28448 38304 28560 38416 0 FreeSans 448 0 0 0 E6BEG[1]
port 51 nsew signal output
flabel metal3 s 28448 38752 28560 38864 0 FreeSans 448 0 0 0 E6BEG[2]
port 52 nsew signal output
flabel metal3 s 28448 39200 28560 39312 0 FreeSans 448 0 0 0 E6BEG[3]
port 53 nsew signal output
flabel metal3 s 28448 39648 28560 39760 0 FreeSans 448 0 0 0 E6BEG[4]
port 54 nsew signal output
flabel metal3 s 28448 40096 28560 40208 0 FreeSans 448 0 0 0 E6BEG[5]
port 55 nsew signal output
flabel metal3 s 28448 40544 28560 40656 0 FreeSans 448 0 0 0 E6BEG[6]
port 56 nsew signal output
flabel metal3 s 28448 40992 28560 41104 0 FreeSans 448 0 0 0 E6BEG[7]
port 57 nsew signal output
flabel metal3 s 28448 41440 28560 41552 0 FreeSans 448 0 0 0 E6BEG[8]
port 58 nsew signal output
flabel metal3 s 28448 41888 28560 42000 0 FreeSans 448 0 0 0 E6BEG[9]
port 59 nsew signal output
flabel metal3 s 28448 30688 28560 30800 0 FreeSans 448 0 0 0 EE4BEG[0]
port 60 nsew signal output
flabel metal3 s 28448 35168 28560 35280 0 FreeSans 448 0 0 0 EE4BEG[10]
port 61 nsew signal output
flabel metal3 s 28448 35616 28560 35728 0 FreeSans 448 0 0 0 EE4BEG[11]
port 62 nsew signal output
flabel metal3 s 28448 36064 28560 36176 0 FreeSans 448 0 0 0 EE4BEG[12]
port 63 nsew signal output
flabel metal3 s 28448 36512 28560 36624 0 FreeSans 448 0 0 0 EE4BEG[13]
port 64 nsew signal output
flabel metal3 s 28448 36960 28560 37072 0 FreeSans 448 0 0 0 EE4BEG[14]
port 65 nsew signal output
flabel metal3 s 28448 37408 28560 37520 0 FreeSans 448 0 0 0 EE4BEG[15]
port 66 nsew signal output
flabel metal3 s 28448 31136 28560 31248 0 FreeSans 448 0 0 0 EE4BEG[1]
port 67 nsew signal output
flabel metal3 s 28448 31584 28560 31696 0 FreeSans 448 0 0 0 EE4BEG[2]
port 68 nsew signal output
flabel metal3 s 28448 32032 28560 32144 0 FreeSans 448 0 0 0 EE4BEG[3]
port 69 nsew signal output
flabel metal3 s 28448 32480 28560 32592 0 FreeSans 448 0 0 0 EE4BEG[4]
port 70 nsew signal output
flabel metal3 s 28448 32928 28560 33040 0 FreeSans 448 0 0 0 EE4BEG[5]
port 71 nsew signal output
flabel metal3 s 28448 33376 28560 33488 0 FreeSans 448 0 0 0 EE4BEG[6]
port 72 nsew signal output
flabel metal3 s 28448 33824 28560 33936 0 FreeSans 448 0 0 0 EE4BEG[7]
port 73 nsew signal output
flabel metal3 s 28448 34272 28560 34384 0 FreeSans 448 0 0 0 EE4BEG[8]
port 74 nsew signal output
flabel metal3 s 28448 34720 28560 34832 0 FreeSans 448 0 0 0 EE4BEG[9]
port 75 nsew signal output
flabel metal3 s 0 27328 112 27440 0 FreeSans 448 0 0 0 FrameData[0]
port 76 nsew signal input
flabel metal3 s 0 36288 112 36400 0 FreeSans 448 0 0 0 FrameData[10]
port 77 nsew signal input
flabel metal3 s 0 37184 112 37296 0 FreeSans 448 0 0 0 FrameData[11]
port 78 nsew signal input
flabel metal3 s 0 38080 112 38192 0 FreeSans 448 0 0 0 FrameData[12]
port 79 nsew signal input
flabel metal3 s 0 38976 112 39088 0 FreeSans 448 0 0 0 FrameData[13]
port 80 nsew signal input
flabel metal3 s 0 39872 112 39984 0 FreeSans 448 0 0 0 FrameData[14]
port 81 nsew signal input
flabel metal3 s 0 40768 112 40880 0 FreeSans 448 0 0 0 FrameData[15]
port 82 nsew signal input
flabel metal3 s 0 41664 112 41776 0 FreeSans 448 0 0 0 FrameData[16]
port 83 nsew signal input
flabel metal3 s 0 42560 112 42672 0 FreeSans 448 0 0 0 FrameData[17]
port 84 nsew signal input
flabel metal3 s 0 43456 112 43568 0 FreeSans 448 0 0 0 FrameData[18]
port 85 nsew signal input
flabel metal3 s 0 44352 112 44464 0 FreeSans 448 0 0 0 FrameData[19]
port 86 nsew signal input
flabel metal3 s 0 28224 112 28336 0 FreeSans 448 0 0 0 FrameData[1]
port 87 nsew signal input
flabel metal3 s 0 45248 112 45360 0 FreeSans 448 0 0 0 FrameData[20]
port 88 nsew signal input
flabel metal3 s 0 46144 112 46256 0 FreeSans 448 0 0 0 FrameData[21]
port 89 nsew signal input
flabel metal3 s 0 47040 112 47152 0 FreeSans 448 0 0 0 FrameData[22]
port 90 nsew signal input
flabel metal3 s 0 47936 112 48048 0 FreeSans 448 0 0 0 FrameData[23]
port 91 nsew signal input
flabel metal3 s 0 48832 112 48944 0 FreeSans 448 0 0 0 FrameData[24]
port 92 nsew signal input
flabel metal3 s 0 49728 112 49840 0 FreeSans 448 0 0 0 FrameData[25]
port 93 nsew signal input
flabel metal3 s 0 50624 112 50736 0 FreeSans 448 0 0 0 FrameData[26]
port 94 nsew signal input
flabel metal3 s 0 51520 112 51632 0 FreeSans 448 0 0 0 FrameData[27]
port 95 nsew signal input
flabel metal3 s 0 52416 112 52528 0 FreeSans 448 0 0 0 FrameData[28]
port 96 nsew signal input
flabel metal3 s 0 53312 112 53424 0 FreeSans 448 0 0 0 FrameData[29]
port 97 nsew signal input
flabel metal3 s 0 29120 112 29232 0 FreeSans 448 0 0 0 FrameData[2]
port 98 nsew signal input
flabel metal3 s 0 54208 112 54320 0 FreeSans 448 0 0 0 FrameData[30]
port 99 nsew signal input
flabel metal3 s 0 55104 112 55216 0 FreeSans 448 0 0 0 FrameData[31]
port 100 nsew signal input
flabel metal3 s 0 30016 112 30128 0 FreeSans 448 0 0 0 FrameData[3]
port 101 nsew signal input
flabel metal3 s 0 30912 112 31024 0 FreeSans 448 0 0 0 FrameData[4]
port 102 nsew signal input
flabel metal3 s 0 31808 112 31920 0 FreeSans 448 0 0 0 FrameData[5]
port 103 nsew signal input
flabel metal3 s 0 32704 112 32816 0 FreeSans 448 0 0 0 FrameData[6]
port 104 nsew signal input
flabel metal3 s 0 33600 112 33712 0 FreeSans 448 0 0 0 FrameData[7]
port 105 nsew signal input
flabel metal3 s 0 34496 112 34608 0 FreeSans 448 0 0 0 FrameData[8]
port 106 nsew signal input
flabel metal3 s 0 35392 112 35504 0 FreeSans 448 0 0 0 FrameData[9]
port 107 nsew signal input
flabel metal3 s 28448 43232 28560 43344 0 FreeSans 448 0 0 0 FrameData_O[0]
port 108 nsew signal output
flabel metal3 s 28448 47712 28560 47824 0 FreeSans 448 0 0 0 FrameData_O[10]
port 109 nsew signal output
flabel metal3 s 28448 48160 28560 48272 0 FreeSans 448 0 0 0 FrameData_O[11]
port 110 nsew signal output
flabel metal3 s 28448 48608 28560 48720 0 FreeSans 448 0 0 0 FrameData_O[12]
port 111 nsew signal output
flabel metal3 s 28448 49056 28560 49168 0 FreeSans 448 0 0 0 FrameData_O[13]
port 112 nsew signal output
flabel metal3 s 28448 49504 28560 49616 0 FreeSans 448 0 0 0 FrameData_O[14]
port 113 nsew signal output
flabel metal3 s 28448 49952 28560 50064 0 FreeSans 448 0 0 0 FrameData_O[15]
port 114 nsew signal output
flabel metal3 s 28448 50400 28560 50512 0 FreeSans 448 0 0 0 FrameData_O[16]
port 115 nsew signal output
flabel metal3 s 28448 50848 28560 50960 0 FreeSans 448 0 0 0 FrameData_O[17]
port 116 nsew signal output
flabel metal3 s 28448 51296 28560 51408 0 FreeSans 448 0 0 0 FrameData_O[18]
port 117 nsew signal output
flabel metal3 s 28448 51744 28560 51856 0 FreeSans 448 0 0 0 FrameData_O[19]
port 118 nsew signal output
flabel metal3 s 28448 43680 28560 43792 0 FreeSans 448 0 0 0 FrameData_O[1]
port 119 nsew signal output
flabel metal3 s 28448 52192 28560 52304 0 FreeSans 448 0 0 0 FrameData_O[20]
port 120 nsew signal output
flabel metal3 s 28448 52640 28560 52752 0 FreeSans 448 0 0 0 FrameData_O[21]
port 121 nsew signal output
flabel metal3 s 28448 53088 28560 53200 0 FreeSans 448 0 0 0 FrameData_O[22]
port 122 nsew signal output
flabel metal3 s 28448 53536 28560 53648 0 FreeSans 448 0 0 0 FrameData_O[23]
port 123 nsew signal output
flabel metal3 s 28448 53984 28560 54096 0 FreeSans 448 0 0 0 FrameData_O[24]
port 124 nsew signal output
flabel metal3 s 28448 54432 28560 54544 0 FreeSans 448 0 0 0 FrameData_O[25]
port 125 nsew signal output
flabel metal3 s 28448 54880 28560 54992 0 FreeSans 448 0 0 0 FrameData_O[26]
port 126 nsew signal output
flabel metal3 s 28448 55328 28560 55440 0 FreeSans 448 0 0 0 FrameData_O[27]
port 127 nsew signal output
flabel metal3 s 28448 55776 28560 55888 0 FreeSans 448 0 0 0 FrameData_O[28]
port 128 nsew signal output
flabel metal3 s 28448 56224 28560 56336 0 FreeSans 448 0 0 0 FrameData_O[29]
port 129 nsew signal output
flabel metal3 s 28448 44128 28560 44240 0 FreeSans 448 0 0 0 FrameData_O[2]
port 130 nsew signal output
flabel metal3 s 28448 56672 28560 56784 0 FreeSans 448 0 0 0 FrameData_O[30]
port 131 nsew signal output
flabel metal3 s 28448 57120 28560 57232 0 FreeSans 448 0 0 0 FrameData_O[31]
port 132 nsew signal output
flabel metal3 s 28448 44576 28560 44688 0 FreeSans 448 0 0 0 FrameData_O[3]
port 133 nsew signal output
flabel metal3 s 28448 45024 28560 45136 0 FreeSans 448 0 0 0 FrameData_O[4]
port 134 nsew signal output
flabel metal3 s 28448 45472 28560 45584 0 FreeSans 448 0 0 0 FrameData_O[5]
port 135 nsew signal output
flabel metal3 s 28448 45920 28560 46032 0 FreeSans 448 0 0 0 FrameData_O[6]
port 136 nsew signal output
flabel metal3 s 28448 46368 28560 46480 0 FreeSans 448 0 0 0 FrameData_O[7]
port 137 nsew signal output
flabel metal3 s 28448 46816 28560 46928 0 FreeSans 448 0 0 0 FrameData_O[8]
port 138 nsew signal output
flabel metal3 s 28448 47264 28560 47376 0 FreeSans 448 0 0 0 FrameData_O[9]
port 139 nsew signal output
flabel metal2 s 2016 0 2128 112 0 FreeSans 448 0 0 0 FrameStrobe[0]
port 140 nsew signal input
flabel metal2 s 15456 0 15568 112 0 FreeSans 448 0 0 0 FrameStrobe[10]
port 141 nsew signal input
flabel metal2 s 16800 0 16912 112 0 FreeSans 448 0 0 0 FrameStrobe[11]
port 142 nsew signal input
flabel metal2 s 18144 0 18256 112 0 FreeSans 448 0 0 0 FrameStrobe[12]
port 143 nsew signal input
flabel metal2 s 19488 0 19600 112 0 FreeSans 448 0 0 0 FrameStrobe[13]
port 144 nsew signal input
flabel metal2 s 20832 0 20944 112 0 FreeSans 448 0 0 0 FrameStrobe[14]
port 145 nsew signal input
flabel metal2 s 22176 0 22288 112 0 FreeSans 448 0 0 0 FrameStrobe[15]
port 146 nsew signal input
flabel metal2 s 23520 0 23632 112 0 FreeSans 448 0 0 0 FrameStrobe[16]
port 147 nsew signal input
flabel metal2 s 24864 0 24976 112 0 FreeSans 448 0 0 0 FrameStrobe[17]
port 148 nsew signal input
flabel metal2 s 26208 0 26320 112 0 FreeSans 448 0 0 0 FrameStrobe[18]
port 149 nsew signal input
flabel metal2 s 27552 0 27664 112 0 FreeSans 448 0 0 0 FrameStrobe[19]
port 150 nsew signal input
flabel metal2 s 3360 0 3472 112 0 FreeSans 448 0 0 0 FrameStrobe[1]
port 151 nsew signal input
flabel metal2 s 4704 0 4816 112 0 FreeSans 448 0 0 0 FrameStrobe[2]
port 152 nsew signal input
flabel metal2 s 6048 0 6160 112 0 FreeSans 448 0 0 0 FrameStrobe[3]
port 153 nsew signal input
flabel metal2 s 7392 0 7504 112 0 FreeSans 448 0 0 0 FrameStrobe[4]
port 154 nsew signal input
flabel metal2 s 8736 0 8848 112 0 FreeSans 448 0 0 0 FrameStrobe[5]
port 155 nsew signal input
flabel metal2 s 10080 0 10192 112 0 FreeSans 448 0 0 0 FrameStrobe[6]
port 156 nsew signal input
flabel metal2 s 11424 0 11536 112 0 FreeSans 448 0 0 0 FrameStrobe[7]
port 157 nsew signal input
flabel metal2 s 12768 0 12880 112 0 FreeSans 448 0 0 0 FrameStrobe[8]
port 158 nsew signal input
flabel metal2 s 14112 0 14224 112 0 FreeSans 448 0 0 0 FrameStrobe[9]
port 159 nsew signal input
flabel metal2 s 2016 57344 2128 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[0]
port 160 nsew signal output
flabel metal2 s 15456 57344 15568 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[10]
port 161 nsew signal output
flabel metal2 s 16800 57344 16912 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[11]
port 162 nsew signal output
flabel metal2 s 18144 57344 18256 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[12]
port 163 nsew signal output
flabel metal2 s 19488 57344 19600 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[13]
port 164 nsew signal output
flabel metal2 s 20832 57344 20944 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[14]
port 165 nsew signal output
flabel metal2 s 22176 57344 22288 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[15]
port 166 nsew signal output
flabel metal2 s 23520 57344 23632 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[16]
port 167 nsew signal output
flabel metal2 s 24864 57344 24976 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[17]
port 168 nsew signal output
flabel metal2 s 26208 57344 26320 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[18]
port 169 nsew signal output
flabel metal2 s 27552 57344 27664 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[19]
port 170 nsew signal output
flabel metal2 s 3360 57344 3472 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[1]
port 171 nsew signal output
flabel metal2 s 4704 57344 4816 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[2]
port 172 nsew signal output
flabel metal2 s 6048 57344 6160 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[3]
port 173 nsew signal output
flabel metal2 s 7392 57344 7504 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[4]
port 174 nsew signal output
flabel metal2 s 8736 57344 8848 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[5]
port 175 nsew signal output
flabel metal2 s 10080 57344 10192 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[6]
port 176 nsew signal output
flabel metal2 s 11424 57344 11536 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[7]
port 177 nsew signal output
flabel metal2 s 12768 57344 12880 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[8]
port 178 nsew signal output
flabel metal2 s 14112 57344 14224 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[9]
port 179 nsew signal output
flabel metal2 s 672 0 784 112 0 FreeSans 448 0 0 0 UserCLK
port 180 nsew signal input
flabel metal2 s 672 57344 784 57456 0 FreeSans 448 0 0 0 UserCLKo
port 181 nsew signal output
flabel metal4 s 3776 0 4096 57456 0 FreeSans 1472 90 0 0 VDD
port 182 nsew power bidirectional
flabel metal4 s 3776 0 4096 56 0 FreeSans 368 0 0 0 VDD
port 182 nsew power bidirectional
flabel metal4 s 3776 57400 4096 57456 0 FreeSans 368 0 0 0 VDD
port 182 nsew power bidirectional
flabel metal4 s 23776 0 24096 57456 0 FreeSans 1472 90 0 0 VDD
port 182 nsew power bidirectional
flabel metal4 s 23776 0 24096 56 0 FreeSans 368 0 0 0 VDD
port 182 nsew power bidirectional
flabel metal4 s 23776 57400 24096 57456 0 FreeSans 368 0 0 0 VDD
port 182 nsew power bidirectional
flabel metal4 s 4436 0 4756 57456 0 FreeSans 1472 90 0 0 VSS
port 183 nsew ground bidirectional
flabel metal4 s 4436 0 4756 56 0 FreeSans 368 0 0 0 VSS
port 183 nsew ground bidirectional
flabel metal4 s 4436 57400 4756 57456 0 FreeSans 368 0 0 0 VSS
port 183 nsew ground bidirectional
flabel metal4 s 24436 0 24756 57456 0 FreeSans 1472 90 0 0 VSS
port 183 nsew ground bidirectional
flabel metal4 s 24436 0 24756 56 0 FreeSans 368 0 0 0 VSS
port 183 nsew ground bidirectional
flabel metal4 s 24436 57400 24756 57456 0 FreeSans 368 0 0 0 VSS
port 183 nsew ground bidirectional
flabel metal3 s 28448 224 28560 336 0 FreeSans 448 0 0 0 W1END[0]
port 184 nsew signal input
flabel metal3 s 28448 672 28560 784 0 FreeSans 448 0 0 0 W1END[1]
port 185 nsew signal input
flabel metal3 s 28448 1120 28560 1232 0 FreeSans 448 0 0 0 W1END[2]
port 186 nsew signal input
flabel metal3 s 28448 1568 28560 1680 0 FreeSans 448 0 0 0 W1END[3]
port 187 nsew signal input
flabel metal3 s 28448 5600 28560 5712 0 FreeSans 448 0 0 0 W2END[0]
port 188 nsew signal input
flabel metal3 s 28448 6048 28560 6160 0 FreeSans 448 0 0 0 W2END[1]
port 189 nsew signal input
flabel metal3 s 28448 6496 28560 6608 0 FreeSans 448 0 0 0 W2END[2]
port 190 nsew signal input
flabel metal3 s 28448 6944 28560 7056 0 FreeSans 448 0 0 0 W2END[3]
port 191 nsew signal input
flabel metal3 s 28448 7392 28560 7504 0 FreeSans 448 0 0 0 W2END[4]
port 192 nsew signal input
flabel metal3 s 28448 7840 28560 7952 0 FreeSans 448 0 0 0 W2END[5]
port 193 nsew signal input
flabel metal3 s 28448 8288 28560 8400 0 FreeSans 448 0 0 0 W2END[6]
port 194 nsew signal input
flabel metal3 s 28448 8736 28560 8848 0 FreeSans 448 0 0 0 W2END[7]
port 195 nsew signal input
flabel metal3 s 28448 2016 28560 2128 0 FreeSans 448 0 0 0 W2MID[0]
port 196 nsew signal input
flabel metal3 s 28448 2464 28560 2576 0 FreeSans 448 0 0 0 W2MID[1]
port 197 nsew signal input
flabel metal3 s 28448 2912 28560 3024 0 FreeSans 448 0 0 0 W2MID[2]
port 198 nsew signal input
flabel metal3 s 28448 3360 28560 3472 0 FreeSans 448 0 0 0 W2MID[3]
port 199 nsew signal input
flabel metal3 s 28448 3808 28560 3920 0 FreeSans 448 0 0 0 W2MID[4]
port 200 nsew signal input
flabel metal3 s 28448 4256 28560 4368 0 FreeSans 448 0 0 0 W2MID[5]
port 201 nsew signal input
flabel metal3 s 28448 4704 28560 4816 0 FreeSans 448 0 0 0 W2MID[6]
port 202 nsew signal input
flabel metal3 s 28448 5152 28560 5264 0 FreeSans 448 0 0 0 W2MID[7]
port 203 nsew signal input
flabel metal3 s 28448 16352 28560 16464 0 FreeSans 448 0 0 0 W6END[0]
port 204 nsew signal input
flabel metal3 s 28448 20832 28560 20944 0 FreeSans 448 0 0 0 W6END[10]
port 205 nsew signal input
flabel metal3 s 28448 21280 28560 21392 0 FreeSans 448 0 0 0 W6END[11]
port 206 nsew signal input
flabel metal3 s 28448 16800 28560 16912 0 FreeSans 448 0 0 0 W6END[1]
port 207 nsew signal input
flabel metal3 s 28448 17248 28560 17360 0 FreeSans 448 0 0 0 W6END[2]
port 208 nsew signal input
flabel metal3 s 28448 17696 28560 17808 0 FreeSans 448 0 0 0 W6END[3]
port 209 nsew signal input
flabel metal3 s 28448 18144 28560 18256 0 FreeSans 448 0 0 0 W6END[4]
port 210 nsew signal input
flabel metal3 s 28448 18592 28560 18704 0 FreeSans 448 0 0 0 W6END[5]
port 211 nsew signal input
flabel metal3 s 28448 19040 28560 19152 0 FreeSans 448 0 0 0 W6END[6]
port 212 nsew signal input
flabel metal3 s 28448 19488 28560 19600 0 FreeSans 448 0 0 0 W6END[7]
port 213 nsew signal input
flabel metal3 s 28448 19936 28560 20048 0 FreeSans 448 0 0 0 W6END[8]
port 214 nsew signal input
flabel metal3 s 28448 20384 28560 20496 0 FreeSans 448 0 0 0 W6END[9]
port 215 nsew signal input
flabel metal3 s 28448 9184 28560 9296 0 FreeSans 448 0 0 0 WW4END[0]
port 216 nsew signal input
flabel metal3 s 28448 13664 28560 13776 0 FreeSans 448 0 0 0 WW4END[10]
port 217 nsew signal input
flabel metal3 s 28448 14112 28560 14224 0 FreeSans 448 0 0 0 WW4END[11]
port 218 nsew signal input
flabel metal3 s 28448 14560 28560 14672 0 FreeSans 448 0 0 0 WW4END[12]
port 219 nsew signal input
flabel metal3 s 28448 15008 28560 15120 0 FreeSans 448 0 0 0 WW4END[13]
port 220 nsew signal input
flabel metal3 s 28448 15456 28560 15568 0 FreeSans 448 0 0 0 WW4END[14]
port 221 nsew signal input
flabel metal3 s 28448 15904 28560 16016 0 FreeSans 448 0 0 0 WW4END[15]
port 222 nsew signal input
flabel metal3 s 28448 9632 28560 9744 0 FreeSans 448 0 0 0 WW4END[1]
port 223 nsew signal input
flabel metal3 s 28448 10080 28560 10192 0 FreeSans 448 0 0 0 WW4END[2]
port 224 nsew signal input
flabel metal3 s 28448 10528 28560 10640 0 FreeSans 448 0 0 0 WW4END[3]
port 225 nsew signal input
flabel metal3 s 28448 10976 28560 11088 0 FreeSans 448 0 0 0 WW4END[4]
port 226 nsew signal input
flabel metal3 s 28448 11424 28560 11536 0 FreeSans 448 0 0 0 WW4END[5]
port 227 nsew signal input
flabel metal3 s 28448 11872 28560 11984 0 FreeSans 448 0 0 0 WW4END[6]
port 228 nsew signal input
flabel metal3 s 28448 12320 28560 12432 0 FreeSans 448 0 0 0 WW4END[7]
port 229 nsew signal input
flabel metal3 s 28448 12768 28560 12880 0 FreeSans 448 0 0 0 WW4END[8]
port 230 nsew signal input
flabel metal3 s 28448 13216 28560 13328 0 FreeSans 448 0 0 0 WW4END[9]
port 231 nsew signal input
rlabel metal1 14280 56448 14280 56448 0 VDD
rlabel metal1 14280 55664 14280 55664 0 VSS
rlabel metal3 686 3192 686 3192 0 A_I_top
rlabel metal3 574 2296 574 2296 0 A_O_top
rlabel metal3 798 4088 798 4088 0 A_T_top
rlabel metal2 3080 11088 3080 11088 0 A_config_C_bit0
rlabel metal2 1512 7980 1512 7980 0 A_config_C_bit1
rlabel metal3 1694 14840 1694 14840 0 A_config_C_bit2
rlabel metal3 1470 15736 1470 15736 0 A_config_C_bit3
rlabel metal3 1470 5880 1470 5880 0 B_I_top
rlabel metal2 1064 3864 1064 3864 0 B_O_top
rlabel metal3 798 6776 798 6776 0 B_T_top
rlabel metal3 2702 16632 2702 16632 0 B_config_C_bit0
rlabel metal2 1176 8008 1176 8008 0 B_config_C_bit1
rlabel metal3 1064 9240 1064 9240 0 B_config_C_bit2
rlabel metal3 630 19320 630 19320 0 B_config_C_bit3
rlabel metal2 1624 7112 1624 7112 0 C_I_top
rlabel metal3 686 7672 686 7672 0 C_O_top
rlabel metal3 1526 9464 1526 9464 0 C_T_top
rlabel metal3 2478 20216 2478 20216 0 C_config_C_bit0
rlabel metal3 854 21112 854 21112 0 C_config_C_bit1
rlabel metal3 798 22008 798 22008 0 C_config_C_bit2
rlabel metal2 5544 21560 5544 21560 0 C_config_C_bit3
rlabel metal3 1694 11256 1694 11256 0 D_I_top
rlabel metal2 5152 7448 5152 7448 0 D_O_top
rlabel metal2 1288 8232 1288 8232 0 D_T_top
rlabel metal3 574 23800 574 23800 0 D_config_C_bit0
rlabel metal2 3752 24360 3752 24360 0 D_config_C_bit1
rlabel metal2 5544 25256 5544 25256 0 D_config_C_bit2
rlabel metal3 686 26488 686 26488 0 D_config_C_bit3
rlabel metal2 25704 21952 25704 21952 0 E1BEG[0]
rlabel metal2 27160 21952 27160 21952 0 E1BEG[1]
rlabel metal3 27874 22680 27874 22680 0 E1BEG[2]
rlabel metal2 25704 23408 25704 23408 0 E1BEG[3]
rlabel metal2 27160 23408 27160 23408 0 E2BEG[0]
rlabel metal2 25592 24416 25592 24416 0 E2BEG[1]
rlabel metal3 27874 24472 27874 24472 0 E2BEG[2]
rlabel metal2 25704 25088 25704 25088 0 E2BEG[3]
rlabel metal2 27160 25088 27160 25088 0 E2BEG[4]
rlabel metal3 27874 25816 27874 25816 0 E2BEG[5]
rlabel metal2 25704 26544 25704 26544 0 E2BEG[6]
rlabel metal2 27272 26600 27272 26600 0 E2BEG[7]
rlabel metal2 25704 27552 25704 27552 0 E2BEGb[0]
rlabel metal2 27048 27384 27048 27384 0 E2BEGb[1]
rlabel metal2 27160 28000 27160 28000 0 E2BEGb[2]
rlabel metal3 27818 28504 27818 28504 0 E2BEGb[3]
rlabel metal3 27762 28952 27762 28952 0 E2BEGb[4]
rlabel metal3 27818 29400 27818 29400 0 E2BEGb[5]
rlabel metal3 27762 29848 27762 29848 0 E2BEGb[6]
rlabel metal3 27818 30296 27818 30296 0 E2BEGb[7]
rlabel metal3 27090 37912 27090 37912 0 E6BEG[0]
rlabel metal3 27090 42392 27090 42392 0 E6BEG[10]
rlabel metal3 27874 42840 27874 42840 0 E6BEG[11]
rlabel metal3 27874 38360 27874 38360 0 E6BEG[1]
rlabel metal3 27762 38808 27762 38808 0 E6BEG[2]
rlabel metal3 27090 39256 27090 39256 0 E6BEG[3]
rlabel metal3 27874 39704 27874 39704 0 E6BEG[4]
rlabel metal3 27090 40152 27090 40152 0 E6BEG[5]
rlabel metal3 27762 40600 27762 40600 0 E6BEG[6]
rlabel metal3 27090 41048 27090 41048 0 E6BEG[7]
rlabel metal3 27874 41496 27874 41496 0 E6BEG[8]
rlabel metal3 27706 41944 27706 41944 0 E6BEG[9]
rlabel metal2 25480 30800 25480 30800 0 EE4BEG[0]
rlabel metal3 27874 35224 27874 35224 0 EE4BEG[10]
rlabel metal3 27818 35672 27818 35672 0 EE4BEG[11]
rlabel metal2 25704 36176 25704 36176 0 EE4BEG[12]
rlabel metal3 27706 36568 27706 36568 0 EE4BEG[13]
rlabel metal2 25480 37072 25480 37072 0 EE4BEG[14]
rlabel metal3 27762 37464 27762 37464 0 EE4BEG[15]
rlabel metal3 27762 31192 27762 31192 0 EE4BEG[1]
rlabel metal3 27090 31640 27090 31640 0 EE4BEG[2]
rlabel metal3 27874 32088 27874 32088 0 EE4BEG[3]
rlabel metal3 27818 32536 27818 32536 0 EE4BEG[4]
rlabel metal2 25704 33040 25704 33040 0 EE4BEG[5]
rlabel metal3 27874 33432 27874 33432 0 EE4BEG[6]
rlabel metal2 25704 34048 25704 34048 0 EE4BEG[7]
rlabel metal3 27762 34328 27762 34328 0 EE4BEG[8]
rlabel metal3 27090 34776 27090 34776 0 EE4BEG[9]
rlabel metal3 126 27384 126 27384 0 FrameData[0]
rlabel metal2 840 41720 840 41720 0 FrameData[10]
rlabel metal2 784 42728 784 42728 0 FrameData[11]
rlabel metal3 1470 38136 1470 38136 0 FrameData[12]
rlabel metal3 238 39032 238 39032 0 FrameData[13]
rlabel metal3 1078 39928 1078 39928 0 FrameData[14]
rlabel metal3 966 40824 966 40824 0 FrameData[15]
rlabel metal3 1022 41720 1022 41720 0 FrameData[16]
rlabel metal3 630 42616 630 42616 0 FrameData[17]
rlabel metal3 518 43512 518 43512 0 FrameData[18]
rlabel metal3 630 44408 630 44408 0 FrameData[19]
rlabel metal3 1722 28280 1722 28280 0 FrameData[1]
rlabel metal3 518 45304 518 45304 0 FrameData[20]
rlabel metal3 1022 46200 1022 46200 0 FrameData[21]
rlabel metal3 574 47096 574 47096 0 FrameData[22]
rlabel metal3 574 47992 574 47992 0 FrameData[23]
rlabel metal3 574 48888 574 48888 0 FrameData[24]
rlabel metal3 574 49784 574 49784 0 FrameData[25]
rlabel metal3 518 50680 518 50680 0 FrameData[26]
rlabel metal3 574 51576 574 51576 0 FrameData[27]
rlabel metal3 574 52472 574 52472 0 FrameData[28]
rlabel metal3 574 53368 574 53368 0 FrameData[29]
rlabel metal3 574 29176 574 29176 0 FrameData[2]
rlabel metal3 574 54264 574 54264 0 FrameData[30]
rlabel metal3 574 55160 574 55160 0 FrameData[31]
rlabel metal3 574 30072 574 30072 0 FrameData[3]
rlabel metal3 574 30968 574 30968 0 FrameData[4]
rlabel metal3 518 31864 518 31864 0 FrameData[5]
rlabel metal3 966 32760 966 32760 0 FrameData[6]
rlabel metal2 1064 37352 1064 37352 0 FrameData[7]
rlabel metal3 630 34552 630 34552 0 FrameData[8]
rlabel metal2 952 41160 952 41160 0 FrameData[9]
rlabel metal3 27090 43288 27090 43288 0 FrameData_O[0]
rlabel metal3 27874 47768 27874 47768 0 FrameData_O[10]
rlabel metal3 27818 48216 27818 48216 0 FrameData_O[11]
rlabel metal3 27090 48664 27090 48664 0 FrameData_O[12]
rlabel metal3 27874 49112 27874 49112 0 FrameData_O[13]
rlabel metal3 27090 49560 27090 49560 0 FrameData_O[14]
rlabel metal3 27762 50008 27762 50008 0 FrameData_O[15]
rlabel metal3 27090 50456 27090 50456 0 FrameData_O[16]
rlabel metal3 27874 50904 27874 50904 0 FrameData_O[17]
rlabel metal3 27818 51352 27818 51352 0 FrameData_O[18]
rlabel metal3 27090 51800 27090 51800 0 FrameData_O[19]
rlabel metal3 27762 43736 27762 43736 0 FrameData_O[1]
rlabel metal3 27874 52248 27874 52248 0 FrameData_O[20]
rlabel metal3 26978 52696 26978 52696 0 FrameData_O[21]
rlabel metal3 27762 53144 27762 53144 0 FrameData_O[22]
rlabel metal3 27090 53592 27090 53592 0 FrameData_O[23]
rlabel metal3 27874 54040 27874 54040 0 FrameData_O[24]
rlabel metal3 27090 54488 27090 54488 0 FrameData_O[25]
rlabel metal3 27314 54936 27314 54936 0 FrameData_O[26]
rlabel metal2 23576 54544 23576 54544 0 FrameData_O[27]
rlabel metal3 25074 55832 25074 55832 0 FrameData_O[28]
rlabel metal3 27370 56280 27370 56280 0 FrameData_O[29]
rlabel metal3 27090 44184 27090 44184 0 FrameData_O[2]
rlabel metal2 25760 51576 25760 51576 0 FrameData_O[30]
rlabel metal3 24360 52696 24360 52696 0 FrameData_O[31]
rlabel metal3 27874 44632 27874 44632 0 FrameData_O[3]
rlabel metal3 27818 45080 27818 45080 0 FrameData_O[4]
rlabel metal3 27090 45528 27090 45528 0 FrameData_O[5]
rlabel metal3 27874 45976 27874 45976 0 FrameData_O[6]
rlabel metal3 27090 46424 27090 46424 0 FrameData_O[7]
rlabel metal3 27762 46872 27762 46872 0 FrameData_O[8]
rlabel metal3 27090 47320 27090 47320 0 FrameData_O[9]
rlabel metal2 2072 2198 2072 2198 0 FrameStrobe[0]
rlabel metal2 27832 6636 27832 6636 0 FrameStrobe[10]
rlabel metal2 16856 854 16856 854 0 FrameStrobe[11]
rlabel metal2 26040 1624 26040 1624 0 FrameStrobe[12]
rlabel metal2 26936 1064 26936 1064 0 FrameStrobe[13]
rlabel metal2 20888 854 20888 854 0 FrameStrobe[14]
rlabel metal2 22232 1022 22232 1022 0 FrameStrobe[15]
rlabel metal2 23576 574 23576 574 0 FrameStrobe[16]
rlabel metal2 24920 238 24920 238 0 FrameStrobe[17]
rlabel metal2 26264 350 26264 350 0 FrameStrobe[18]
rlabel metal2 27608 1134 27608 1134 0 FrameStrobe[19]
rlabel metal2 3416 854 3416 854 0 FrameStrobe[1]
rlabel metal2 4760 238 4760 238 0 FrameStrobe[2]
rlabel metal2 6104 1638 6104 1638 0 FrameStrobe[3]
rlabel metal2 7448 518 7448 518 0 FrameStrobe[4]
rlabel metal3 20944 19320 20944 19320 0 FrameStrobe[5]
rlabel metal2 10136 518 10136 518 0 FrameStrobe[6]
rlabel metal2 11480 574 11480 574 0 FrameStrobe[7]
rlabel metal2 12824 686 12824 686 0 FrameStrobe[8]
rlabel metal2 14168 518 14168 518 0 FrameStrobe[9]
rlabel metal2 2520 55300 2520 55300 0 FrameStrobe_O[0]
rlabel metal3 16016 56280 16016 56280 0 FrameStrobe_O[10]
rlabel metal2 17304 55300 17304 55300 0 FrameStrobe_O[11]
rlabel metal2 18368 56280 18368 56280 0 FrameStrobe_O[12]
rlabel metal2 20328 56840 20328 56840 0 FrameStrobe_O[13]
rlabel metal2 20888 56826 20888 56826 0 FrameStrobe_O[14]
rlabel metal2 23016 56448 23016 56448 0 FrameStrobe_O[15]
rlabel metal2 23576 56826 23576 56826 0 FrameStrobe_O[16]
rlabel metal2 24920 56826 24920 56826 0 FrameStrobe_O[17]
rlabel metal2 26264 57330 26264 57330 0 FrameStrobe_O[18]
rlabel metal2 23800 52472 23800 52472 0 FrameStrobe_O[19]
rlabel metal2 3416 56826 3416 56826 0 FrameStrobe_O[1]
rlabel metal2 5208 56448 5208 56448 0 FrameStrobe_O[2]
rlabel metal3 6496 55160 6496 55160 0 FrameStrobe_O[3]
rlabel metal2 7448 56770 7448 56770 0 FrameStrobe_O[4]
rlabel metal2 9016 56448 9016 56448 0 FrameStrobe_O[5]
rlabel metal2 10584 56504 10584 56504 0 FrameStrobe_O[6]
rlabel metal3 11704 55160 11704 55160 0 FrameStrobe_O[7]
rlabel metal2 13048 56448 13048 56448 0 FrameStrobe_O[8]
rlabel metal2 14616 56504 14616 56504 0 FrameStrobe_O[9]
rlabel metal2 6888 39592 6888 39592 0 Inst_A_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 21560 29232 21560 29232 0 Inst_B_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 15512 16072 15512 16072 0 Inst_C_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 13608 19600 13608 19600 0 Inst_D_IO_1_bidirectional_frame_config_pass.Q
rlabel metal3 9184 34104 9184 34104 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 9128 34384 9128 34384 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit1.Q
rlabel metal3 16072 9576 16072 9576 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 18088 10752 18088 10752 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 19320 14560 19320 14560 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 16072 13832 16072 13832 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit13.Q
rlabel metal3 17528 12152 17528 12152 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 7784 14560 7784 14560 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit15.Q
rlabel metal3 2996 15288 2996 15288 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 7112 15512 7112 15512 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 18312 17528 18312 17528 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit18.Q
rlabel metal3 18928 17640 18928 17640 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 16352 40152 16352 40152 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 17304 17304 17304 17304 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 18760 16688 18760 16688 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 11144 10752 11144 10752 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 11480 11648 11480 11648 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 12040 11088 12040 11088 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 21000 15456 21000 15456 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q
rlabel metal3 21672 15288 21672 15288 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit26.Q
rlabel metal3 20160 15288 20160 15288 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 19544 13496 19544 13496 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 7784 10528 7784 10528 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 15512 39088 15512 39088 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit3.Q
rlabel metal3 8736 11480 8736 11480 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 9016 11704 9016 11704 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 18536 21336 18536 21336 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 19096 21728 19096 21728 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 19656 29176 19656 29176 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 19656 24304 19656 24304 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 16520 9632 16520 9632 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit8.Q
rlabel metal3 16016 7336 16016 7336 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 7448 25368 7448 25368 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit0.Q
rlabel metal3 8344 24696 8344 24696 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 13888 19208 13888 19208 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 12320 19320 12320 19320 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 4984 29904 4984 29904 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 3640 29512 3640 29512 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit13.Q
rlabel metal3 16016 30856 16016 30856 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 15848 31640 15848 31640 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 2856 23240 2856 23240 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 4032 23352 4032 23352 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit17.Q
rlabel metal3 21616 24136 21616 24136 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 22400 24696 22400 24696 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 3136 34888 3136 34888 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 10136 30240 10136 30240 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 9744 27608 9744 27608 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 21280 25704 21280 25704 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 19936 26488 19936 26488 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 9912 15736 9912 15736 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 8232 16576 8232 16576 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 16072 24976 16072 24976 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 14896 24696 14896 24696 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 2856 17696 2856 17696 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 3304 20132 3304 20132 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 4312 36008 4312 36008 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 12936 30128 12936 30128 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit30.Q
rlabel metal3 13104 30184 13104 30184 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 8120 37744 8120 37744 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 9464 39872 9464 39872 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 21000 31024 21000 31024 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit6.Q
rlabel metal3 20944 30968 20944 30968 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 12824 16576 12824 16576 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 16184 17136 16184 17136 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 7112 22400 7112 22400 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 8120 22232 8120 22232 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 14280 6944 14280 6944 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 14952 5544 14952 5544 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 2912 25480 2912 25480 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 4088 25368 4088 25368 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 1288 35336 1288 35336 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 2912 34104 2912 34104 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 6104 39032 6104 39032 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 7000 39200 7000 39200 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 20888 31080 20888 31080 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit18.Q
rlabel metal3 22456 30184 22456 30184 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 14728 33208 14728 33208 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 9072 26824 9072 26824 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 10696 25984 10696 25984 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 10808 21224 10808 21224 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 12040 21840 12040 21840 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit23.Q
rlabel metal3 13832 15288 13832 15288 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 16184 15568 16184 15568 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 14616 19320 14616 19320 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 12152 18704 12152 18704 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 2800 32760 2800 32760 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 3696 33320 3696 33320 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 15904 41720 15904 41720 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit3.Q
rlabel metal3 6832 29624 6832 29624 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit30.Q
rlabel metal3 4872 31192 4872 31192 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit31.Q
rlabel metal3 10696 38248 10696 38248 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 14280 39480 14280 39480 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 17752 28504 17752 28504 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 18984 27720 18984 27720 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 9632 9240 9632 9240 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 10864 7672 10864 7672 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit9.Q
rlabel metal3 13552 27272 13552 27272 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 15344 27272 15344 27272 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit11.Q
rlabel metal3 5040 19208 5040 19208 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit12.Q
rlabel metal2 6552 19936 6552 19936 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 5208 16632 5208 16632 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit14.Q
rlabel metal2 6552 17808 6552 17808 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit15.Q
rlabel metal3 5824 19992 5824 19992 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit16.Q
rlabel metal2 8456 20440 8456 20440 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit17.Q
rlabel metal3 13496 21560 13496 21560 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 16184 21840 16184 21840 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit19.Q
rlabel metal3 11536 28616 11536 28616 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 13048 28504 13048 28504 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit21.Q
rlabel metal3 16688 23352 16688 23352 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 18144 23912 18144 23912 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 9352 13776 9352 13776 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 10864 12264 10864 12264 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 14168 12656 14168 12656 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 13832 13384 13832 13384 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 4480 27048 4480 27048 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 3640 26768 3640 26768 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 3304 16184 3304 16184 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 2968 16968 2968 16968 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 12936 31976 12936 31976 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit4.Q
rlabel metal2 11760 31752 11760 31752 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit5.Q
rlabel metal2 18984 34608 18984 34608 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit6.Q
rlabel metal2 19880 35560 19880 35560 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 7672 19712 7672 19712 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 12936 24584 12936 24584 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit9.Q
rlabel metal3 11816 31864 11816 31864 0 Inst_W_IO4_switch_matrix.E1BEG0
rlabel metal2 19544 34552 19544 34552 0 Inst_W_IO4_switch_matrix.E1BEG1
rlabel metal3 12544 24136 12544 24136 0 Inst_W_IO4_switch_matrix.E1BEG2
rlabel metal3 14952 26264 14952 26264 0 Inst_W_IO4_switch_matrix.E1BEG3
rlabel metal2 5544 18592 5544 18592 0 Inst_W_IO4_switch_matrix.E2BEG0
rlabel metal3 7504 17752 7504 17752 0 Inst_W_IO4_switch_matrix.E2BEG1
rlabel metal2 8008 20328 8008 20328 0 Inst_W_IO4_switch_matrix.E2BEG2
rlabel metal2 15512 22680 15512 22680 0 Inst_W_IO4_switch_matrix.E2BEG3
rlabel metal2 12600 29008 12600 29008 0 Inst_W_IO4_switch_matrix.E2BEG4
rlabel metal2 17752 24304 17752 24304 0 Inst_W_IO4_switch_matrix.E2BEG5
rlabel metal2 9968 13608 9968 13608 0 Inst_W_IO4_switch_matrix.E2BEG6
rlabel metal2 15176 14224 15176 14224 0 Inst_W_IO4_switch_matrix.E2BEG7
rlabel metal3 4648 27272 4648 27272 0 Inst_W_IO4_switch_matrix.E2BEGb0
rlabel metal2 3416 17304 3416 17304 0 Inst_W_IO4_switch_matrix.E2BEGb1
rlabel metal2 7560 22176 7560 22176 0 Inst_W_IO4_switch_matrix.E2BEGb2
rlabel metal2 15456 29176 15456 29176 0 Inst_W_IO4_switch_matrix.E2BEGb3
rlabel metal3 13608 38696 13608 38696 0 Inst_W_IO4_switch_matrix.E2BEGb4
rlabel metal2 18536 27160 18536 27160 0 Inst_W_IO4_switch_matrix.E2BEGb5
rlabel metal2 10136 8288 10136 8288 0 Inst_W_IO4_switch_matrix.E2BEGb6
rlabel metal2 15400 5488 15400 5488 0 Inst_W_IO4_switch_matrix.E2BEGb7
rlabel metal2 4536 30240 4536 30240 0 Inst_W_IO4_switch_matrix.E6BEG0
rlabel metal2 16520 31304 16520 31304 0 Inst_W_IO4_switch_matrix.E6BEG1
rlabel metal2 9800 34440 9800 34440 0 Inst_W_IO4_switch_matrix.E6BEG10
rlabel metal2 16184 36848 16184 36848 0 Inst_W_IO4_switch_matrix.E6BEG11
rlabel metal2 1624 23352 1624 23352 0 Inst_W_IO4_switch_matrix.E6BEG2
rlabel metal2 21672 25032 21672 25032 0 Inst_W_IO4_switch_matrix.E6BEG3
rlabel metal2 11256 31024 11256 31024 0 Inst_W_IO4_switch_matrix.E6BEG4
rlabel metal2 20664 28280 20664 28280 0 Inst_W_IO4_switch_matrix.E6BEG5
rlabel metal2 10024 16352 10024 16352 0 Inst_W_IO4_switch_matrix.E6BEG6
rlabel metal2 15624 24304 15624 24304 0 Inst_W_IO4_switch_matrix.E6BEG7
rlabel metal3 2520 20888 2520 20888 0 Inst_W_IO4_switch_matrix.E6BEG8
rlabel metal2 13608 29848 13608 29848 0 Inst_W_IO4_switch_matrix.E6BEG9
rlabel metal3 4312 25704 4312 25704 0 Inst_W_IO4_switch_matrix.EE4BEG0
rlabel metal2 2128 33992 2128 33992 0 Inst_W_IO4_switch_matrix.EE4BEG1
rlabel metal2 8064 24584 8064 24584 0 Inst_W_IO4_switch_matrix.EE4BEG10
rlabel metal2 2632 35896 2632 35896 0 Inst_W_IO4_switch_matrix.EE4BEG11
rlabel metal2 9016 39144 9016 39144 0 Inst_W_IO4_switch_matrix.EE4BEG12
rlabel metal2 21672 31696 21672 31696 0 Inst_W_IO4_switch_matrix.EE4BEG13
rlabel metal2 15736 17192 15736 17192 0 Inst_W_IO4_switch_matrix.EE4BEG14
rlabel metal2 13496 20384 13496 20384 0 Inst_W_IO4_switch_matrix.EE4BEG15
rlabel metal2 7056 40152 7056 40152 0 Inst_W_IO4_switch_matrix.EE4BEG2
rlabel metal2 21280 31976 21280 31976 0 Inst_W_IO4_switch_matrix.EE4BEG3
rlabel metal3 10360 24696 10360 24696 0 Inst_W_IO4_switch_matrix.EE4BEG4
rlabel metal2 11368 21896 11368 21896 0 Inst_W_IO4_switch_matrix.EE4BEG5
rlabel metal2 15680 15176 15680 15176 0 Inst_W_IO4_switch_matrix.EE4BEG6
rlabel metal2 13832 21392 13832 21392 0 Inst_W_IO4_switch_matrix.EE4BEG7
rlabel metal2 3416 32984 3416 32984 0 Inst_W_IO4_switch_matrix.EE4BEG8
rlabel metal2 6048 30968 6048 30968 0 Inst_W_IO4_switch_matrix.EE4BEG9
rlabel metal2 728 350 728 350 0 UserCLK
rlabel metal2 13608 36008 13608 36008 0 UserCLK_regs
rlabel metal2 896 55944 896 55944 0 UserCLKo
rlabel metal3 27426 280 27426 280 0 W1END[0]
rlabel metal3 26922 728 26922 728 0 W1END[1]
rlabel metal3 27034 1176 27034 1176 0 W1END[2]
rlabel metal2 27160 1400 27160 1400 0 W1END[3]
rlabel metal3 27202 5656 27202 5656 0 W2END[0]
rlabel metal2 26712 6664 26712 6664 0 W2END[1]
rlabel metal2 26600 6608 26600 6608 0 W2END[2]
rlabel metal3 27986 7000 27986 7000 0 W2END[3]
rlabel metal3 27930 7448 27930 7448 0 W2END[4]
rlabel metal4 27496 7616 27496 7616 0 W2END[5]
rlabel metal3 27874 8344 27874 8344 0 W2END[6]
rlabel metal3 27202 8792 27202 8792 0 W2END[7]
rlabel metal3 27146 2072 27146 2072 0 W2MID[0]
rlabel metal3 27538 2520 27538 2520 0 W2MID[1]
rlabel metal3 27538 2968 27538 2968 0 W2MID[2]
rlabel metal2 27496 3080 27496 3080 0 W2MID[3]
rlabel metal3 27986 3864 27986 3864 0 W2MID[4]
rlabel metal3 27986 4312 27986 4312 0 W2MID[5]
rlabel metal3 27986 4760 27986 4760 0 W2MID[6]
rlabel metal3 27930 5208 27930 5208 0 W2MID[7]
rlabel metal2 27384 15848 27384 15848 0 W6END[0]
rlabel metal3 28042 20888 28042 20888 0 W6END[10]
rlabel metal2 27496 20664 27496 20664 0 W6END[11]
rlabel metal3 27538 16856 27538 16856 0 W6END[1]
rlabel metal3 28042 17304 28042 17304 0 W6END[2]
rlabel metal3 27538 17752 27538 17752 0 W6END[3]
rlabel metal2 27384 17528 27384 17528 0 W6END[4]
rlabel metal3 26740 18424 26740 18424 0 W6END[5]
rlabel metal3 28042 19096 28042 19096 0 W6END[6]
rlabel metal2 27384 18984 27384 18984 0 W6END[7]
rlabel metal2 25592 20440 25592 20440 0 W6END[8]
rlabel metal2 26600 20216 26600 20216 0 W6END[9]
rlabel metal2 25704 9520 25704 9520 0 WW4END[0]
rlabel metal3 27538 13720 27538 13720 0 WW4END[10]
rlabel metal3 27986 14168 27986 14168 0 WW4END[11]
rlabel metal2 27384 14168 27384 14168 0 WW4END[12]
rlabel metal3 27538 15064 27538 15064 0 WW4END[13]
rlabel metal2 27552 14728 27552 14728 0 WW4END[14]
rlabel metal2 26600 16016 26600 16016 0 WW4END[15]
rlabel metal2 26600 9744 26600 9744 0 WW4END[1]
rlabel metal2 26600 10248 26600 10248 0 WW4END[2]
rlabel metal3 28042 10584 28042 10584 0 WW4END[3]
rlabel metal2 26600 11200 26600 11200 0 WW4END[4]
rlabel metal2 27384 11032 27384 11032 0 WW4END[5]
rlabel metal3 27538 11928 27538 11928 0 WW4END[6]
rlabel metal3 28042 12376 28042 12376 0 WW4END[7]
rlabel metal2 26600 12880 26600 12880 0 WW4END[8]
rlabel metal2 27384 12712 27384 12712 0 WW4END[9]
rlabel metal2 18200 15960 18200 15960 0 _000_
rlabel metal2 9352 12040 9352 12040 0 _001_
rlabel metal2 16632 7728 16632 7728 0 _002_
rlabel metal2 15176 10024 15176 10024 0 _003_
rlabel metal2 15400 8120 15400 8120 0 _004_
rlabel metal2 3640 13832 3640 13832 0 _005_
rlabel metal2 12264 7952 12264 7952 0 _006_
rlabel metal2 8344 11704 8344 11704 0 _007_
rlabel metal2 17304 16128 17304 16128 0 _008_
rlabel metal2 19544 18032 19544 18032 0 _009_
rlabel metal2 17640 12208 17640 12208 0 _010_
rlabel metal2 19656 21672 19656 21672 0 _011_
rlabel metal2 15736 10472 15736 10472 0 _012_
rlabel metal3 16128 8232 16128 8232 0 _013_
rlabel metal3 16464 8008 16464 8008 0 _014_
rlabel metal3 17080 7672 17080 7672 0 _015_
rlabel metal2 17192 9968 17192 9968 0 _016_
rlabel metal2 15960 9016 15960 9016 0 _017_
rlabel metal2 17584 8344 17584 8344 0 _018_
rlabel metal3 8624 15848 8624 15848 0 _019_
rlabel metal2 7560 12936 7560 12936 0 _020_
rlabel metal3 6048 14280 6048 14280 0 _021_
rlabel metal2 7952 13160 7952 13160 0 _022_
rlabel metal3 8400 15176 8400 15176 0 _023_
rlabel metal3 7784 14840 7784 14840 0 _024_
rlabel metal3 8512 14504 8512 14504 0 _025_
rlabel metal2 12152 10696 12152 10696 0 _026_
rlabel metal2 12264 10472 12264 10472 0 _027_
rlabel metal2 12768 10024 12768 10024 0 _028_
rlabel metal2 13944 10304 13944 10304 0 _029_
rlabel metal2 10920 10752 10920 10752 0 _030_
rlabel metal2 10752 10472 10752 10472 0 _031_
rlabel metal3 12488 10360 12488 10360 0 _032_
rlabel metal2 7896 9856 7896 9856 0 _033_
rlabel metal2 7448 10304 7448 10304 0 _034_
rlabel metal2 7224 10864 7224 10864 0 _035_
rlabel metal3 8680 10584 8680 10584 0 _036_
rlabel metal3 8680 9128 8680 9128 0 _037_
rlabel metal2 8288 8008 8288 8008 0 _038_
rlabel metal3 8848 10360 8848 10360 0 _039_
rlabel metal2 20552 10248 20552 10248 0 _040_
rlabel metal3 20272 13496 20272 13496 0 _041_
rlabel metal2 20664 11872 20664 11872 0 _042_
rlabel metal2 20776 12488 20776 12488 0 _043_
rlabel metal3 20888 15176 20888 15176 0 _044_
rlabel metal2 19992 14504 19992 14504 0 _045_
rlabel metal2 16688 16072 16688 16072 0 _046_
rlabel metal2 18648 16352 18648 16352 0 _047_
rlabel metal2 17360 15848 17360 15848 0 _048_
rlabel metal2 17136 15624 17136 15624 0 _049_
rlabel metal2 19992 17472 19992 17472 0 _050_
rlabel metal2 18984 16576 18984 16576 0 _051_
rlabel metal2 19992 16576 19992 16576 0 _052_
rlabel metal2 19376 16856 19376 16856 0 _053_
rlabel metal2 17864 19096 17864 19096 0 _054_
rlabel metal3 18648 17080 18648 17080 0 _055_
rlabel metal3 18200 17752 18200 17752 0 _056_
rlabel metal3 17864 17080 17864 17080 0 _057_
rlabel metal3 18424 10024 18424 10024 0 _058_
rlabel metal3 18200 10696 18200 10696 0 _059_
rlabel metal2 18760 11648 18760 11648 0 _060_
rlabel metal2 19264 12152 19264 12152 0 _061_
rlabel metal2 18760 13832 18760 13832 0 _062_
rlabel metal2 18368 12376 18368 12376 0 _063_
rlabel metal2 16912 12152 16912 12152 0 _064_
rlabel metal3 17640 15288 17640 15288 0 _065_
rlabel metal2 17528 13720 17528 13720 0 _066_
rlabel metal2 17752 11984 17752 11984 0 _067_
rlabel metal2 20664 20160 20664 20160 0 _068_
rlabel metal3 21616 20104 21616 20104 0 _069_
rlabel metal2 19768 21336 19768 21336 0 _070_
rlabel metal2 19880 23128 19880 23128 0 _071_
rlabel metal2 20328 19656 20328 19656 0 _072_
rlabel metal2 19992 20160 19992 20160 0 _073_
rlabel metal3 18424 21000 18424 21000 0 _074_
rlabel metal2 17752 20440 17752 20440 0 _075_
rlabel metal3 18368 21560 18368 21560 0 _076_
rlabel metal3 20160 21336 20160 21336 0 _077_
rlabel metal2 14056 37296 14056 37296 0 clknet_0_UserCLK
rlabel metal2 14840 34048 14840 34048 0 clknet_0_UserCLK_regs
rlabel metal2 10584 38080 10584 38080 0 clknet_1_0__leaf_UserCLK
rlabel metal2 12600 32984 12600 32984 0 clknet_1_0__leaf_UserCLK_regs
rlabel metal3 9184 37240 9184 37240 0 clknet_1_1__leaf_UserCLK_regs
rlabel metal2 1624 3808 1624 3808 0 net1
rlabel metal2 2576 41048 2576 41048 0 net10
rlabel metal3 19208 17136 19208 17136 0 net100
rlabel metal2 7392 19208 7392 19208 0 net101
rlabel metal3 18200 12432 18200 12432 0 net102
rlabel metal3 21028 12040 21028 12040 0 net103
rlabel metal2 22008 9016 22008 9016 0 net104
rlabel metal2 17528 6160 17528 6160 0 net105
rlabel metal2 6888 15876 6888 15876 0 net106
rlabel metal2 2296 7728 2296 7728 0 net107
rlabel metal2 23688 13048 23688 13048 0 net108
rlabel metal2 17024 9240 17024 9240 0 net109
rlabel metal2 1736 15848 1736 15848 0 net11
rlabel metal2 17080 11704 17080 11704 0 net110
rlabel metal2 2016 5096 2016 5096 0 net111
rlabel metal3 6944 6104 6944 6104 0 net112
rlabel metal2 2408 7952 2408 7952 0 net113
rlabel metal2 2408 10304 2408 10304 0 net114
rlabel metal2 2408 12432 2408 12432 0 net115
rlabel metal2 14392 15624 14392 15624 0 net116
rlabel metal3 8736 7448 8736 7448 0 net117
rlabel metal3 4200 13608 4200 13608 0 net118
rlabel metal3 4368 12376 4368 12376 0 net119
rlabel metal3 2352 22456 2352 22456 0 net12
rlabel metal3 1792 11592 1792 11592 0 net120
rlabel metal2 5600 16408 5600 16408 0 net121
rlabel metal3 9912 13944 9912 13944 0 net122
rlabel metal2 2016 9352 2016 9352 0 net123
rlabel metal2 2352 23576 2352 23576 0 net124
rlabel metal2 4312 24612 4312 24612 0 net125
rlabel metal2 3864 38192 3864 38192 0 net126
rlabel metal2 2184 26180 2184 26180 0 net127
rlabel metal2 24976 22344 24976 22344 0 net128
rlabel metal3 24920 21560 24920 21560 0 net129
rlabel metal2 2744 23072 2744 23072 0 net13
rlabel metal3 18312 22624 18312 22624 0 net130
rlabel metal2 24696 24080 24696 24080 0 net131
rlabel metal4 18648 20776 18648 20776 0 net132
rlabel metal2 24920 23968 24920 23968 0 net133
rlabel metal4 20664 23408 20664 23408 0 net134
rlabel metal2 16072 24248 16072 24248 0 net135
rlabel metal2 26208 24696 26208 24696 0 net136
rlabel metal2 18816 24808 18816 24808 0 net137
rlabel metal2 24248 23156 24248 23156 0 net138
rlabel metal3 16072 17080 16072 17080 0 net139
rlabel metal3 8400 41216 8400 41216 0 net14
rlabel metal2 24920 27552 24920 27552 0 net140
rlabel metal3 4032 16968 4032 16968 0 net141
rlabel metal4 26264 26264 26264 26264 0 net142
rlabel metal3 21168 28616 21168 28616 0 net143
rlabel metal2 12768 40264 12768 40264 0 net144
rlabel metal3 22680 28504 22680 28504 0 net145
rlabel metal2 26264 30632 26264 30632 0 net146
rlabel metal3 27496 9352 27496 9352 0 net147
rlabel metal3 20104 36176 20104 36176 0 net148
rlabel metal2 24696 42672 24696 42672 0 net149
rlabel metal2 7448 39032 7448 39032 0 net15
rlabel metal3 25928 44296 25928 44296 0 net150
rlabel metal2 26264 39312 26264 39312 0 net151
rlabel metal2 1176 22680 1176 22680 0 net152
rlabel metal3 23520 39592 23520 39592 0 net153
rlabel metal2 26488 38080 26488 38080 0 net154
rlabel metal2 24472 40264 24472 40264 0 net155
rlabel metal3 21504 41832 21504 41832 0 net156
rlabel metal2 24808 40656 24808 40656 0 net157
rlabel metal2 1400 22792 1400 22792 0 net158
rlabel metal2 26152 42392 26152 42392 0 net159
rlabel metal2 7112 25424 7112 25424 0 net16
rlabel metal2 24808 31416 24808 31416 0 net160
rlabel metal2 26264 36176 26264 36176 0 net161
rlabel metal2 26152 36736 26152 36736 0 net162
rlabel metal2 9576 39816 9576 39816 0 net163
rlabel metal2 20776 35336 20776 35336 0 net164
rlabel metal2 15288 19376 15288 19376 0 net165
rlabel metal3 23128 38696 23128 38696 0 net166
rlabel metal2 1736 37240 1736 37240 0 net167
rlabel metal2 23688 34832 23688 34832 0 net168
rlabel metal3 24192 32648 24192 32648 0 net169
rlabel metal2 9464 19376 9464 19376 0 net17
rlabel metal2 26152 33376 26152 33376 0 net170
rlabel metal2 24920 32256 24920 32256 0 net171
rlabel metal2 17864 24584 17864 24584 0 net172
rlabel metal2 25032 34104 25032 34104 0 net173
rlabel metal2 26152 34944 26152 34944 0 net174
rlabel metal2 24696 34384 24696 34384 0 net175
rlabel metal2 24920 40880 24920 40880 0 net176
rlabel metal2 26264 48944 26264 48944 0 net177
rlabel metal2 26264 49448 26264 49448 0 net178
rlabel metal2 2184 18536 2184 18536 0 net179
rlabel metal2 2744 46536 2744 46536 0 net18
rlabel metal3 18536 50680 18536 50680 0 net180
rlabel metal3 16968 49672 16968 49672 0 net181
rlabel metal2 2912 21560 2912 21560 0 net182
rlabel metal2 24696 50512 24696 50512 0 net183
rlabel metal2 26264 52304 26264 52304 0 net184
rlabel metal2 27272 44408 27272 44408 0 net185
rlabel metal3 25760 52136 25760 52136 0 net186
rlabel metal3 17416 44968 17416 44968 0 net187
rlabel metal2 26264 53424 26264 53424 0 net188
rlabel metal3 18648 52808 18648 52808 0 net189
rlabel metal2 8344 41944 8344 41944 0 net19
rlabel metal2 26320 43848 26320 43848 0 net190
rlabel metal2 24696 53648 24696 53648 0 net191
rlabel metal3 26208 55272 26208 55272 0 net192
rlabel metal3 25144 55272 25144 55272 0 net193
rlabel metal3 22960 54488 22960 54488 0 net194
rlabel metal3 14672 46984 14672 46984 0 net195
rlabel metal2 20888 54544 20888 54544 0 net196
rlabel metal2 3192 13104 3192 13104 0 net197
rlabel metal3 22456 44296 22456 44296 0 net198
rlabel metal3 16240 51240 16240 51240 0 net199
rlabel metal3 952 2856 952 2856 0 net2
rlabel metal2 840 45864 840 45864 0 net20
rlabel metal2 23240 48300 23240 48300 0 net200
rlabel metal2 26040 45864 26040 45864 0 net201
rlabel metal2 26264 46312 26264 46312 0 net202
rlabel metal3 20216 45864 20216 45864 0 net203
rlabel metal3 24920 47376 24920 47376 0 net204
rlabel metal3 21336 46536 21336 46536 0 net205
rlabel metal2 26488 45948 26488 45948 0 net206
rlabel metal3 22008 47432 22008 47432 0 net207
rlabel metal3 5432 39704 5432 39704 0 net208
rlabel metal3 22120 37352 22120 37352 0 net209
rlabel metal3 6020 42504 6020 42504 0 net21
rlabel metal3 19432 55272 19432 55272 0 net210
rlabel metal2 26488 2240 26488 2240 0 net211
rlabel metal2 27496 2128 27496 2128 0 net212
rlabel metal2 21896 52248 21896 52248 0 net213
rlabel metal3 15904 2072 15904 2072 0 net214
rlabel metal2 22008 53816 22008 53816 0 net215
rlabel metal2 23576 51744 23576 51744 0 net216
rlabel metal2 24920 54208 24920 54208 0 net217
rlabel metal4 22792 29288 22792 29288 0 net218
rlabel metal2 3024 30072 3024 30072 0 net219
rlabel metal3 2016 50456 2016 50456 0 net22
rlabel metal2 6216 55888 6216 55888 0 net220
rlabel metal2 6328 49476 6328 49476 0 net221
rlabel metal2 8120 49392 8120 49392 0 net222
rlabel metal3 18480 39704 18480 39704 0 net223
rlabel metal3 16408 54488 16408 54488 0 net224
rlabel metal2 12824 49476 12824 49476 0 net225
rlabel metal3 16856 55944 16856 55944 0 net226
rlabel metal3 20832 41720 20832 41720 0 net227
rlabel metal2 1400 55552 1400 55552 0 net228
rlabel metal2 16520 7392 16520 7392 0 net229
rlabel metal3 3752 51240 3752 51240 0 net23
rlabel metal2 2184 7140 2184 7140 0 net230
rlabel metal2 9128 48720 9128 48720 0 net24
rlabel metal2 2688 24584 2688 24584 0 net25
rlabel metal2 1624 52584 1624 52584 0 net26
rlabel metal2 1624 30072 1624 30072 0 net27
rlabel metal2 1344 54600 1344 54600 0 net28
rlabel metal3 1008 22120 1008 22120 0 net29
rlabel metal2 3136 7000 3136 7000 0 net3
rlabel metal2 11816 39144 11816 39144 0 net30
rlabel metal2 16408 35392 16408 35392 0 net31
rlabel metal3 10528 41272 10528 41272 0 net32
rlabel metal2 2520 34496 2520 34496 0 net33
rlabel metal3 7112 38920 7112 38920 0 net34
rlabel metal3 1064 18480 1064 18480 0 net35
rlabel metal3 952 41048 952 41048 0 net36
rlabel metal2 3192 11760 3192 11760 0 net37
rlabel metal2 2072 10528 2072 10528 0 net38
rlabel metal2 3080 18816 3080 18816 0 net39
rlabel metal2 12040 24472 12040 24472 0 net4
rlabel metal3 2464 21672 2464 21672 0 net40
rlabel metal2 1400 16184 1400 16184 0 net41
rlabel metal2 17416 32032 17416 32032 0 net42
rlabel metal2 9352 22960 9352 22960 0 net43
rlabel metal3 2072 35784 2072 35784 0 net44
rlabel metal2 5432 39088 5432 39088 0 net45
rlabel metal2 3528 39424 3528 39424 0 net46
rlabel metal3 1792 28504 1792 28504 0 net47
rlabel metal3 17752 26376 17752 26376 0 net48
rlabel metal3 17472 31752 17472 31752 0 net49
rlabel metal3 6552 24080 6552 24080 0 net5
rlabel metal2 2632 29176 2632 29176 0 net50
rlabel metal2 14392 21560 14392 21560 0 net51
rlabel metal2 23128 16324 23128 16324 0 net52
rlabel metal3 9912 9016 9912 9016 0 net53
rlabel metal2 18088 29344 18088 29344 0 net54
rlabel metal2 7896 40432 7896 40432 0 net55
rlabel metal2 25704 1736 25704 1736 0 net56
rlabel metal2 24920 3584 24920 3584 0 net57
rlabel metal3 23464 1848 23464 1848 0 net58
rlabel metal2 26600 1344 26600 1344 0 net59
rlabel metal3 6440 41832 6440 41832 0 net6
rlabel metal3 23128 18424 23128 18424 0 net60
rlabel metal2 19544 8400 19544 8400 0 net61
rlabel metal3 18256 25928 18256 25928 0 net62
rlabel metal2 26936 7224 26936 7224 0 net63
rlabel metal3 16912 26712 16912 26712 0 net64
rlabel metal3 27608 7560 27608 7560 0 net65
rlabel metal2 1848 17530 1848 17530 0 net66
rlabel metal2 19544 20944 19544 20944 0 net67
rlabel metal2 20888 18144 20888 18144 0 net68
rlabel metal2 26152 3024 26152 3024 0 net69
rlabel metal2 1400 41328 1400 41328 0 net7
rlabel metal3 23688 15400 23688 15400 0 net70
rlabel metal2 27104 2856 27104 2856 0 net71
rlabel metal3 27272 3640 27272 3640 0 net72
rlabel metal2 18872 18256 18872 18256 0 net73
rlabel metal2 18032 9912 18032 9912 0 net74
rlabel metal2 17976 18256 17976 18256 0 net75
rlabel metal2 10024 25088 10024 25088 0 net76
rlabel metal2 2296 33488 2296 33488 0 net77
rlabel metal2 20944 23352 20944 23352 0 net78
rlabel metal2 11032 38752 11032 38752 0 net79
rlabel metal3 2016 23016 2016 23016 0 net8
rlabel metal2 17528 23800 17528 23800 0 net80
rlabel metal2 8232 39704 8232 39704 0 net81
rlabel metal2 2632 25088 2632 25088 0 net82
rlabel metal2 6104 40264 6104 40264 0 net83
rlabel metal3 21000 17696 21000 17696 0 net84
rlabel metal2 23240 31584 23240 31584 0 net85
rlabel metal3 22232 21728 22232 21728 0 net86
rlabel metal3 24416 19992 24416 19992 0 net87
rlabel metal3 15680 21000 15680 21000 0 net88
rlabel metal3 21448 23800 21448 23800 0 net89
rlabel metal4 2408 23072 2408 23072 0 net9
rlabel metal2 27104 12824 27104 12824 0 net90
rlabel metal3 27104 13832 27104 13832 0 net91
rlabel metal4 19656 15624 19656 15624 0 net92
rlabel metal2 2744 17696 2744 17696 0 net93
rlabel metal3 15848 18816 15848 18816 0 net94
rlabel metal2 26040 9408 26040 9408 0 net95
rlabel metal2 18760 22456 18760 22456 0 net96
rlabel metal3 27328 10920 27328 10920 0 net97
rlabel metal2 16464 21560 16464 21560 0 net98
rlabel metal2 27048 11648 27048 11648 0 net99
<< properties >>
string FIXED_BBOX 0 0 28560 57456
<< end >>
