VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO LUT4AB
  CLASS BLOCK ;
  FOREIGN LUT4AB ;
  ORIGIN 0.000 0.000 ;
  SIZE 287.280 BY 287.280 ;
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.015500 ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 0.000 120.400 0.560 ;
    END
  END Ci
  PIN Co
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 286.720 120.400 287.280 ;
    END
  END Co
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 108.640 287.280 109.200 ;
    END
  END E1BEG[0]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 110.880 287.280 111.440 ;
    END
  END E1BEG[1]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 113.120 287.280 113.680 ;
    END
  END E1BEG[2]
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 115.360 287.280 115.920 ;
    END
  END E1BEG[3]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.513500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 108.640 0.560 109.200 ;
    END
  END E1END[0]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.513500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 0.560 111.440 ;
    END
  END E1END[1]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.516500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 113.120 0.560 113.680 ;
    END
  END E1END[2]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.516500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 115.360 0.560 115.920 ;
    END
  END E1END[3]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 117.600 287.280 118.160 ;
    END
  END E2BEG[0]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 119.840 287.280 120.400 ;
    END
  END E2BEG[1]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 122.080 287.280 122.640 ;
    END
  END E2BEG[2]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 124.320 287.280 124.880 ;
    END
  END E2BEG[3]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 126.560 287.280 127.120 ;
    END
  END E2BEG[4]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 128.800 287.280 129.360 ;
    END
  END E2BEG[5]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 131.040 287.280 131.600 ;
    END
  END E2BEG[6]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 133.280 287.280 133.840 ;
    END
  END E2BEG[7]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 135.520 287.280 136.080 ;
    END
  END E2BEGb[0]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 137.760 287.280 138.320 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 140.000 287.280 140.560 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 142.240 287.280 142.800 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 144.480 287.280 145.040 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 146.720 287.280 147.280 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 148.960 287.280 149.520 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 151.200 287.280 151.760 ;
    END
  END E2BEGb[7]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.006000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 135.520 0.560 136.080 ;
    END
  END E2END[0]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.006000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 0.560 138.320 ;
    END
  END E2END[1]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.510500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.000 0.560 140.560 ;
    END
  END E2END[2]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.510500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 142.240 0.560 142.800 ;
    END
  END E2END[3]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.480 0.560 145.040 ;
    END
  END E2END[4]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.009000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 146.720 0.560 147.280 ;
    END
  END E2END[5]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.609500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 148.960 0.560 149.520 ;
    END
  END E2END[6]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 0.560 151.760 ;
    END
  END E2END[7]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 0.560 118.160 ;
    END
  END E2MID[0]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 119.840 0.560 120.400 ;
    END
  END E2MID[1]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 122.080 0.560 122.640 ;
    END
  END E2MID[2]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.705500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 0.560 124.880 ;
    END
  END E2MID[3]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.901000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.560 0.560 127.120 ;
    END
  END E2MID[4]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 128.800 0.560 129.360 ;
    END
  END E2MID[5]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.204000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.040 0.560 131.600 ;
    END
  END E2MID[6]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.102500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 133.280 0.560 133.840 ;
    END
  END E2MID[7]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 189.280 287.280 189.840 ;
    END
  END E6BEG[0]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 211.680 287.280 212.240 ;
    END
  END E6BEG[10]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 213.920 287.280 214.480 ;
    END
  END E6BEG[11]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 191.520 287.280 192.080 ;
    END
  END E6BEG[1]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 193.760 287.280 194.320 ;
    END
  END E6BEG[2]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 196.000 287.280 196.560 ;
    END
  END E6BEG[3]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 198.240 287.280 198.800 ;
    END
  END E6BEG[4]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 200.480 287.280 201.040 ;
    END
  END E6BEG[5]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 202.720 287.280 203.280 ;
    END
  END E6BEG[6]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 204.960 287.280 205.520 ;
    END
  END E6BEG[7]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 207.200 287.280 207.760 ;
    END
  END E6BEG[8]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 209.440 287.280 210.000 ;
    END
  END E6BEG[9]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.018000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 189.280 0.560 189.840 ;
    END
  END E6END[0]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.680 0.560 212.240 ;
    END
  END E6END[10]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 213.920 0.560 214.480 ;
    END
  END E6END[11]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.916000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 191.520 0.560 192.080 ;
    END
  END E6END[1]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 193.760 0.560 194.320 ;
    END
  END E6END[2]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 196.000 0.560 196.560 ;
    END
  END E6END[3]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.240 0.560 198.800 ;
    END
  END E6END[4]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 200.480 0.560 201.040 ;
    END
  END E6END[5]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 202.720 0.560 203.280 ;
    END
  END E6END[6]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.960 0.560 205.520 ;
    END
  END E6END[7]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.200 0.560 207.760 ;
    END
  END E6END[8]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 209.440 0.560 210.000 ;
    END
  END E6END[9]
  PIN EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 153.440 287.280 154.000 ;
    END
  END EE4BEG[0]
  PIN EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 175.840 287.280 176.400 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 178.080 287.280 178.640 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 180.320 287.280 180.880 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 182.560 287.280 183.120 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 184.800 287.280 185.360 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 187.040 287.280 187.600 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 155.680 287.280 156.240 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 157.920 287.280 158.480 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 160.160 287.280 160.720 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 162.400 287.280 162.960 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 164.640 287.280 165.200 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 166.880 287.280 167.440 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 169.120 287.280 169.680 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 171.360 287.280 171.920 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 173.600 287.280 174.160 ;
    END
  END EE4BEG[9]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 153.440 0.560 154.000 ;
    END
  END EE4END[0]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 175.840 0.560 176.400 ;
    END
  END EE4END[10]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 178.080 0.560 178.640 ;
    END
  END EE4END[11]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 180.320 0.560 180.880 ;
    END
  END EE4END[12]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.560 0.560 183.120 ;
    END
  END EE4END[13]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.800 0.560 185.360 ;
    END
  END EE4END[14]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 187.040 0.560 187.600 ;
    END
  END EE4END[15]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 155.680 0.560 156.240 ;
    END
  END EE4END[1]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.920 0.560 158.480 ;
    END
  END EE4END[2]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.105000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 160.160 0.560 160.720 ;
    END
  END EE4END[3]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 162.400 0.560 162.960 ;
    END
  END EE4END[4]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 0.560 165.200 ;
    END
  END EE4END[5]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.880 0.560 167.440 ;
    END
  END EE4END[6]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 169.120 0.560 169.680 ;
    END
  END EE4END[7]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 171.360 0.560 171.920 ;
    END
  END EE4END[8]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 173.600 0.560 174.160 ;
    END
  END EE4END[9]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 216.160 0.560 216.720 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 238.560 0.560 239.120 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 240.800 0.560 241.360 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 243.040 0.560 243.600 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 245.280 0.560 245.840 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 247.520 0.560 248.080 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 249.760 0.560 250.320 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 252.000 0.560 252.560 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.240 0.560 254.800 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 256.480 0.560 257.040 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 258.720 0.560 259.280 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 218.400 0.560 218.960 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 260.960 0.560 261.520 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 263.200 0.560 263.760 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 265.440 0.560 266.000 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 267.680 0.560 268.240 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 11.538500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 269.920 0.560 270.480 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 11.538500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 272.160 0.560 272.720 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 11.538500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 274.400 0.560 274.960 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 11.538500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 276.640 0.560 277.200 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 11.538500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.880 0.560 279.440 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 11.538500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 281.120 0.560 281.680 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 220.640 0.560 221.200 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 11.538500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 283.360 0.560 283.920 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 11.538500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.600 0.560 286.160 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 222.880 0.560 223.440 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 225.120 0.560 225.680 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 227.360 0.560 227.920 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 229.600 0.560 230.160 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 231.840 0.560 232.400 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 234.080 0.560 234.640 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.986500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 236.320 0.560 236.880 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 216.160 287.280 216.720 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 238.560 287.280 239.120 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 240.800 287.280 241.360 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 243.040 287.280 243.600 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 245.280 287.280 245.840 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 247.520 287.280 248.080 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 249.760 287.280 250.320 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 252.000 287.280 252.560 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 254.240 287.280 254.800 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 256.480 287.280 257.040 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 258.720 287.280 259.280 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 218.400 287.280 218.960 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 260.960 287.280 261.520 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 263.200 287.280 263.760 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 265.440 287.280 266.000 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 267.680 287.280 268.240 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 269.920 287.280 270.480 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 272.160 287.280 272.720 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 274.400 287.280 274.960 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 276.640 287.280 277.200 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 278.880 287.280 279.440 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 281.120 287.280 281.680 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 220.640 287.280 221.200 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 283.360 287.280 283.920 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 285.600 287.280 286.160 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 222.880 287.280 223.440 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 225.120 287.280 225.680 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 227.360 287.280 227.920 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 229.600 287.280 230.160 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 231.840 287.280 232.400 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 234.080 287.280 234.640 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 236.320 287.280 236.880 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 240.800 0.000 241.360 0.560 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 0.000 263.760 0.560 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 0.000 266.000 0.560 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 0.000 268.240 0.560 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 0.000 270.480 0.560 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 0.000 272.720 0.560 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 274.400 0.000 274.960 0.560 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 0.000 277.200 0.560 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 0.000 279.440 0.560 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 0.000 281.680 0.560 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.386500 ;
    PORT
      LAYER Metal2 ;
        RECT 283.360 0.000 283.920 0.560 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 243.040 0.000 243.600 0.560 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 0.000 245.840 0.560 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 0.000 248.080 0.560 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 0.000 250.320 0.560 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 0.000 252.560 0.560 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 254.240 0.000 254.800 0.560 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 0.000 257.040 0.560 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 0.000 259.280 0.560 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.050499 ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 0.000 261.520 0.560 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 240.800 286.720 241.360 287.280 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 286.720 263.760 287.280 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 286.720 266.000 287.280 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 286.720 268.240 287.280 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 286.720 270.480 287.280 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 286.720 272.720 287.280 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 274.400 286.720 274.960 287.280 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 286.720 277.200 287.280 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 286.720 279.440 287.280 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 286.720 281.680 287.280 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 283.360 286.720 283.920 287.280 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 243.040 286.720 243.600 287.280 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 286.720 245.840 287.280 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 286.720 248.080 287.280 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 286.720 250.320 287.280 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 286.720 252.560 287.280 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 254.240 286.720 254.800 287.280 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 286.720 257.040 287.280 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 286.720 259.280 287.280 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 286.720 261.520 287.280 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 286.720 3.920 287.280 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 5.600 286.720 6.160 287.280 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 7.840 286.720 8.400 287.280 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 286.720 10.640 287.280 ;
    END
  END N1BEG[3]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.015000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 0.560 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.015000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.600 0.000 6.160 0.560 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.015000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.840 0.000 8.400 0.560 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.015000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 0.000 10.640 0.560 ;
    END
  END N1END[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 12.320 286.720 12.880 287.280 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 14.560 286.720 15.120 287.280 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 286.720 17.360 287.280 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 19.040 286.720 19.600 287.280 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 21.280 286.720 21.840 287.280 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 286.720 24.080 287.280 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 286.720 26.320 287.280 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 286.720 28.560 287.280 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 286.720 30.800 287.280 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 286.720 33.040 287.280 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 286.720 35.280 287.280 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 286.720 37.520 287.280 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 286.720 39.760 287.280 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 286.720 42.000 287.280 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 286.720 44.240 287.280 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 286.720 46.480 287.280 ;
    END
  END N2BEGb[7]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.009000 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 0.560 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.108000 ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 0.000 33.040 0.560 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 0.000 35.280 0.560 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.009000 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 0.560 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.009000 ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 0.000 39.760 0.560 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 0.000 42.000 0.560 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 0.560 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.009000 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 0.000 46.480 0.560 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.003000 ;
    PORT
      LAYER Metal2 ;
        RECT 12.320 0.000 12.880 0.560 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.504500 ;
    PORT
      LAYER Metal2 ;
        RECT 14.560 0.000 15.120 0.560 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.003000 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 0.000 17.360 0.560 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.705500 ;
    PORT
      LAYER Metal2 ;
        RECT 19.040 0.000 19.600 0.560 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.952000 ;
    PORT
      LAYER Metal2 ;
        RECT 21.280 0.000 21.840 0.560 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.504500 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 0.560 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.603500 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 0.000 26.320 0.560 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.901000 ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 0.000 28.560 0.560 ;
    END
  END N2MID[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 286.720 48.720 287.280 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 286.720 71.120 287.280 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 286.720 73.360 287.280 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 286.720 75.600 287.280 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 286.720 77.840 287.280 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 286.720 80.080 287.280 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 286.720 82.320 287.280 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 286.720 50.960 287.280 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 286.720 53.200 287.280 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 286.720 55.440 287.280 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 286.720 57.680 287.280 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 286.720 59.920 287.280 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 286.720 62.160 287.280 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 286.720 64.400 287.280 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 286.720 66.640 287.280 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 286.720 68.880 287.280 ;
    END
  END N4BEG[9]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 0.000 48.720 0.560 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 0.560 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 0.000 73.360 0.560 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 0.000 75.600 0.560 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 0.560 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 0.000 80.080 0.560 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 0.000 82.320 0.560 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.456500 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 0.560 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 0.000 53.200 0.560 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 0.000 55.440 0.560 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 0.000 57.680 0.560 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 0.000 59.920 0.560 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 0.000 62.160 0.560 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 0.560 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 0.000 66.640 0.560 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 0.000 68.880 0.560 ;
    END
  END N4END[9]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 286.720 84.560 287.280 ;
    END
  END NN4BEG[0]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 286.720 106.960 287.280 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 286.720 109.200 287.280 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 286.720 111.440 287.280 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 286.720 113.680 287.280 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 286.720 115.920 287.280 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 286.720 118.160 287.280 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 286.720 86.800 287.280 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 286.720 89.040 287.280 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 286.720 91.280 287.280 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 286.720 93.520 287.280 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 286.720 95.760 287.280 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 286.720 98.000 287.280 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 286.720 100.240 287.280 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 286.720 102.480 287.280 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 286.720 104.720 287.280 ;
    END
  END NN4BEG[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 0.560 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 0.000 106.960 0.560 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 0.000 109.200 0.560 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 0.560 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 0.000 113.680 0.560 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 0.000 115.920 0.560 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 0.000 118.160 0.560 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 0.000 86.800 0.560 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 0.000 89.040 0.560 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.105000 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 0.560 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 0.000 93.520 0.560 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 0.000 95.760 0.560 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 0.560 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 0.000 100.240 0.560 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 0.000 102.480 0.560 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 0.560 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 0.000 122.640 0.560 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 0.560 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 0.000 127.120 0.560 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 0.000 129.360 0.560 ;
    END
  END S1BEG[3]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.012000 ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 286.720 122.640 287.280 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.012000 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 286.720 124.880 287.280 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.012000 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 286.720 127.120 287.280 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.012000 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 286.720 129.360 287.280 ;
    END
  END S1END[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 0.560 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 0.000 133.840 0.560 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 0.000 136.080 0.560 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 0.000 138.320 0.560 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 0.000 140.560 0.560 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 0.000 142.800 0.560 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 0.560 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 0.000 147.280 0.560 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 0.000 149.520 0.560 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 0.000 151.760 0.560 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 0.000 154.000 0.560 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 0.000 156.240 0.560 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 0.560 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 0.000 160.720 0.560 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 0.000 162.960 0.560 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 0.560 ;
    END
  END S2BEGb[7]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.009000 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 286.720 149.520 287.280 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405500 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 286.720 151.760 287.280 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.009000 ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 286.720 154.000 287.280 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 286.720 156.240 287.280 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 286.720 158.480 287.280 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 286.720 160.720 287.280 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.904000 ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 286.720 162.960 287.280 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.009000 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 286.720 165.200 287.280 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.003000 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 286.720 131.600 287.280 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.504500 ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 286.720 133.840 287.280 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.003000 ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 286.720 136.080 287.280 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.399500 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 286.720 138.320 287.280 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.003000 ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 286.720 140.560 287.280 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.504500 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 286.720 142.800 287.280 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 286.720 145.040 287.280 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.901000 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 286.720 147.280 287.280 ;
    END
  END S2MID[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 0.560 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 0.000 189.840 0.560 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 0.000 192.080 0.560 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 0.000 194.320 0.560 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 0.000 196.560 0.560 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 0.000 198.800 0.560 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 200.480 0.000 201.040 0.560 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 169.120 0.000 169.680 0.560 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 0.000 171.920 0.560 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 0.000 174.160 0.560 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 0.000 176.400 0.560 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 0.000 178.640 0.560 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 0.000 180.880 0.560 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 0.000 183.120 0.560 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 0.000 185.360 0.560 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 0.000 187.600 0.560 ;
    END
  END S4BEG[9]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 286.720 167.440 287.280 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 286.720 189.840 287.280 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 286.720 192.080 287.280 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 286.720 194.320 287.280 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 286.720 196.560 287.280 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 286.720 198.800 287.280 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 200.480 286.720 201.040 287.280 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 169.120 286.720 169.680 287.280 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 286.720 171.920 287.280 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 286.720 174.160 287.280 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 286.720 176.400 287.280 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 286.720 178.640 287.280 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 286.720 180.880 287.280 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 286.720 183.120 287.280 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 286.720 185.360 287.280 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 286.720 187.600 287.280 ;
    END
  END S4END[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 0.000 203.280 0.560 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 0.000 225.680 0.560 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 0.000 227.920 0.560 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 0.000 230.160 0.560 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 0.000 232.400 0.560 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 0.000 234.640 0.560 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 0.000 236.880 0.560 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 0.000 205.520 0.560 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 0.000 207.760 0.560 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 0.000 210.000 0.560 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 0.560 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 0.000 214.480 0.560 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 216.160 0.000 216.720 0.560 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 0.000 218.960 0.560 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 220.640 0.000 221.200 0.560 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 0.000 223.440 0.560 ;
    END
  END SS4BEG[9]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 286.720 203.280 287.280 ;
    END
  END SS4END[0]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 286.720 225.680 287.280 ;
    END
  END SS4END[10]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 286.720 227.920 287.280 ;
    END
  END SS4END[11]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 286.720 230.160 287.280 ;
    END
  END SS4END[12]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 286.720 232.400 287.280 ;
    END
  END SS4END[13]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 286.720 234.640 287.280 ;
    END
  END SS4END[14]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 286.720 236.880 287.280 ;
    END
  END SS4END[15]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 286.720 205.520 287.280 ;
    END
  END SS4END[1]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 286.720 207.760 287.280 ;
    END
  END SS4END[2]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 286.720 210.000 287.280 ;
    END
  END SS4END[3]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 286.720 212.240 287.280 ;
    END
  END SS4END[4]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 286.720 214.480 287.280 ;
    END
  END SS4END[5]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 216.160 286.720 216.720 287.280 ;
    END
  END SS4END[6]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 286.720 218.960 287.280 ;
    END
  END SS4END[7]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 220.640 286.720 221.200 287.280 ;
    END
  END SS4END[8]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 286.720 223.440 287.280 ;
    END
  END SS4END[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 0.000 239.120 0.560 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 286.720 239.120 287.280 ;
    END
  END UserCLKo
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.880 0.000 20.480 287.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 118.880 0.000 120.480 287.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.880 0.000 220.480 287.280 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.180 0.000 23.780 287.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.180 0.000 123.780 287.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 222.180 0.000 223.780 287.280 ;
    END
  END VSS
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1.120 0.560 1.680 ;
    END
  END W1BEG[0]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3.360 0.560 3.920 ;
    END
  END W1BEG[1]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 5.600 0.560 6.160 ;
    END
  END W1BEG[2]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 7.840 0.560 8.400 ;
    END
  END W1BEG[3]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.012000 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 1.120 287.280 1.680 ;
    END
  END W1END[0]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.513500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 3.360 287.280 3.920 ;
    END
  END W1END[1]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.516500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 5.600 287.280 6.160 ;
    END
  END W1END[2]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.516500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 7.840 287.280 8.400 ;
    END
  END W1END[3]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 10.080 0.560 10.640 ;
    END
  END W2BEG[0]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 12.320 0.560 12.880 ;
    END
  END W2BEG[1]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 14.560 0.560 15.120 ;
    END
  END W2BEG[2]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 16.800 0.560 17.360 ;
    END
  END W2BEG[3]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.040 0.560 19.600 ;
    END
  END W2BEG[4]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 21.280 0.560 21.840 ;
    END
  END W2BEG[5]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.520 0.560 24.080 ;
    END
  END W2BEG[6]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 25.760 0.560 26.320 ;
    END
  END W2BEG[7]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 28.000 0.560 28.560 ;
    END
  END W2BEGb[0]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.240 0.560 30.800 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 32.480 0.560 33.040 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 34.720 0.560 35.280 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 36.960 0.560 37.520 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.200 0.560 39.760 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 41.440 0.560 42.000 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.680 0.560 44.240 ;
    END
  END W2BEGb[7]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 28.000 287.280 28.560 ;
    END
  END W2END[0]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.564500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 30.240 287.280 30.800 ;
    END
  END W2END[1]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.009000 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 32.480 287.280 33.040 ;
    END
  END W2END[2]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.009000 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 34.720 287.280 35.280 ;
    END
  END W2END[3]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.510500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 36.960 287.280 37.520 ;
    END
  END W2END[4]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 39.200 287.280 39.760 ;
    END
  END W2END[5]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.558500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 41.440 287.280 42.000 ;
    END
  END W2END[6]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 43.680 287.280 44.240 ;
    END
  END W2END[7]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 10.080 287.280 10.640 ;
    END
  END W2MID[0]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 12.320 287.280 12.880 ;
    END
  END W2MID[1]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 14.560 287.280 15.120 ;
    END
  END W2MID[2]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.615500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 16.800 287.280 17.360 ;
    END
  END W2MID[3]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.105000 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 19.040 287.280 19.600 ;
    END
  END W2MID[4]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.504500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 21.280 287.280 21.840 ;
    END
  END W2MID[5]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.399500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 23.520 287.280 24.080 ;
    END
  END W2MID[6]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.060000 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 25.760 287.280 26.320 ;
    END
  END W2MID[7]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 81.760 0.560 82.320 ;
    END
  END W6BEG[0]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.160 0.560 104.720 ;
    END
  END W6BEG[10]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.400 0.560 106.960 ;
    END
  END W6BEG[11]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.000 0.560 84.560 ;
    END
  END W6BEG[1]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.240 0.560 86.800 ;
    END
  END W6BEG[2]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 88.480 0.560 89.040 ;
    END
  END W6BEG[3]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 0.560 91.280 ;
    END
  END W6BEG[4]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 92.960 0.560 93.520 ;
    END
  END W6BEG[5]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 95.200 0.560 95.760 ;
    END
  END W6BEG[6]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 97.440 0.560 98.000 ;
    END
  END W6BEG[7]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 99.680 0.560 100.240 ;
    END
  END W6BEG[8]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 101.920 0.560 102.480 ;
    END
  END W6BEG[9]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.012000 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 81.760 287.280 82.320 ;
    END
  END W6END[0]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 104.160 287.280 104.720 ;
    END
  END W6END[10]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 106.400 287.280 106.960 ;
    END
  END W6END[11]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.117000 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 84.000 287.280 84.560 ;
    END
  END W6END[1]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 86.240 287.280 86.800 ;
    END
  END W6END[2]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 88.480 287.280 89.040 ;
    END
  END W6END[3]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 90.720 287.280 91.280 ;
    END
  END W6END[4]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 92.960 287.280 93.520 ;
    END
  END W6END[5]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 95.200 287.280 95.760 ;
    END
  END W6END[6]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 97.440 287.280 98.000 ;
    END
  END W6END[7]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 99.680 287.280 100.240 ;
    END
  END W6END[8]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 101.920 287.280 102.480 ;
    END
  END W6END[9]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 45.920 0.560 46.480 ;
    END
  END WW4BEG[0]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 68.320 0.560 68.880 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.560 0.560 71.120 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 72.800 0.560 73.360 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 75.040 0.560 75.600 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 77.280 0.560 77.840 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 79.520 0.560 80.080 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.160 0.560 48.720 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.400 0.560 50.960 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 52.640 0.560 53.200 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 54.880 0.560 55.440 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 0.560 57.680 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.360 0.560 59.920 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.600 0.560 62.160 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 63.840 0.560 64.400 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.080 0.560 66.640 ;
    END
  END WW4BEG[9]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 45.920 287.280 46.480 ;
    END
  END WW4END[0]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 68.320 287.280 68.880 ;
    END
  END WW4END[10]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 70.560 287.280 71.120 ;
    END
  END WW4END[11]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 72.800 287.280 73.360 ;
    END
  END WW4END[12]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 75.040 287.280 75.600 ;
    END
  END WW4END[13]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 77.280 287.280 77.840 ;
    END
  END WW4END[14]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 79.520 287.280 80.080 ;
    END
  END WW4END[15]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 48.160 287.280 48.720 ;
    END
  END WW4END[1]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.006000 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 50.400 287.280 50.960 ;
    END
  END WW4END[2]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 52.640 287.280 53.200 ;
    END
  END WW4END[3]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 54.880 287.280 55.440 ;
    END
  END WW4END[4]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 57.120 287.280 57.680 ;
    END
  END WW4END[5]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 59.360 287.280 59.920 ;
    END
  END WW4END[6]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 61.600 287.280 62.160 ;
    END
  END WW4END[7]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 63.840 287.280 64.400 ;
    END
  END WW4END[8]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 66.080 287.280 66.640 ;
    END
  END WW4END[9]
  OBS
      LAYER Nwell ;
        RECT 2.930 3.490 284.350 282.670 ;
      LAYER Metal1 ;
        RECT 3.360 3.620 283.920 282.540 ;
      LAYER Metal2 ;
        RECT 0.140 286.420 3.060 286.720 ;
        RECT 4.220 286.420 5.300 286.720 ;
        RECT 6.460 286.420 7.540 286.720 ;
        RECT 8.700 286.420 9.780 286.720 ;
        RECT 10.940 286.420 12.020 286.720 ;
        RECT 13.180 286.420 14.260 286.720 ;
        RECT 15.420 286.420 16.500 286.720 ;
        RECT 17.660 286.420 18.740 286.720 ;
        RECT 19.900 286.420 20.980 286.720 ;
        RECT 22.140 286.420 23.220 286.720 ;
        RECT 24.380 286.420 25.460 286.720 ;
        RECT 26.620 286.420 27.700 286.720 ;
        RECT 28.860 286.420 29.940 286.720 ;
        RECT 31.100 286.420 32.180 286.720 ;
        RECT 33.340 286.420 34.420 286.720 ;
        RECT 35.580 286.420 36.660 286.720 ;
        RECT 37.820 286.420 38.900 286.720 ;
        RECT 40.060 286.420 41.140 286.720 ;
        RECT 42.300 286.420 43.380 286.720 ;
        RECT 44.540 286.420 45.620 286.720 ;
        RECT 46.780 286.420 47.860 286.720 ;
        RECT 49.020 286.420 50.100 286.720 ;
        RECT 51.260 286.420 52.340 286.720 ;
        RECT 53.500 286.420 54.580 286.720 ;
        RECT 55.740 286.420 56.820 286.720 ;
        RECT 57.980 286.420 59.060 286.720 ;
        RECT 60.220 286.420 61.300 286.720 ;
        RECT 62.460 286.420 63.540 286.720 ;
        RECT 64.700 286.420 65.780 286.720 ;
        RECT 66.940 286.420 68.020 286.720 ;
        RECT 69.180 286.420 70.260 286.720 ;
        RECT 71.420 286.420 72.500 286.720 ;
        RECT 73.660 286.420 74.740 286.720 ;
        RECT 75.900 286.420 76.980 286.720 ;
        RECT 78.140 286.420 79.220 286.720 ;
        RECT 80.380 286.420 81.460 286.720 ;
        RECT 82.620 286.420 83.700 286.720 ;
        RECT 84.860 286.420 85.940 286.720 ;
        RECT 87.100 286.420 88.180 286.720 ;
        RECT 89.340 286.420 90.420 286.720 ;
        RECT 91.580 286.420 92.660 286.720 ;
        RECT 93.820 286.420 94.900 286.720 ;
        RECT 96.060 286.420 97.140 286.720 ;
        RECT 98.300 286.420 99.380 286.720 ;
        RECT 100.540 286.420 101.620 286.720 ;
        RECT 102.780 286.420 103.860 286.720 ;
        RECT 105.020 286.420 106.100 286.720 ;
        RECT 107.260 286.420 108.340 286.720 ;
        RECT 109.500 286.420 110.580 286.720 ;
        RECT 111.740 286.420 112.820 286.720 ;
        RECT 113.980 286.420 115.060 286.720 ;
        RECT 116.220 286.420 117.300 286.720 ;
        RECT 118.460 286.420 119.540 286.720 ;
        RECT 120.700 286.420 121.780 286.720 ;
        RECT 122.940 286.420 124.020 286.720 ;
        RECT 125.180 286.420 126.260 286.720 ;
        RECT 127.420 286.420 128.500 286.720 ;
        RECT 129.660 286.420 130.740 286.720 ;
        RECT 131.900 286.420 132.980 286.720 ;
        RECT 134.140 286.420 135.220 286.720 ;
        RECT 136.380 286.420 137.460 286.720 ;
        RECT 138.620 286.420 139.700 286.720 ;
        RECT 140.860 286.420 141.940 286.720 ;
        RECT 143.100 286.420 144.180 286.720 ;
        RECT 145.340 286.420 146.420 286.720 ;
        RECT 147.580 286.420 148.660 286.720 ;
        RECT 149.820 286.420 150.900 286.720 ;
        RECT 152.060 286.420 153.140 286.720 ;
        RECT 154.300 286.420 155.380 286.720 ;
        RECT 156.540 286.420 157.620 286.720 ;
        RECT 158.780 286.420 159.860 286.720 ;
        RECT 161.020 286.420 162.100 286.720 ;
        RECT 163.260 286.420 164.340 286.720 ;
        RECT 165.500 286.420 166.580 286.720 ;
        RECT 167.740 286.420 168.820 286.720 ;
        RECT 169.980 286.420 171.060 286.720 ;
        RECT 172.220 286.420 173.300 286.720 ;
        RECT 174.460 286.420 175.540 286.720 ;
        RECT 176.700 286.420 177.780 286.720 ;
        RECT 178.940 286.420 180.020 286.720 ;
        RECT 181.180 286.420 182.260 286.720 ;
        RECT 183.420 286.420 184.500 286.720 ;
        RECT 185.660 286.420 186.740 286.720 ;
        RECT 187.900 286.420 188.980 286.720 ;
        RECT 190.140 286.420 191.220 286.720 ;
        RECT 192.380 286.420 193.460 286.720 ;
        RECT 194.620 286.420 195.700 286.720 ;
        RECT 196.860 286.420 197.940 286.720 ;
        RECT 199.100 286.420 200.180 286.720 ;
        RECT 201.340 286.420 202.420 286.720 ;
        RECT 203.580 286.420 204.660 286.720 ;
        RECT 205.820 286.420 206.900 286.720 ;
        RECT 208.060 286.420 209.140 286.720 ;
        RECT 210.300 286.420 211.380 286.720 ;
        RECT 212.540 286.420 213.620 286.720 ;
        RECT 214.780 286.420 215.860 286.720 ;
        RECT 217.020 286.420 218.100 286.720 ;
        RECT 219.260 286.420 220.340 286.720 ;
        RECT 221.500 286.420 222.580 286.720 ;
        RECT 223.740 286.420 224.820 286.720 ;
        RECT 225.980 286.420 227.060 286.720 ;
        RECT 228.220 286.420 229.300 286.720 ;
        RECT 230.460 286.420 231.540 286.720 ;
        RECT 232.700 286.420 233.780 286.720 ;
        RECT 234.940 286.420 236.020 286.720 ;
        RECT 237.180 286.420 238.260 286.720 ;
        RECT 239.420 286.420 240.500 286.720 ;
        RECT 241.660 286.420 242.740 286.720 ;
        RECT 243.900 286.420 244.980 286.720 ;
        RECT 246.140 286.420 247.220 286.720 ;
        RECT 248.380 286.420 249.460 286.720 ;
        RECT 250.620 286.420 251.700 286.720 ;
        RECT 252.860 286.420 253.940 286.720 ;
        RECT 255.100 286.420 256.180 286.720 ;
        RECT 257.340 286.420 258.420 286.720 ;
        RECT 259.580 286.420 260.660 286.720 ;
        RECT 261.820 286.420 262.900 286.720 ;
        RECT 264.060 286.420 265.140 286.720 ;
        RECT 266.300 286.420 267.380 286.720 ;
        RECT 268.540 286.420 269.620 286.720 ;
        RECT 270.780 286.420 271.860 286.720 ;
        RECT 273.020 286.420 274.100 286.720 ;
        RECT 275.260 286.420 276.340 286.720 ;
        RECT 277.500 286.420 278.580 286.720 ;
        RECT 279.740 286.420 280.820 286.720 ;
        RECT 281.980 286.420 283.060 286.720 ;
        RECT 284.220 286.420 287.140 286.720 ;
        RECT 0.140 0.860 287.140 286.420 ;
        RECT 0.140 0.090 3.060 0.860 ;
        RECT 4.220 0.090 5.300 0.860 ;
        RECT 6.460 0.090 7.540 0.860 ;
        RECT 8.700 0.090 9.780 0.860 ;
        RECT 10.940 0.090 12.020 0.860 ;
        RECT 13.180 0.090 14.260 0.860 ;
        RECT 15.420 0.090 16.500 0.860 ;
        RECT 17.660 0.090 18.740 0.860 ;
        RECT 19.900 0.090 20.980 0.860 ;
        RECT 22.140 0.090 23.220 0.860 ;
        RECT 24.380 0.090 25.460 0.860 ;
        RECT 26.620 0.090 27.700 0.860 ;
        RECT 28.860 0.090 29.940 0.860 ;
        RECT 31.100 0.090 32.180 0.860 ;
        RECT 33.340 0.090 34.420 0.860 ;
        RECT 35.580 0.090 36.660 0.860 ;
        RECT 37.820 0.090 38.900 0.860 ;
        RECT 40.060 0.090 41.140 0.860 ;
        RECT 42.300 0.090 43.380 0.860 ;
        RECT 44.540 0.090 45.620 0.860 ;
        RECT 46.780 0.090 47.860 0.860 ;
        RECT 49.020 0.090 50.100 0.860 ;
        RECT 51.260 0.090 52.340 0.860 ;
        RECT 53.500 0.090 54.580 0.860 ;
        RECT 55.740 0.090 56.820 0.860 ;
        RECT 57.980 0.090 59.060 0.860 ;
        RECT 60.220 0.090 61.300 0.860 ;
        RECT 62.460 0.090 63.540 0.860 ;
        RECT 64.700 0.090 65.780 0.860 ;
        RECT 66.940 0.090 68.020 0.860 ;
        RECT 69.180 0.090 70.260 0.860 ;
        RECT 71.420 0.090 72.500 0.860 ;
        RECT 73.660 0.090 74.740 0.860 ;
        RECT 75.900 0.090 76.980 0.860 ;
        RECT 78.140 0.090 79.220 0.860 ;
        RECT 80.380 0.090 81.460 0.860 ;
        RECT 82.620 0.090 83.700 0.860 ;
        RECT 84.860 0.090 85.940 0.860 ;
        RECT 87.100 0.090 88.180 0.860 ;
        RECT 89.340 0.090 90.420 0.860 ;
        RECT 91.580 0.090 92.660 0.860 ;
        RECT 93.820 0.090 94.900 0.860 ;
        RECT 96.060 0.090 97.140 0.860 ;
        RECT 98.300 0.090 99.380 0.860 ;
        RECT 100.540 0.090 101.620 0.860 ;
        RECT 102.780 0.090 103.860 0.860 ;
        RECT 105.020 0.090 106.100 0.860 ;
        RECT 107.260 0.090 108.340 0.860 ;
        RECT 109.500 0.090 110.580 0.860 ;
        RECT 111.740 0.090 112.820 0.860 ;
        RECT 113.980 0.090 115.060 0.860 ;
        RECT 116.220 0.090 117.300 0.860 ;
        RECT 118.460 0.090 119.540 0.860 ;
        RECT 120.700 0.090 121.780 0.860 ;
        RECT 122.940 0.090 124.020 0.860 ;
        RECT 125.180 0.090 126.260 0.860 ;
        RECT 127.420 0.090 128.500 0.860 ;
        RECT 129.660 0.090 130.740 0.860 ;
        RECT 131.900 0.090 132.980 0.860 ;
        RECT 134.140 0.090 135.220 0.860 ;
        RECT 136.380 0.090 137.460 0.860 ;
        RECT 138.620 0.090 139.700 0.860 ;
        RECT 140.860 0.090 141.940 0.860 ;
        RECT 143.100 0.090 144.180 0.860 ;
        RECT 145.340 0.090 146.420 0.860 ;
        RECT 147.580 0.090 148.660 0.860 ;
        RECT 149.820 0.090 150.900 0.860 ;
        RECT 152.060 0.090 153.140 0.860 ;
        RECT 154.300 0.090 155.380 0.860 ;
        RECT 156.540 0.090 157.620 0.860 ;
        RECT 158.780 0.090 159.860 0.860 ;
        RECT 161.020 0.090 162.100 0.860 ;
        RECT 163.260 0.090 164.340 0.860 ;
        RECT 165.500 0.090 166.580 0.860 ;
        RECT 167.740 0.090 168.820 0.860 ;
        RECT 169.980 0.090 171.060 0.860 ;
        RECT 172.220 0.090 173.300 0.860 ;
        RECT 174.460 0.090 175.540 0.860 ;
        RECT 176.700 0.090 177.780 0.860 ;
        RECT 178.940 0.090 180.020 0.860 ;
        RECT 181.180 0.090 182.260 0.860 ;
        RECT 183.420 0.090 184.500 0.860 ;
        RECT 185.660 0.090 186.740 0.860 ;
        RECT 187.900 0.090 188.980 0.860 ;
        RECT 190.140 0.090 191.220 0.860 ;
        RECT 192.380 0.090 193.460 0.860 ;
        RECT 194.620 0.090 195.700 0.860 ;
        RECT 196.860 0.090 197.940 0.860 ;
        RECT 199.100 0.090 200.180 0.860 ;
        RECT 201.340 0.090 202.420 0.860 ;
        RECT 203.580 0.090 204.660 0.860 ;
        RECT 205.820 0.090 206.900 0.860 ;
        RECT 208.060 0.090 209.140 0.860 ;
        RECT 210.300 0.090 211.380 0.860 ;
        RECT 212.540 0.090 213.620 0.860 ;
        RECT 214.780 0.090 215.860 0.860 ;
        RECT 217.020 0.090 218.100 0.860 ;
        RECT 219.260 0.090 220.340 0.860 ;
        RECT 221.500 0.090 222.580 0.860 ;
        RECT 223.740 0.090 224.820 0.860 ;
        RECT 225.980 0.090 227.060 0.860 ;
        RECT 228.220 0.090 229.300 0.860 ;
        RECT 230.460 0.090 231.540 0.860 ;
        RECT 232.700 0.090 233.780 0.860 ;
        RECT 234.940 0.090 236.020 0.860 ;
        RECT 237.180 0.090 238.260 0.860 ;
        RECT 239.420 0.090 240.500 0.860 ;
        RECT 241.660 0.090 242.740 0.860 ;
        RECT 243.900 0.090 244.980 0.860 ;
        RECT 246.140 0.090 247.220 0.860 ;
        RECT 248.380 0.090 249.460 0.860 ;
        RECT 250.620 0.090 251.700 0.860 ;
        RECT 252.860 0.090 253.940 0.860 ;
        RECT 255.100 0.090 256.180 0.860 ;
        RECT 257.340 0.090 258.420 0.860 ;
        RECT 259.580 0.090 260.660 0.860 ;
        RECT 261.820 0.090 262.900 0.860 ;
        RECT 264.060 0.090 265.140 0.860 ;
        RECT 266.300 0.090 267.380 0.860 ;
        RECT 268.540 0.090 269.620 0.860 ;
        RECT 270.780 0.090 271.860 0.860 ;
        RECT 273.020 0.090 274.100 0.860 ;
        RECT 275.260 0.090 276.340 0.860 ;
        RECT 277.500 0.090 278.580 0.860 ;
        RECT 279.740 0.090 280.820 0.860 ;
        RECT 281.980 0.090 283.060 0.860 ;
        RECT 284.220 0.090 287.140 0.860 ;
      LAYER Metal3 ;
        RECT 0.090 286.460 287.190 287.140 ;
        RECT 0.860 285.300 286.420 286.460 ;
        RECT 0.090 284.220 287.190 285.300 ;
        RECT 0.860 283.060 286.420 284.220 ;
        RECT 0.090 281.980 287.190 283.060 ;
        RECT 0.860 280.820 286.420 281.980 ;
        RECT 0.090 279.740 287.190 280.820 ;
        RECT 0.860 278.580 286.420 279.740 ;
        RECT 0.090 277.500 287.190 278.580 ;
        RECT 0.860 276.340 286.420 277.500 ;
        RECT 0.090 275.260 287.190 276.340 ;
        RECT 0.860 274.100 286.420 275.260 ;
        RECT 0.090 273.020 287.190 274.100 ;
        RECT 0.860 271.860 286.420 273.020 ;
        RECT 0.090 270.780 287.190 271.860 ;
        RECT 0.860 269.620 286.420 270.780 ;
        RECT 0.090 268.540 287.190 269.620 ;
        RECT 0.860 267.380 286.420 268.540 ;
        RECT 0.090 266.300 287.190 267.380 ;
        RECT 0.860 265.140 286.420 266.300 ;
        RECT 0.090 264.060 287.190 265.140 ;
        RECT 0.860 262.900 286.420 264.060 ;
        RECT 0.090 261.820 287.190 262.900 ;
        RECT 0.860 260.660 286.420 261.820 ;
        RECT 0.090 259.580 287.190 260.660 ;
        RECT 0.860 258.420 286.420 259.580 ;
        RECT 0.090 257.340 287.190 258.420 ;
        RECT 0.860 256.180 286.420 257.340 ;
        RECT 0.090 255.100 287.190 256.180 ;
        RECT 0.860 253.940 286.420 255.100 ;
        RECT 0.090 252.860 287.190 253.940 ;
        RECT 0.860 251.700 286.420 252.860 ;
        RECT 0.090 250.620 287.190 251.700 ;
        RECT 0.860 249.460 286.420 250.620 ;
        RECT 0.090 248.380 287.190 249.460 ;
        RECT 0.860 247.220 286.420 248.380 ;
        RECT 0.090 246.140 287.190 247.220 ;
        RECT 0.860 244.980 286.420 246.140 ;
        RECT 0.090 243.900 287.190 244.980 ;
        RECT 0.860 242.740 286.420 243.900 ;
        RECT 0.090 241.660 287.190 242.740 ;
        RECT 0.860 240.500 286.420 241.660 ;
        RECT 0.090 239.420 287.190 240.500 ;
        RECT 0.860 238.260 286.420 239.420 ;
        RECT 0.090 237.180 287.190 238.260 ;
        RECT 0.860 236.020 286.420 237.180 ;
        RECT 0.090 234.940 287.190 236.020 ;
        RECT 0.860 233.780 286.420 234.940 ;
        RECT 0.090 232.700 287.190 233.780 ;
        RECT 0.860 231.540 286.420 232.700 ;
        RECT 0.090 230.460 287.190 231.540 ;
        RECT 0.860 229.300 286.420 230.460 ;
        RECT 0.090 228.220 287.190 229.300 ;
        RECT 0.860 227.060 286.420 228.220 ;
        RECT 0.090 225.980 287.190 227.060 ;
        RECT 0.860 224.820 286.420 225.980 ;
        RECT 0.090 223.740 287.190 224.820 ;
        RECT 0.860 222.580 286.420 223.740 ;
        RECT 0.090 221.500 287.190 222.580 ;
        RECT 0.860 220.340 286.420 221.500 ;
        RECT 0.090 219.260 287.190 220.340 ;
        RECT 0.860 218.100 286.420 219.260 ;
        RECT 0.090 217.020 287.190 218.100 ;
        RECT 0.860 215.860 286.420 217.020 ;
        RECT 0.090 214.780 287.190 215.860 ;
        RECT 0.860 213.620 286.420 214.780 ;
        RECT 0.090 212.540 287.190 213.620 ;
        RECT 0.860 211.380 286.420 212.540 ;
        RECT 0.090 210.300 287.190 211.380 ;
        RECT 0.860 209.140 286.420 210.300 ;
        RECT 0.090 208.060 287.190 209.140 ;
        RECT 0.860 206.900 286.420 208.060 ;
        RECT 0.090 205.820 287.190 206.900 ;
        RECT 0.860 204.660 286.420 205.820 ;
        RECT 0.090 203.580 287.190 204.660 ;
        RECT 0.860 202.420 286.420 203.580 ;
        RECT 0.090 201.340 287.190 202.420 ;
        RECT 0.860 200.180 286.420 201.340 ;
        RECT 0.090 199.100 287.190 200.180 ;
        RECT 0.860 197.940 286.420 199.100 ;
        RECT 0.090 196.860 287.190 197.940 ;
        RECT 0.860 195.700 286.420 196.860 ;
        RECT 0.090 194.620 287.190 195.700 ;
        RECT 0.860 193.460 286.420 194.620 ;
        RECT 0.090 192.380 287.190 193.460 ;
        RECT 0.860 191.220 286.420 192.380 ;
        RECT 0.090 190.140 287.190 191.220 ;
        RECT 0.860 188.980 286.420 190.140 ;
        RECT 0.090 187.900 287.190 188.980 ;
        RECT 0.860 186.740 286.420 187.900 ;
        RECT 0.090 185.660 287.190 186.740 ;
        RECT 0.860 184.500 286.420 185.660 ;
        RECT 0.090 183.420 287.190 184.500 ;
        RECT 0.860 182.260 286.420 183.420 ;
        RECT 0.090 181.180 287.190 182.260 ;
        RECT 0.860 180.020 286.420 181.180 ;
        RECT 0.090 178.940 287.190 180.020 ;
        RECT 0.860 177.780 286.420 178.940 ;
        RECT 0.090 176.700 287.190 177.780 ;
        RECT 0.860 175.540 286.420 176.700 ;
        RECT 0.090 174.460 287.190 175.540 ;
        RECT 0.860 173.300 286.420 174.460 ;
        RECT 0.090 172.220 287.190 173.300 ;
        RECT 0.860 171.060 286.420 172.220 ;
        RECT 0.090 169.980 287.190 171.060 ;
        RECT 0.860 168.820 286.420 169.980 ;
        RECT 0.090 167.740 287.190 168.820 ;
        RECT 0.860 166.580 286.420 167.740 ;
        RECT 0.090 165.500 287.190 166.580 ;
        RECT 0.860 164.340 286.420 165.500 ;
        RECT 0.090 163.260 287.190 164.340 ;
        RECT 0.860 162.100 286.420 163.260 ;
        RECT 0.090 161.020 287.190 162.100 ;
        RECT 0.860 159.860 286.420 161.020 ;
        RECT 0.090 158.780 287.190 159.860 ;
        RECT 0.860 157.620 286.420 158.780 ;
        RECT 0.090 156.540 287.190 157.620 ;
        RECT 0.860 155.380 286.420 156.540 ;
        RECT 0.090 154.300 287.190 155.380 ;
        RECT 0.860 153.140 286.420 154.300 ;
        RECT 0.090 152.060 287.190 153.140 ;
        RECT 0.860 150.900 286.420 152.060 ;
        RECT 0.090 149.820 287.190 150.900 ;
        RECT 0.860 148.660 286.420 149.820 ;
        RECT 0.090 147.580 287.190 148.660 ;
        RECT 0.860 146.420 286.420 147.580 ;
        RECT 0.090 145.340 287.190 146.420 ;
        RECT 0.860 144.180 286.420 145.340 ;
        RECT 0.090 143.100 287.190 144.180 ;
        RECT 0.860 141.940 286.420 143.100 ;
        RECT 0.090 140.860 287.190 141.940 ;
        RECT 0.860 139.700 286.420 140.860 ;
        RECT 0.090 138.620 287.190 139.700 ;
        RECT 0.860 137.460 286.420 138.620 ;
        RECT 0.090 136.380 287.190 137.460 ;
        RECT 0.860 135.220 286.420 136.380 ;
        RECT 0.090 134.140 287.190 135.220 ;
        RECT 0.860 132.980 286.420 134.140 ;
        RECT 0.090 131.900 287.190 132.980 ;
        RECT 0.860 130.740 286.420 131.900 ;
        RECT 0.090 129.660 287.190 130.740 ;
        RECT 0.860 128.500 286.420 129.660 ;
        RECT 0.090 127.420 287.190 128.500 ;
        RECT 0.860 126.260 286.420 127.420 ;
        RECT 0.090 125.180 287.190 126.260 ;
        RECT 0.860 124.020 286.420 125.180 ;
        RECT 0.090 122.940 287.190 124.020 ;
        RECT 0.860 121.780 286.420 122.940 ;
        RECT 0.090 120.700 287.190 121.780 ;
        RECT 0.860 119.540 286.420 120.700 ;
        RECT 0.090 118.460 287.190 119.540 ;
        RECT 0.860 117.300 286.420 118.460 ;
        RECT 0.090 116.220 287.190 117.300 ;
        RECT 0.860 115.060 286.420 116.220 ;
        RECT 0.090 113.980 287.190 115.060 ;
        RECT 0.860 112.820 286.420 113.980 ;
        RECT 0.090 111.740 287.190 112.820 ;
        RECT 0.860 110.580 286.420 111.740 ;
        RECT 0.090 109.500 287.190 110.580 ;
        RECT 0.860 108.340 286.420 109.500 ;
        RECT 0.090 107.260 287.190 108.340 ;
        RECT 0.860 106.100 286.420 107.260 ;
        RECT 0.090 105.020 287.190 106.100 ;
        RECT 0.860 103.860 286.420 105.020 ;
        RECT 0.090 102.780 287.190 103.860 ;
        RECT 0.860 101.620 286.420 102.780 ;
        RECT 0.090 100.540 287.190 101.620 ;
        RECT 0.860 99.380 286.420 100.540 ;
        RECT 0.090 98.300 287.190 99.380 ;
        RECT 0.860 97.140 286.420 98.300 ;
        RECT 0.090 96.060 287.190 97.140 ;
        RECT 0.860 94.900 286.420 96.060 ;
        RECT 0.090 93.820 287.190 94.900 ;
        RECT 0.860 92.660 286.420 93.820 ;
        RECT 0.090 91.580 287.190 92.660 ;
        RECT 0.860 90.420 286.420 91.580 ;
        RECT 0.090 89.340 287.190 90.420 ;
        RECT 0.860 88.180 286.420 89.340 ;
        RECT 0.090 87.100 287.190 88.180 ;
        RECT 0.860 85.940 286.420 87.100 ;
        RECT 0.090 84.860 287.190 85.940 ;
        RECT 0.860 83.700 286.420 84.860 ;
        RECT 0.090 82.620 287.190 83.700 ;
        RECT 0.860 81.460 286.420 82.620 ;
        RECT 0.090 80.380 287.190 81.460 ;
        RECT 0.860 79.220 286.420 80.380 ;
        RECT 0.090 78.140 287.190 79.220 ;
        RECT 0.860 76.980 286.420 78.140 ;
        RECT 0.090 75.900 287.190 76.980 ;
        RECT 0.860 74.740 286.420 75.900 ;
        RECT 0.090 73.660 287.190 74.740 ;
        RECT 0.860 72.500 286.420 73.660 ;
        RECT 0.090 71.420 287.190 72.500 ;
        RECT 0.860 70.260 286.420 71.420 ;
        RECT 0.090 69.180 287.190 70.260 ;
        RECT 0.860 68.020 286.420 69.180 ;
        RECT 0.090 66.940 287.190 68.020 ;
        RECT 0.860 65.780 286.420 66.940 ;
        RECT 0.090 64.700 287.190 65.780 ;
        RECT 0.860 63.540 286.420 64.700 ;
        RECT 0.090 62.460 287.190 63.540 ;
        RECT 0.860 61.300 286.420 62.460 ;
        RECT 0.090 60.220 287.190 61.300 ;
        RECT 0.860 59.060 286.420 60.220 ;
        RECT 0.090 57.980 287.190 59.060 ;
        RECT 0.860 56.820 286.420 57.980 ;
        RECT 0.090 55.740 287.190 56.820 ;
        RECT 0.860 54.580 286.420 55.740 ;
        RECT 0.090 53.500 287.190 54.580 ;
        RECT 0.860 52.340 286.420 53.500 ;
        RECT 0.090 51.260 287.190 52.340 ;
        RECT 0.860 50.100 286.420 51.260 ;
        RECT 0.090 49.020 287.190 50.100 ;
        RECT 0.860 47.860 286.420 49.020 ;
        RECT 0.090 46.780 287.190 47.860 ;
        RECT 0.860 45.620 286.420 46.780 ;
        RECT 0.090 44.540 287.190 45.620 ;
        RECT 0.860 43.380 286.420 44.540 ;
        RECT 0.090 42.300 287.190 43.380 ;
        RECT 0.860 41.140 286.420 42.300 ;
        RECT 0.090 40.060 287.190 41.140 ;
        RECT 0.860 38.900 286.420 40.060 ;
        RECT 0.090 37.820 287.190 38.900 ;
        RECT 0.860 36.660 286.420 37.820 ;
        RECT 0.090 35.580 287.190 36.660 ;
        RECT 0.860 34.420 286.420 35.580 ;
        RECT 0.090 33.340 287.190 34.420 ;
        RECT 0.860 32.180 286.420 33.340 ;
        RECT 0.090 31.100 287.190 32.180 ;
        RECT 0.860 29.940 286.420 31.100 ;
        RECT 0.090 28.860 287.190 29.940 ;
        RECT 0.860 27.700 286.420 28.860 ;
        RECT 0.090 26.620 287.190 27.700 ;
        RECT 0.860 25.460 286.420 26.620 ;
        RECT 0.090 24.380 287.190 25.460 ;
        RECT 0.860 23.220 286.420 24.380 ;
        RECT 0.090 22.140 287.190 23.220 ;
        RECT 0.860 20.980 286.420 22.140 ;
        RECT 0.090 19.900 287.190 20.980 ;
        RECT 0.860 18.740 286.420 19.900 ;
        RECT 0.090 17.660 287.190 18.740 ;
        RECT 0.860 16.500 286.420 17.660 ;
        RECT 0.090 15.420 287.190 16.500 ;
        RECT 0.860 14.260 286.420 15.420 ;
        RECT 0.090 13.180 287.190 14.260 ;
        RECT 0.860 12.020 286.420 13.180 ;
        RECT 0.090 10.940 287.190 12.020 ;
        RECT 0.860 9.780 286.420 10.940 ;
        RECT 0.090 8.700 287.190 9.780 ;
        RECT 0.860 7.540 286.420 8.700 ;
        RECT 0.090 6.460 287.190 7.540 ;
        RECT 0.860 5.300 286.420 6.460 ;
        RECT 0.090 4.220 287.190 5.300 ;
        RECT 0.860 3.060 286.420 4.220 ;
        RECT 0.090 1.980 287.190 3.060 ;
        RECT 0.860 0.820 286.420 1.980 ;
        RECT 0.090 0.140 287.190 0.820 ;
      LAYER Metal4 ;
        RECT 0.700 0.090 18.580 287.190 ;
        RECT 20.780 0.090 21.880 287.190 ;
        RECT 24.080 0.090 118.580 287.190 ;
        RECT 120.780 0.090 121.880 287.190 ;
        RECT 124.080 0.090 218.580 287.190 ;
        RECT 220.780 0.090 221.880 287.190 ;
        RECT 224.080 0.090 287.140 287.190 ;
  END
END LUT4AB
END LIBRARY

