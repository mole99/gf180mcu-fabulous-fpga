module LUT4AB (Ci,
    Co,
    UserCLK,
    UserCLKo,
    E1BEG,
    E1END,
    E2BEG,
    E2BEGb,
    E2END,
    E2MID,
    E6BEG,
    E6END,
    EE4BEG,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    NN4BEG,
    NN4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    SS4BEG,
    SS4END,
    W1BEG,
    W1END,
    W2BEG,
    W2BEGb,
    W2END,
    W2MID,
    W6BEG,
    W6END,
    WW4BEG,
    WW4END);
 input Ci;
 output Co;
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 input [3:0] E1END;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 input [7:0] E2END;
 input [7:0] E2MID;
 output [11:0] E6BEG;
 input [11:0] E6END;
 output [15:0] EE4BEG;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [15:0] NN4BEG;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [15:0] SS4BEG;
 input [15:0] SS4END;
 output [3:0] W1BEG;
 input [3:0] W1END;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 input [7:0] W2END;
 input [7:0] W2MID;
 output [11:0] W6BEG;
 input [11:0] W6END;
 output [15:0] WW4BEG;
 input [15:0] WW4END;

 wire A;
 wire B;
 wire C;
 wire net1;
 wire D;
 wire E;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire F;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire G;
 wire H;
 wire \Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.E6BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E6BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.M_AB ;
 wire \Inst_LUT4AB_switch_matrix.M_AD ;
 wire \Inst_LUT4AB_switch_matrix.M_AH ;
 wire \Inst_LUT4AB_switch_matrix.M_EF ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.W6BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.W6BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG3 ;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire UserCLK_regs;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_0_UserCLK_regs;
 wire clknet_1_0__leaf_UserCLK_regs;
 wire clknet_1_1__leaf_UserCLK_regs;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0859_ (.I(S2MID[6]),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0860_ (.I(W2MID[6]),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0861_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0862_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0863_ (.I(N2MID[7]),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0864_ (.I(S2MID[7]),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0865_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0866_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0867_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0868_ (.I(S2MID[3]),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0869_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0870_ (.I(E2MID[4]),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0871_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0872_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0873_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0874_ (.I(E6END[1]),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0875_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0876_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0877_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0878_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0879_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0880_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0881_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0882_ (.I(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0883_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0884_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0885_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0886_ (.I(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0887_ (.I(\Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0888_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0889_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0890_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0891_ (.I(S2END[6]),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0892_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0893_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0894_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0895_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0896_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0897_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0898_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0899_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0900_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0901_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0902_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0903_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0904_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0905_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0906_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0907_ (.I(\Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0908_ (.I(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0909_ (.I(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0910_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0911_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0912_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0913_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0914_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0915_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0916_ (.I(S2END[1]),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0917_ (.I(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0918_ (.I(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0919_ (.I(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0920_ (.I(\Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0921_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0922_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0923_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0924_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0925_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0926_ (.I(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0927_ (.I(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0928_ (.I(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0929_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0930_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0931_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0932_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0933_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0934_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0935_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0936_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0937_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0938_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0939_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0940_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ),
    .A2(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0941_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0942_ (.A1(_0715_),
    .A2(_0789_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0943_ (.I0(N1END[2]),
    .I1(N2END[4]),
    .I2(N4END[0]),
    .I3(E2END[4]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0944_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ),
    .A2(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0945_ (.I0(E6END[0]),
    .I1(S2END[4]),
    .I2(W2END[4]),
    .I3(W6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0946_ (.A1(_0715_),
    .A2(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0947_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ),
    .A2(_0792_),
    .A3(_0794_),
    .B1(_0788_),
    .B2(_0790_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0948_ (.I0(E2MID[2]),
    .I1(S2MID[2]),
    .I2(W2MID[2]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0949_ (.I0(N2MID[3]),
    .I1(E2MID[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0950_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ),
    .A2(W2MID[3]),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0951_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ),
    .A2(_0716_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ),
    .C(_0797_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0952_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ),
    .A2(_0796_),
    .B(_0798_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0953_ (.I(_0799_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0954_ (.I0(A),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0955_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .A2(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0956_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0957_ (.A1(_0717_),
    .A2(_0803_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0958_ (.I0(N1END[0]),
    .I1(N2END[2]),
    .I2(N4END[2]),
    .I3(E2END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0959_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .A2(_0805_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0960_ (.I0(E6END[0]),
    .I1(S2END[2]),
    .I2(W2END[2]),
    .I3(WW4END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0961_ (.A1(_0717_),
    .A2(_0807_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0962_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ),
    .A2(_0806_),
    .A3(_0808_),
    .B1(_0802_),
    .B2(_0804_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0963_ (.I0(EE4END[2]),
    .I1(S4END[2]),
    .I2(W2END[7]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0964_ (.I0(NN4END[0]),
    .I1(S2END[2]),
    .I2(E2END[2]),
    .I3(W2END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0965_ (.I0(_0795_),
    .I1(_0800_),
    .I2(_0810_),
    .I3(_0809_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0966_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0967_ (.A1(_0709_),
    .A2(_0812_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0968_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0969_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .A2(_0814_),
    .B(_0710_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0970_ (.I0(E6END[0]),
    .I1(S2END[4]),
    .I2(W2END[4]),
    .I3(W6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0971_ (.I0(N2END[4]),
    .I1(E1END[2]),
    .I2(N4END[0]),
    .I3(E2END[4]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0972_ (.A1(_0709_),
    .A2(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0973_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .A2(_0816_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0974_ (.A1(_0813_),
    .A2(_0815_),
    .B1(_0818_),
    .B2(_0819_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0975_ (.I0(N2MID[6]),
    .I1(S2MID[6]),
    .I2(W2MID[6]),
    .I3(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0976_ (.I0(N2MID[7]),
    .I1(E2MID[7]),
    .I2(S2MID[7]),
    .I3(W2MID[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0977_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0978_ (.I0(A),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0979_ (.A1(_0713_),
    .A2(_0823_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0980_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .A2(_0822_),
    .B(_0714_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0981_ (.I0(E6END[0]),
    .I1(S2END[2]),
    .I2(W2END[2]),
    .I3(W6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0982_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .A2(_0826_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0983_ (.I0(N2END[2]),
    .I1(E1END[0]),
    .I2(N4END[2]),
    .I3(E2END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0984_ (.A1(_0713_),
    .A2(_0828_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0985_ (.A1(_0824_),
    .A2(_0825_),
    .B1(_0827_),
    .B2(_0829_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0986_ (.I0(NN4END[3]),
    .I1(WW4END[0]),
    .I2(S4END[3]),
    .I3(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0987_ (.I0(N2END[6]),
    .I1(SS4END[3]),
    .I2(E2END[6]),
    .I3(W2END[6]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0988_ (.I(_0831_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0989_ (.I0(_0820_),
    .I1(_0821_),
    .I2(_0831_),
    .I3(_0830_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0990_ (.I0(_0833_),
    .I1(Ci),
    .S(\Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0991_ (.I0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .I1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .S(_0834_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0992_ (.A1(N4END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0993_ (.A1(_0722_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ),
    .C(_0836_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0994_ (.I0(A),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0995_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0996_ (.A1(_0723_),
    .A2(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0997_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ),
    .A2(_0838_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0998_ (.I0(NN4END[2]),
    .I1(EE4END[2]),
    .I2(E1END[0]),
    .I3(E6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0999_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ),
    .A2(_0842_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1000_ (.I0(S4END[2]),
    .I1(SS4END[2]),
    .I2(W2END[2]),
    .I3(W6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1001_ (.A1(_0723_),
    .A2(_0844_),
    .B(_0724_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1002_ (.A1(_0840_),
    .A2(_0841_),
    .B1(_0843_),
    .B2(_0845_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1003_ (.A1(_0840_),
    .A2(_0841_),
    .B1(_0843_),
    .B2(_0845_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1004_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .A2(W6END[1]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1005_ (.I(_0847_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1006_ (.I0(N4END[1]),
    .I1(E6END[1]),
    .I2(W6END[1]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1007_ (.A1(_0846_),
    .A2(_0848_),
    .B(_0721_),
    .C(_0837_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1008_ (.I0(N2END[4]),
    .I1(S2END[4]),
    .I2(EE4END[0]),
    .I3(W2END[4]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1009_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ),
    .A2(_0851_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1010_ (.A1(_0725_),
    .A2(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1011_ (.I(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1012_ (.A1(_0850_),
    .A2(_0854_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1013_ (.A1(N2MID[4]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1014_ (.A1(_0718_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ),
    .C(_0856_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1015_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1016_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1017_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .A2(_0008_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1018_ (.A1(_0719_),
    .A2(_0858_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1019_ (.I0(S2END[4]),
    .I1(W2END[4]),
    .I2(S4END[0]),
    .I3(WW4END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1020_ (.A1(_0719_),
    .A2(_0011_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1021_ (.I0(N2END[4]),
    .I1(E1END[2]),
    .I2(E2END[4]),
    .I3(E6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1022_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .A2(_0013_),
    .B(_0720_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1023_ (.A1(_0009_),
    .A2(_0010_),
    .B1(_0012_),
    .B2(_0014_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1024_ (.A1(_0009_),
    .A2(_0010_),
    .B1(_0012_),
    .B2(_0014_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1025_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .A2(W2MID[4]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1026_ (.I(_0016_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1027_ (.I0(N2MID[4]),
    .I1(E2MID[4]),
    .I2(W2MID[4]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1028_ (.A1(_0015_),
    .A2(_0017_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ),
    .C(_0857_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1029_ (.I0(N2MID[5]),
    .I1(E2MID[5]),
    .I2(S2MID[5]),
    .I3(W2MID[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1030_ (.A1(_0721_),
    .A2(_0020_),
    .B(_0725_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1031_ (.A1(_0019_),
    .A2(_0021_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1032_ (.A1(_0855_),
    .A2(_0022_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1033_ (.A1(_0850_),
    .A2(_0854_),
    .B1(_0019_),
    .B2(_0021_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1034_ (.I0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .I1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .S(_0834_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1035_ (.I0(_0835_),
    .I1(_0025_),
    .S(_0811_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1036_ (.I0(A),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1037_ (.A1(_0728_),
    .A2(_0027_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1038_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1039_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .A2(_0029_),
    .B(_0729_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1040_ (.I0(N1END[0]),
    .I1(E2END[2]),
    .I2(N2END[2]),
    .I3(E6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1041_ (.I0(S2END[2]),
    .I1(W2END[2]),
    .I2(S4END[2]),
    .I3(W6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1042_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .A2(_0032_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1043_ (.A1(_0728_),
    .A2(_0031_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1044_ (.A1(_0028_),
    .A2(_0030_),
    .B1(_0033_),
    .B2(_0034_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1045_ (.I0(N4END[0]),
    .I1(E6END[0]),
    .I2(S4END[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1046_ (.I0(N2END[0]),
    .I1(S2END[0]),
    .I2(E2END[0]),
    .I3(WW4END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1047_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1048_ (.A1(_0726_),
    .A2(_0037_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1049_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1050_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .A2(_0039_),
    .B(_0727_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1051_ (.I0(N1END[2]),
    .I1(E2END[4]),
    .I2(N2END[4]),
    .I3(E6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1052_ (.I0(S2END[4]),
    .I1(W2END[4]),
    .I2(S4END[0]),
    .I3(WW4END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1053_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .A2(_0042_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1054_ (.A1(_0726_),
    .A2(_0041_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1055_ (.A1(_0038_),
    .A2(_0040_),
    .B1(_0043_),
    .B2(_0044_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1056_ (.I0(N2MID[0]),
    .I1(E2MID[0]),
    .I2(S2MID[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1057_ (.I0(N2MID[1]),
    .I1(E2MID[1]),
    .I2(S2MID[1]),
    .I3(W2MID[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1058_ (.I(_0046_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1059_ (.I0(_0045_),
    .I1(_0046_),
    .I2(_0036_),
    .I3(_0035_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1060_ (.I0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .I1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .S(_0834_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1061_ (.I0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .I1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .S(_0834_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1062_ (.I0(_0049_),
    .I1(_0050_),
    .S(_0811_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1063_ (.I0(_0026_),
    .I1(_0051_),
    .S(_0023_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1064_ (.A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A2(_0834_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1065_ (.I0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .I1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S(_0834_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1066_ (.A1(_0730_),
    .A2(_0834_),
    .B(_0811_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1067_ (.A1(_0811_),
    .A2(_0054_),
    .B1(_0055_),
    .B2(_0053_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1068_ (.A1(_0023_),
    .A2(_0056_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1069_ (.I0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .I1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .S(_0834_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1070_ (.I0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .I1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .S(_0834_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1071_ (.I0(_0059_),
    .I1(_0058_),
    .S(_0811_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1072_ (.A1(_0023_),
    .A2(_0060_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1073_ (.A1(_0048_),
    .A2(_0061_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1074_ (.A1(_0048_),
    .A2(_0052_),
    .B1(_0057_),
    .B2(_0062_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1075_ (.A1(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .A2(\Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1076_ (.A1(\Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ),
    .A2(_0063_),
    .B(_0064_),
    .ZN(A));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1077_ (.A1(_0736_),
    .A2(_0045_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1078_ (.A1(_0736_),
    .A2(_0047_),
    .B(_0065_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1079_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ),
    .A2(_0035_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1080_ (.A1(_0736_),
    .A2(_0036_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1081_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ),
    .A2(_0067_),
    .A3(_0068_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1082_ (.A1(_0066_),
    .A2(_0069_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1083_ (.A1(_0066_),
    .A2(_0069_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1084_ (.I0(_0018_),
    .I1(_0020_),
    .I2(_0851_),
    .I3(_0849_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1085_ (.I(_0072_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1086_ (.I0(_0795_),
    .I1(_0800_),
    .I2(_0810_),
    .I3(_0809_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1087_ (.I(_0074_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1088_ (.A1(_0073_),
    .A2(_0074_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1089_ (.A1(_0072_),
    .A2(_0075_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1090_ (.A1(_0072_),
    .A2(_0074_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1091_ (.A1(_0073_),
    .A2(_0075_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1092_ (.A1(_0072_),
    .A2(_0074_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1093_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A2(_0077_),
    .B1(_0079_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1094_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(_0076_),
    .B1(_0080_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .C(_0071_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1095_ (.I0(_0820_),
    .I1(_0821_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1096_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ),
    .A2(_0832_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1097_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ),
    .A2(_0830_),
    .B(_0084_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1098_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ),
    .A2(_0083_),
    .B(_0735_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1099_ (.A1(_0811_),
    .A2(_0024_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1100_ (.A1(_0811_),
    .A2(_0024_),
    .B(Ci),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1101_ (.A1(_0735_),
    .A2(_0087_),
    .A3(_0088_),
    .B1(_0085_),
    .B2(_0086_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _1102_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(_0076_),
    .B1(_0077_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .C1(_0080_),
    .C2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1103_ (.I(_0090_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1104_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A2(_0079_),
    .B(_0091_),
    .C(_0070_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1105_ (.A1(_0081_),
    .A2(_0082_),
    .B(_0092_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1106_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(_0076_),
    .B1(_0077_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1107_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A2(_0079_),
    .B1(_0080_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .C(_0071_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _1108_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(_0076_),
    .B1(_0077_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .C1(_0079_),
    .C2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1109_ (.I(_0096_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1110_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A2(_0080_),
    .B(_0097_),
    .C(_0070_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1111_ (.A1(_0094_),
    .A2(_0095_),
    .B(_0098_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1112_ (.I0(_0093_),
    .I1(_0099_),
    .S(_0089_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1113_ (.I0(_0100_),
    .I1(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ),
    .Z(B));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1114_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1115_ (.A1(_0742_),
    .A2(_0101_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1116_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1117_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .A2(_0103_),
    .B(_0743_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1118_ (.I0(S1END[1]),
    .I1(S2END[5]),
    .I2(S1END[3]),
    .I3(W1END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1119_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .A2(_0105_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1120_ (.I0(N1END[1]),
    .I1(N2END[5]),
    .I2(E1END[1]),
    .I3(E2END[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1121_ (.A1(_0742_),
    .A2(_0107_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1122_ (.A1(_0102_),
    .A2(_0104_),
    .B1(_0106_),
    .B2(_0108_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1123_ (.I0(N2MID[2]),
    .I1(W2MID[2]),
    .I2(E2MID[2]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1124_ (.I0(N2MID[3]),
    .I1(E2MID[3]),
    .I2(S2MID[3]),
    .I3(W2MID[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1125_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1126_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .A2(_0111_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1127_ (.I0(A),
    .I1(B),
    .I2(D),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1128_ (.A1(_0744_),
    .A2(_0113_),
    .B(_0745_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1129_ (.I0(N1END[1]),
    .I1(N4END[3]),
    .I2(N2END[3]),
    .I3(E2END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1130_ (.I0(E6END[1]),
    .I1(S2END[3]),
    .I2(W2END[3]),
    .I3(W6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1131_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .A2(_0116_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1132_ (.A1(_0744_),
    .A2(_0115_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1133_ (.A1(_0112_),
    .A2(_0114_),
    .B1(_0117_),
    .B2(_0118_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1134_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1135_ (.I0(N4END[2]),
    .I1(E2END[2]),
    .I2(W2END[7]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1136_ (.I0(N2END[2]),
    .I1(E2END[2]),
    .I2(S2END[2]),
    .I3(WW4END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1137_ (.I0(_0109_),
    .I1(_0110_),
    .I2(_0121_),
    .I3(_0120_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1138_ (.I(_0122_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1139_ (.I0(A),
    .I1(B),
    .I2(D),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1140_ (.A1(_0748_),
    .A2(_0124_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1141_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1142_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .A2(_0126_),
    .B(_0749_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1143_ (.I0(NN4END[3]),
    .I1(E1END[1]),
    .I2(E2END[3]),
    .I3(E6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1144_ (.A1(_0748_),
    .A2(_0128_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1145_ (.I0(S2END[3]),
    .I1(W2END[3]),
    .I2(S4END[3]),
    .I3(W6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1146_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .A2(_0130_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1147_ (.A1(_0125_),
    .A2(_0127_),
    .B1(_0129_),
    .B2(_0131_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1148_ (.I0(NN4END[1]),
    .I1(EE4END[1]),
    .I2(S4END[1]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1149_ (.I0(N2END[4]),
    .I1(E2END[4]),
    .I2(SS4END[2]),
    .I3(W2END[4]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1150_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1151_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1152_ (.A1(_0746_),
    .A2(_0135_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1153_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .A2(_0134_),
    .B(_0747_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1154_ (.I0(N1END[1]),
    .I1(N2END[5]),
    .I2(E1END[1]),
    .I3(E2END[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1155_ (.I0(S1END[1]),
    .I1(S2END[5]),
    .I2(W1END[1]),
    .I3(W1END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1156_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .A2(_0139_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1157_ (.A1(_0746_),
    .A2(_0138_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1158_ (.A1(_0136_),
    .A2(_0137_),
    .B1(_0140_),
    .B2(_0141_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1159_ (.I0(N2MID[4]),
    .I1(E2MID[4]),
    .I2(S2MID[4]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1160_ (.I0(N2MID[5]),
    .I1(E2MID[5]),
    .I2(S2MID[5]),
    .I3(W2MID[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1161_ (.I0(_0142_),
    .I1(_0143_),
    .I2(_0133_),
    .I3(_0132_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1162_ (.A1(_0122_),
    .A2(_0144_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1163_ (.A1(_0122_),
    .A2(_0144_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1164_ (.A1(_0122_),
    .A2(_0144_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1165_ (.I0(_0109_),
    .I1(_0110_),
    .I2(_0121_),
    .I3(_0120_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1166_ (.I(_0148_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1167_ (.I0(_0142_),
    .I1(_0143_),
    .I2(_0133_),
    .I3(_0132_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1168_ (.A1(_0148_),
    .A2(_0150_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1169_ (.A1(_0148_),
    .A2(_0150_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1170_ (.I(_0152_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1171_ (.A1(_0078_),
    .A2(_0087_),
    .A3(_0088_),
    .B(_0080_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1172_ (.A1(_0151_),
    .A2(_0154_),
    .B(_0152_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1173_ (.A1(_0122_),
    .A2(_0144_),
    .B1(_0151_),
    .B2(_0154_),
    .C(_0152_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1174_ (.I0(N4END[3]),
    .I1(W2END[3]),
    .I2(E2END[3]),
    .I3(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1175_ (.I0(N2END[7]),
    .I1(S2END[7]),
    .I2(EE4END[2]),
    .I3(W2END[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1176_ (.I0(E),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1177_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .A2(_0159_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1178_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1179_ (.A1(_0753_),
    .A2(_0161_),
    .B(_0754_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1180_ (.I0(N1END[2]),
    .I1(N2END[6]),
    .I2(E1END[2]),
    .I3(E2END[6]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1181_ (.I0(S1END[2]),
    .I1(W1END[0]),
    .I2(S2END[6]),
    .I3(W1END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1182_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .A2(_0164_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1183_ (.A1(_0753_),
    .A2(_0163_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1184_ (.A1(_0160_),
    .A2(_0162_),
    .B1(_0165_),
    .B2(_0166_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1185_ (.I0(N2MID[6]),
    .I1(W2MID[6]),
    .I2(E2MID[6]),
    .I3(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1186_ (.A1(W2MID[7]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1187_ (.A1(_0712_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ),
    .C(_0168_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1188_ (.A1(E2MID[7]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1189_ (.A1(_0711_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ),
    .B(_0170_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1190_ (.A1(_0169_),
    .A2(_0171_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1191_ (.A1(_0169_),
    .A2(_0171_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1192_ (.I0(_0167_),
    .I1(_0173_),
    .I2(_0158_),
    .I3(_0157_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1193_ (.A1(_0755_),
    .A2(_0174_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1194_ (.A1(_0755_),
    .A2(_0145_),
    .A3(_0156_),
    .B(_0175_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1195_ (.I0(NN4END[2]),
    .I1(S4END[2]),
    .I2(E2END[2]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1196_ (.I0(N2END[3]),
    .I1(S2END[3]),
    .I2(E2END[3]),
    .I3(WW4END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1197_ (.I0(E),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1198_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1199_ (.A1(_0758_),
    .A2(_0180_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1200_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .A2(_0179_),
    .B(_0759_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1201_ (.I0(S1END[0]),
    .I1(S1END[2]),
    .I2(S2END[6]),
    .I3(W1END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1202_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .A2(_0183_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1203_ (.I0(N1END[2]),
    .I1(N2END[6]),
    .I2(E1END[2]),
    .I3(E2END[6]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1204_ (.A1(_0758_),
    .A2(_0185_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1205_ (.A1(_0181_),
    .A2(_0182_),
    .B1(_0184_),
    .B2(_0186_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1206_ (.I0(N2MID[2]),
    .I1(S2MID[2]),
    .I2(E2MID[2]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1207_ (.A1(W2MID[3]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1208_ (.A1(_0716_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ),
    .C(_0188_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1209_ (.I0(N2MID[3]),
    .I1(E2MID[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1210_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ),
    .A2(_0190_),
    .B(_0189_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1211_ (.I(_0191_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1212_ (.I0(_0187_),
    .I1(_0192_),
    .I2(_0178_),
    .I3(_0177_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1213_ (.I0(N4END[1]),
    .I1(SS4END[1]),
    .I2(W2END[4]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1214_ (.I0(N2END[5]),
    .I1(E2END[5]),
    .I2(SS4END[1]),
    .I3(W2END[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1215_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1216_ (.A1(_0760_),
    .A2(_0196_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1217_ (.I0(E),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1218_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .A2(_0198_),
    .B(_0761_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1219_ (.I0(N1END[2]),
    .I1(N2END[6]),
    .I2(E1END[2]),
    .I3(E2END[6]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1220_ (.I0(S1END[2]),
    .I1(W1END[0]),
    .I2(S2END[6]),
    .I3(W1END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1221_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .A2(_0201_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1222_ (.A1(_0760_),
    .A2(_0200_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1223_ (.A1(_0197_),
    .A2(_0199_),
    .B1(_0202_),
    .B2(_0203_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1224_ (.I0(N2MID[4]),
    .I1(W2MID[4]),
    .I2(S2MID[4]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1225_ (.I0(N2MID[5]),
    .I1(E2MID[5]),
    .I2(S2MID[5]),
    .I3(W2MID[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1226_ (.I0(_0204_),
    .I1(_0205_),
    .I2(_0195_),
    .I3(_0194_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1227_ (.I(_0206_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1228_ (.A1(_0193_),
    .A2(_0206_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1229_ (.A1(_0193_),
    .A2(_0207_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1230_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A2(_0193_),
    .A3(_0207_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1231_ (.A1(_0193_),
    .A2(_0206_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1232_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(_0209_),
    .B1(_0211_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1233_ (.A1(_0756_),
    .A2(_0208_),
    .B(_0210_),
    .C(_0212_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1234_ (.I0(EE4END[3]),
    .I1(WW4END[1]),
    .I2(S4END[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1235_ (.I0(NN4END[2]),
    .I1(E2END[1]),
    .I2(S2END[1]),
    .I3(W2END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1236_ (.I(_0215_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1237_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1238_ (.I0(E),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1239_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .A2(_0218_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1240_ (.A1(_0762_),
    .A2(_0217_),
    .B(_0763_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1241_ (.I0(N1END[2]),
    .I1(N2END[6]),
    .I2(E1END[2]),
    .I3(E2END[6]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1242_ (.I0(S1END[0]),
    .I1(S1END[2]),
    .I2(S2END[6]),
    .I3(W1END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1243_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .A2(_0222_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1244_ (.A1(_0762_),
    .A2(_0221_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1245_ (.A1(_0219_),
    .A2(_0220_),
    .B1(_0223_),
    .B2(_0224_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1246_ (.I0(E2MID[0]),
    .I1(S2MID[0]),
    .I2(W2MID[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1247_ (.I0(N2MID[1]),
    .I1(E2MID[1]),
    .I2(S2MID[1]),
    .I3(W2MID[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1248_ (.I(_0226_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1249_ (.I0(_0225_),
    .I1(_0226_),
    .I2(_0215_),
    .I3(_0214_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1250_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A2(_0193_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1251_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(_0209_),
    .B1(_0211_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1252_ (.A1(_0757_),
    .A2(_0208_),
    .B1(_0229_),
    .B2(_0206_),
    .C(_0230_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1253_ (.I0(_0231_),
    .I1(_0213_),
    .S(_0176_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1254_ (.I0(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .I1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .I2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .I3(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S0(_0193_),
    .S1(_0206_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1255_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A2(_0193_),
    .A3(_0207_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1256_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(_0209_),
    .B1(_0211_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .C(_0234_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1257_ (.A1(_0765_),
    .A2(_0208_),
    .B(_0235_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1258_ (.I0(_0236_),
    .I1(_0233_),
    .S(_0176_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1259_ (.I0(_0232_),
    .I1(_0237_),
    .S(_0228_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1260_ (.I0(_0238_),
    .I1(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ),
    .Z(E));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1261_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1262_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1263_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .A2(_0240_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1264_ (.A1(_0737_),
    .A2(_0239_),
    .B(_0738_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1265_ (.I0(S1END[1]),
    .I1(S2END[5]),
    .I2(W1END[1]),
    .I3(W1END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1266_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .A2(_0243_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1267_ (.I0(N1END[1]),
    .I1(N2END[5]),
    .I2(E1END[1]),
    .I3(E2END[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1268_ (.A1(_0737_),
    .A2(_0245_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1269_ (.A1(_0241_),
    .A2(_0242_),
    .B1(_0244_),
    .B2(_0246_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1270_ (.I0(E2MID[6]),
    .I1(S2MID[6]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1271_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1272_ (.A1(_0708_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ),
    .C(_0248_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1273_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ),
    .A2(_0247_),
    .B(_0249_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1274_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .A2(_0250_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1275_ (.I0(N2MID[7]),
    .I1(E2MID[7]),
    .I2(S2MID[7]),
    .I3(W2MID[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1276_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .A2(_0252_),
    .B(_0251_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1277_ (.I0(A),
    .I1(B),
    .I2(D),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1278_ (.A1(_0740_),
    .A2(_0254_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1279_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1280_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ),
    .A2(_0256_),
    .B(_0741_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1281_ (.I0(N2END[3]),
    .I1(N4END[3]),
    .I2(E1END[1]),
    .I3(E2END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1282_ (.I0(E6END[1]),
    .I1(S2END[3]),
    .I2(W2END[3]),
    .I3(WW4END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1283_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ),
    .A2(_0259_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1284_ (.A1(_0740_),
    .A2(_0258_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1285_ (.A1(_0255_),
    .A2(_0257_),
    .B1(_0260_),
    .B2(_0261_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1286_ (.I0(E2END[3]),
    .I1(WW4END[2]),
    .I2(SS4END[3]),
    .I3(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1287_ (.A1(W2END[6]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1288_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ),
    .A2(_0739_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ),
    .C(_0263_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1289_ (.I0(NN4END[3]),
    .I1(E2END[6]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1290_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ),
    .A2(_0265_),
    .B(_0264_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1291_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .A2(_0266_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1292_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .A2(_0262_),
    .B(_0267_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1293_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ),
    .A2(_0253_),
    .A3(_0268_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1294_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ),
    .A2(_0154_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1295_ (.A1(_0269_),
    .A2(_0270_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1296_ (.A1(_0149_),
    .A2(_0150_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1297_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A2(_0151_),
    .B1(_0272_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1298_ (.A1(_0149_),
    .A2(_0150_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1299_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(_0153_),
    .B1(_0274_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1300_ (.A1(_0273_),
    .A2(_0275_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1301_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A2(_0151_),
    .B1(_0274_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1302_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(_0153_),
    .B1(_0272_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1303_ (.A1(_0277_),
    .A2(_0278_),
    .B(_0271_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1304_ (.I0(A),
    .I1(B),
    .I2(D),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1305_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1306_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .A2(_0281_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1307_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ),
    .A2(_0282_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1308_ (.A1(_0752_),
    .A2(_0280_),
    .B(_0283_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1309_ (.I0(N1END[1]),
    .I1(N2END[3]),
    .I2(EE4END[3]),
    .I3(E6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1310_ (.I0(S4END[3]),
    .I1(W2END[3]),
    .I2(SS4END[3]),
    .I3(W6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1311_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .A2(_0286_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1312_ (.A1(_0752_),
    .A2(_0285_),
    .B(_0287_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1313_ (.A1(_0284_),
    .A2(_0288_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1314_ (.I0(N4END[0]),
    .I1(W6END[0]),
    .I2(SS4END[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1315_ (.I0(N2END[0]),
    .I1(S2END[0]),
    .I2(EE4END[1]),
    .I3(W2END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1316_ (.I(_0290_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1317_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1318_ (.A1(_0750_),
    .A2(_0292_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1319_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1320_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .A2(_0294_),
    .B(_0751_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1321_ (.I0(N1END[1]),
    .I1(N2END[5]),
    .I2(E1END[1]),
    .I3(E2END[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1322_ (.I0(S1END[1]),
    .I1(S2END[5]),
    .I2(S1END[3]),
    .I3(W1END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1323_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .A2(_0297_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1324_ (.A1(_0750_),
    .A2(_0296_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1325_ (.A1(_0293_),
    .A2(_0295_),
    .B1(_0298_),
    .B2(_0299_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1326_ (.I0(N2MID[0]),
    .I1(S2MID[0]),
    .I2(W2MID[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1327_ (.I0(N2MID[1]),
    .I1(E2MID[1]),
    .I2(S2MID[1]),
    .I3(W2MID[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1328_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ),
    .A2(_0289_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1329_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ),
    .A2(_0291_),
    .B(_0302_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1330_ (.I0(_0300_),
    .I1(_0301_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1331_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ),
    .A2(_0304_),
    .B(_0303_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1332_ (.I(_0305_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1333_ (.A1(_0271_),
    .A2(_0276_),
    .B(_0279_),
    .C(_0306_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1334_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0151_),
    .B1(_0274_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1335_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A2(_0153_),
    .B1(_0272_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1336_ (.A1(_0308_),
    .A2(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1337_ (.A1(_0271_),
    .A2(_0310_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1338_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A2(_0153_),
    .B1(_0274_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1339_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A2(_0151_),
    .B1(_0272_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1340_ (.A1(_0312_),
    .A2(_0313_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1341_ (.A1(_0269_),
    .A2(_0270_),
    .A3(_0314_),
    .B(_0305_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1342_ (.A1(_0311_),
    .A2(_0315_),
    .B(_0307_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1343_ (.I0(_0316_),
    .I1(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ),
    .Z(C));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1344_ (.A1(_0145_),
    .A2(_0156_),
    .A3(_0208_),
    .B(_0211_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1345_ (.I0(_0167_),
    .I1(_0173_),
    .I2(_0158_),
    .I3(_0157_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1346_ (.I0(_0318_),
    .I1(_0317_),
    .S(\Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1347_ (.I0(_0204_),
    .I1(_0205_),
    .I2(_0195_),
    .I3(_0194_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1348_ (.I(_0320_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1349_ (.I0(_0187_),
    .I1(_0192_),
    .I2(_0178_),
    .I3(_0177_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1350_ (.A1(_0320_),
    .A2(_0322_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1351_ (.A1(_0320_),
    .A2(_0322_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1352_ (.I(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1353_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A2(_0323_),
    .B1(_0324_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1354_ (.A1(_0321_),
    .A2(_0322_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1355_ (.A1(_0321_),
    .A2(_0322_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1356_ (.I(_0328_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1357_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(_0327_),
    .B1(_0329_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1358_ (.A1(_0326_),
    .A2(_0330_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1359_ (.A1(_0319_),
    .A2(_0331_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1360_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0214_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1361_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0216_),
    .B(_0333_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1362_ (.I0(_0225_),
    .I1(_0226_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1363_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ),
    .A2(_0335_),
    .B(_0334_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1364_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0323_),
    .B1(_0324_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1365_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(_0327_),
    .B1(_0329_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1366_ (.A1(_0337_),
    .A2(_0338_),
    .B(_0319_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1367_ (.A1(_0332_),
    .A2(_0336_),
    .A3(_0339_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1368_ (.A1(_0767_),
    .A2(_0319_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1369_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(_0319_),
    .B(_0324_),
    .C(_0341_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1370_ (.I0(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .I1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .S(_0319_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1371_ (.A1(_0766_),
    .A2(_0319_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1372_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(_0319_),
    .B(_0327_),
    .C(_0344_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1373_ (.I0(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .I1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .S(_0319_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1374_ (.A1(_0329_),
    .A2(_0343_),
    .B1(_0346_),
    .B2(_0323_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1375_ (.A1(_0336_),
    .A2(_0342_),
    .A3(_0345_),
    .A4(_0347_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1376_ (.A1(_0340_),
    .A2(_0348_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1377_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1378_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ),
    .A2(_0349_),
    .B(_0350_),
    .ZN(F));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1379_ (.A1(_0317_),
    .A2(_0323_),
    .B(_0325_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1380_ (.I0(E),
    .I1(H),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1381_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .A2(_0352_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1382_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1383_ (.A1(_0731_),
    .A2(_0354_),
    .B(_0732_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1384_ (.I0(N1END[3]),
    .I1(N2END[7]),
    .I2(E1END[3]),
    .I3(E2END[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1385_ (.I0(S1END[3]),
    .I1(W1END[1]),
    .I2(S2END[7]),
    .I3(W1END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1386_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .A2(_0357_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1387_ (.A1(_0731_),
    .A2(_0356_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1388_ (.A1(_0353_),
    .A2(_0355_),
    .B1(_0358_),
    .B2(_0359_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1389_ (.I0(N2MID[6]),
    .I1(E2MID[6]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1390_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1391_ (.A1(_0707_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ),
    .C(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1392_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ),
    .A2(_0360_),
    .B(_0362_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1393_ (.I0(N2MID[7]),
    .I1(E2MID[7]),
    .I2(S2MID[7]),
    .I3(W2MID[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1394_ (.I0(N4END[3]),
    .I1(EE4END[0]),
    .I2(S4END[3]),
    .I3(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1395_ (.I0(N2END[7]),
    .I1(E2END[7]),
    .I2(S2END[7]),
    .I3(WW4END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1396_ (.I(_0366_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1397_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_0364_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1398_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_0363_),
    .B(_0368_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1399_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_0365_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1400_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_0367_),
    .B(_0370_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1401_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ),
    .A2(_0369_),
    .B(_0371_),
    .C(_0768_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1402_ (.A1(_0768_),
    .A2(_0351_),
    .B(_0372_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1403_ (.I0(N4END[2]),
    .I1(W2END[2]),
    .I2(SS4END[2]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1404_ (.I0(N2END[3]),
    .I1(SS4END[0]),
    .I2(E2END[3]),
    .I3(W2END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1405_ (.I0(E),
    .I1(H),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1406_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1407_ (.A1(_0769_),
    .A2(_0377_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1408_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .A2(_0376_),
    .B(_0770_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1409_ (.I0(S1END[1]),
    .I1(S1END[3]),
    .I2(S2END[7]),
    .I3(W1END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1410_ (.I0(N1END[3]),
    .I1(N2END[7]),
    .I2(E1END[3]),
    .I3(E2END[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1411_ (.A1(_0769_),
    .A2(_0381_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1412_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .A2(_0380_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1413_ (.A1(_0378_),
    .A2(_0379_),
    .B1(_0382_),
    .B2(_0383_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1414_ (.I0(N2MID[2]),
    .I1(W2MID[2]),
    .I2(S2MID[2]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1415_ (.I0(N2MID[3]),
    .I1(E2MID[3]),
    .I2(S2MID[3]),
    .I3(W2MID[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1416_ (.I0(_0384_),
    .I1(_0385_),
    .I2(_0375_),
    .I3(_0374_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1417_ (.I(_0386_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1418_ (.I0(E6END[1]),
    .I1(S4END[1]),
    .I2(WW4END[3]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1419_ (.I0(NN4END[1]),
    .I1(S2END[5]),
    .I2(E2END[5]),
    .I3(W2END[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1420_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1421_ (.A1(_0771_),
    .A2(_0390_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1422_ (.I0(E),
    .I1(H),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1423_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .A2(_0392_),
    .B(_0772_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1424_ (.I0(N1END[3]),
    .I1(N2END[7]),
    .I2(E1END[3]),
    .I3(E2END[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1425_ (.I0(S1END[3]),
    .I1(W1END[1]),
    .I2(S2END[7]),
    .I3(W1END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1426_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .A2(_0395_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1427_ (.A1(_0771_),
    .A2(_0394_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1428_ (.A1(_0391_),
    .A2(_0393_),
    .B1(_0396_),
    .B2(_0397_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1429_ (.I0(E2MID[4]),
    .I1(W2MID[4]),
    .I2(S2MID[4]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1430_ (.I0(N2MID[5]),
    .I1(E2MID[5]),
    .I2(S2MID[5]),
    .I3(W2MID[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1431_ (.I0(_0398_),
    .I1(_0399_),
    .I2(_0389_),
    .I3(_0388_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1432_ (.A1(_0386_),
    .A2(_0400_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1433_ (.A1(_0387_),
    .A2(_0400_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1434_ (.A1(_0386_),
    .A2(_0400_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1435_ (.I0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .I1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .I2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .I3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S0(_0386_),
    .S1(_0400_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1436_ (.I0(NN4END[0]),
    .I1(W2END[0]),
    .I2(E6END[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1437_ (.I0(N2END[1]),
    .I1(EE4END[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1438_ (.A1(W2END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1439_ (.A1(_0764_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ),
    .C(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1440_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ),
    .A2(_0406_),
    .B(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1441_ (.I(_0409_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1442_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1443_ (.A1(_0773_),
    .A2(_0411_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1444_ (.I0(E),
    .I1(H),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1445_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .A2(_0413_),
    .B(_0412_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1446_ (.I0(S1END[1]),
    .I1(S1END[3]),
    .I2(S2END[7]),
    .I3(W1END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1447_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .A2(_0415_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1448_ (.I0(N1END[3]),
    .I1(N2END[7]),
    .I2(E1END[3]),
    .I3(E2END[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1449_ (.A1(_0773_),
    .A2(_0417_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1450_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ),
    .A2(_0414_),
    .B1(_0416_),
    .B2(_0418_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1451_ (.I0(N2MID[0]),
    .I1(E2MID[0]),
    .I2(W2MID[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1452_ (.I0(N2MID[1]),
    .I1(E2MID[1]),
    .I2(S2MID[1]),
    .I3(W2MID[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1453_ (.I0(_0419_),
    .I1(_0420_),
    .I2(_0410_),
    .I3(_0405_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1454_ (.A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(_0387_),
    .A3(_0400_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1455_ (.A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A2(_0402_),
    .B1(_0403_),
    .B2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1456_ (.A1(_0774_),
    .A2(_0401_),
    .B(_0422_),
    .C(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1457_ (.I0(_0424_),
    .I1(_0404_),
    .S(_0373_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1458_ (.I0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .I1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .I2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .I3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .S0(_0386_),
    .S1(_0400_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1459_ (.I0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .I1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .I2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .I3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .S0(_0386_),
    .S1(_0400_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1460_ (.I0(_0427_),
    .I1(_0426_),
    .S(_0373_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1461_ (.I0(_0428_),
    .I1(_0425_),
    .S(_0421_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1462_ (.I0(_0429_),
    .I1(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ),
    .Z(G));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1463_ (.A1(_0317_),
    .A2(_0323_),
    .B1(_0386_),
    .B2(_0400_),
    .C(_0325_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1464_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0364_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1465_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0363_),
    .B(_0431_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1466_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0365_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1467_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0367_),
    .B(_0433_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1468_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ),
    .A2(_0432_),
    .B(_0434_),
    .C(_0775_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1469_ (.A1(_0775_),
    .A2(_0401_),
    .A3(_0430_),
    .B(_0435_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1470_ (.I0(_0398_),
    .I1(_0399_),
    .I2(_0389_),
    .I3(_0388_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1471_ (.I(_0437_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1472_ (.I0(_0384_),
    .I1(_0385_),
    .I2(_0375_),
    .I3(_0374_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1473_ (.I(_0439_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1474_ (.A1(_0437_),
    .A2(_0440_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1475_ (.A1(_0438_),
    .A2(_0439_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1476_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A2(_0441_),
    .B1(_0442_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1477_ (.A1(_0438_),
    .A2(_0440_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1478_ (.A1(_0437_),
    .A2(_0439_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1479_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A2(_0444_),
    .B1(_0445_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1480_ (.A1(_0443_),
    .A2(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1481_ (.I0(_0419_),
    .I1(_0420_),
    .I2(_0410_),
    .I3(_0405_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1482_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A2(_0441_),
    .B1(_0444_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1483_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(_0442_),
    .B1(_0445_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1484_ (.A1(_0449_),
    .A2(_0450_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1485_ (.I0(_0451_),
    .I1(_0447_),
    .S(_0436_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1486_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A2(_0441_),
    .B1(_0445_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1487_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(_0442_),
    .B1(_0444_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1488_ (.A1(_0453_),
    .A2(_0454_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1489_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A2(_0441_),
    .B1(_0444_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1490_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(_0442_),
    .B1(_0445_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1491_ (.A1(_0456_),
    .A2(_0457_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1492_ (.I0(_0458_),
    .I1(_0455_),
    .S(_0436_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1493_ (.I0(_0459_),
    .I1(_0452_),
    .S(_0448_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1494_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ),
    .A2(_0460_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1495_ (.A1(_0776_),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ),
    .B(_0461_),
    .ZN(H));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1496_ (.I0(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .I1(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1497_ (.I0(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .I1(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1498_ (.I0(_0462_),
    .I1(_0463_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1499_ (.I0(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .I1(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .I2(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1500_ (.I0(_0464_),
    .I1(_0465_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1501_ (.I0(E),
    .I1(F),
    .S(_0466_),
    .Z(\Inst_LUT4AB_switch_matrix.M_EF ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1502_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .A2(_0252_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1503_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .A2(_0250_),
    .B(_0467_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1504_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .A2(_0262_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1505_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .A2(_0266_),
    .B(_0469_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1506_ (.A1(_0468_),
    .A2(_0470_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1507_ (.I0(_0471_),
    .I1(_0155_),
    .S(\Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1508_ (.A1(_0123_),
    .A2(_0144_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1509_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A2(_0146_),
    .B1(_0473_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1510_ (.A1(_0123_),
    .A2(_0144_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1511_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(_0147_),
    .B1(_0475_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1512_ (.A1(_0474_),
    .A2(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1513_ (.A1(_0472_),
    .A2(_0477_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1514_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A2(_0146_),
    .B1(_0475_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1515_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(_0147_),
    .B1(_0473_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1516_ (.A1(_0479_),
    .A2(_0480_),
    .B(_0472_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1517_ (.I(_0481_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1518_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ),
    .A2(_0289_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1519_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ),
    .A2(_0291_),
    .B(_0483_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1520_ (.I0(_0300_),
    .I1(_0301_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1521_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ),
    .A2(_0485_),
    .B(_0484_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1522_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A2(_0146_),
    .B1(_0147_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1523_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A2(_0473_),
    .B1(_0475_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1524_ (.A1(_0487_),
    .A2(_0488_),
    .B(_0472_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1525_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0146_),
    .B1(_0147_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1526_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A2(_0473_),
    .B1(_0475_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1527_ (.A1(_0490_),
    .A2(_0491_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1528_ (.A1(_0472_),
    .A2(_0492_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1529_ (.A1(_0486_),
    .A2(_0489_),
    .A3(_0493_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1530_ (.A1(_0478_),
    .A2(_0482_),
    .A3(_0486_),
    .B(_0494_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1531_ (.I0(_0495_),
    .I1(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ),
    .Z(D));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1532_ (.I0(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .I1(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .I2(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1533_ (.I0(_0465_),
    .I1(_0496_),
    .S(_0783_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1534_ (.I0(C),
    .I1(D),
    .S(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1535_ (.I0(\Inst_LUT4AB_switch_matrix.M_AB ),
    .I1(_0498_),
    .S(_0496_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1536_ (.I0(_0498_),
    .I1(_0499_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.M_AD ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1537_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1538_ (.I0(E),
    .I1(G),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1539_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .A2(_0501_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1540_ (.A1(_0781_),
    .A2(_0500_),
    .B(_0782_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1541_ (.I0(N1END[0]),
    .I1(N2END[0]),
    .I2(E1END[0]),
    .I3(E2END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1542_ (.I0(S1END[0]),
    .I1(W1END[0]),
    .I2(S2END[0]),
    .I3(W1END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1543_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .A2(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1544_ (.A1(_0781_),
    .A2(_0504_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1545_ (.A1(_0502_),
    .A2(_0503_),
    .B1(_0506_),
    .B2(_0507_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1546_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1547_ (.I(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1548_ (.I0(E),
    .I1(G),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1549_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .A2(_0510_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1550_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .A2(_0509_),
    .B(_0511_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1551_ (.I0(N1END[0]),
    .I1(NN4END[0]),
    .I2(E1END[0]),
    .I3(E2END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1552_ (.I0(S1END[0]),
    .I1(S1END[2]),
    .I2(S2END[0]),
    .I3(W1END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1553_ (.I0(_0513_),
    .I1(_0514_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1554_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ),
    .A2(_0515_),
    .B(_0512_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1555_ (.I(_0516_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1556_ (.I0(E),
    .I1(G),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1557_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1558_ (.A1(_0777_),
    .A2(_0518_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1559_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .A2(_0517_),
    .B(_0778_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1560_ (.I0(N1END[0]),
    .I1(N2END[0]),
    .I2(E1END[0]),
    .I3(EE4END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1561_ (.A1(_0777_),
    .A2(_0521_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1562_ (.I0(S1END[0]),
    .I1(W1END[0]),
    .I2(S2END[0]),
    .I3(W1END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1563_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .A2(_0523_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1564_ (.A1(_0519_),
    .A2(_0520_),
    .B1(_0522_),
    .B2(_0524_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1565_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1566_ (.I0(E),
    .I1(G),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1567_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1568_ (.A1(_0779_),
    .A2(_0525_),
    .B(_0780_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1569_ (.I0(S1END[0]),
    .I1(S1END[2]),
    .I2(SS4END[0]),
    .I3(WW4END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1570_ (.I0(N1END[0]),
    .I1(N2END[0]),
    .I2(E1END[0]),
    .I3(E2END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1571_ (.A1(_0779_),
    .A2(_0530_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1572_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(_0529_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1573_ (.A1(_0527_),
    .A2(_0528_),
    .B1(_0531_),
    .B2(_0532_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1574_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1575_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1576_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .B(_0534_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1577_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(_0516_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1578_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .B(_0536_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1579_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ),
    .A2(_0535_),
    .B(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1580_ (.I0(_0538_),
    .I1(_0496_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1581_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .A2(_0466_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1582_ (.A1(_0783_),
    .A2(_0539_),
    .B(_0540_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1583_ (.I0(H),
    .I1(G),
    .S(_0541_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1584_ (.I0(\Inst_LUT4AB_switch_matrix.M_EF ),
    .I1(_0542_),
    .S(_0539_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1585_ (.I0(_0499_),
    .I1(_0543_),
    .S(_0538_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1586_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .A2(_0544_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1587_ (.A1(_0783_),
    .A2(_0543_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1588_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .A2(_0542_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1589_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .A2(_0546_),
    .A3(_0547_),
    .B(_0545_),
    .ZN(\Inst_LUT4AB_switch_matrix.M_AH ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1590_ (.I0(A),
    .I1(B),
    .S(_0465_),
    .Z(\Inst_LUT4AB_switch_matrix.M_AB ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1591_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1592_ (.A1(_0784_),
    .A2(_0548_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1593_ (.I0(B),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1594_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .A2(_0550_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1595_ (.I0(S2END[1]),
    .I1(W2END[1]),
    .I2(S4END[1]),
    .I3(W6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1596_ (.A1(_0784_),
    .A2(_0552_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1597_ (.I0(N1END[3]),
    .I1(E2END[1]),
    .I2(N2END[1]),
    .I3(E6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1598_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .A2(_0554_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1599_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0553_),
    .A3(_0555_),
    .B1(_0549_),
    .B2(_0551_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1600_ (.I0(B),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1601_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1602_ (.I(_0557_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1603_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0558_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1604_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0556_),
    .B(_0559_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1605_ (.I0(NN4END[1]),
    .I1(E2END[1]),
    .I2(E1END[3]),
    .I3(E6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1606_ (.I0(S2END[1]),
    .I1(W2END[1]),
    .I2(S4END[1]),
    .I3(W6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1607_ (.I(_0562_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1608_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0563_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1609_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0561_),
    .B(_0564_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1610_ (.A1(_0560_),
    .A2(_0565_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1611_ (.I0(B),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1612_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .A2(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1613_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1614_ (.A1(_0785_),
    .A2(_0568_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1615_ (.I0(N1END[3]),
    .I1(N2END[1]),
    .I2(N4END[1]),
    .I3(EE4END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1616_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .A2(_0570_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1617_ (.I0(E6END[1]),
    .I1(W2END[1]),
    .I2(S2END[1]),
    .I3(W6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1618_ (.A1(_0785_),
    .A2(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1619_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_0571_),
    .A3(_0573_),
    .B1(_0567_),
    .B2(_0569_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1620_ (.I0(B),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1621_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1622_ (.I(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1623_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .A2(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1624_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .A2(_0574_),
    .B(_0577_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1625_ (.I0(E6END[1]),
    .I1(SS4END[1]),
    .I2(W2END[1]),
    .I3(W6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1626_ (.I(_0579_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1627_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .A2(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1628_ (.I0(N2END[1]),
    .I1(E1END[3]),
    .I2(N4END[1]),
    .I3(E2END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1629_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .A2(_0582_),
    .B(_0581_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1630_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ),
    .A2(_0583_),
    .B(_0578_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1631_ (.I0(E1END[2]),
    .I1(W1END[2]),
    .I2(A),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1632_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_0584_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1633_ (.I0(C),
    .I1(D),
    .I2(E),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1634_ (.A1(_0786_),
    .A2(_0586_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1635_ (.I0(_0018_),
    .I1(_0142_),
    .I2(_0204_),
    .I3(_0398_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1636_ (.A1(_0786_),
    .A2(_0588_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1637_ (.I0(G),
    .I1(H),
    .I2(\Inst_LUT4AB_switch_matrix.M_AD ),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1638_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_0590_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1639_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ),
    .A2(_0585_),
    .A3(_0587_),
    .B1(_0589_),
    .B2(_0591_),
    .ZN(\Inst_LUT4AB_switch_matrix.W6BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1640_ (.I0(E1END[3]),
    .I1(W1END[3]),
    .I2(A),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1641_ (.I0(C),
    .I1(D),
    .I2(E),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1642_ (.I0(_0800_),
    .I1(_0110_),
    .I2(_0192_),
    .I3(_0385_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1643_ (.I0(G),
    .I1(H),
    .I2(\Inst_LUT4AB_switch_matrix.M_AB ),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1644_ (.I0(_0592_),
    .I1(_0593_),
    .I2(_0595_),
    .I3(_0594_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.W6BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1645_ (.I0(E),
    .I1(_0204_),
    .I2(_0398_),
    .I3(_0851_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1646_ (.I0(N1END[1]),
    .I1(S1END[1]),
    .I2(W1END[1]),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1647_ (.I0(_0597_),
    .I1(_0596_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.WW4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1648_ (.I0(C),
    .I1(_0192_),
    .I2(_0385_),
    .I3(_0133_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1649_ (.I0(N1END[0]),
    .I1(W1END[0]),
    .I2(S1END[0]),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1650_ (.I0(_0599_),
    .I1(_0598_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.WW4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1651_ (.I0(H),
    .I1(_0018_),
    .I2(_0142_),
    .I3(_0195_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1652_ (.I0(N1END[3]),
    .I1(S1END[3]),
    .I2(W1END[3]),
    .I3(A),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1653_ (.I0(_0601_),
    .I1(_0600_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.WW4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1654_ (.I0(G),
    .I1(_0800_),
    .I2(_0110_),
    .I3(_0389_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1655_ (.I0(N1END[2]),
    .I1(S1END[2]),
    .I2(W1END[2]),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1656_ (.I0(_0603_),
    .I1(_0602_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.WW4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1657_ (.I0(E),
    .I1(_0204_),
    .I2(_0398_),
    .I3(_0036_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1658_ (.I0(N1END[1]),
    .I1(E1END[1]),
    .I2(W1END[1]),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1659_ (.I0(_0605_),
    .I1(_0604_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.SS4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1660_ (.I0(C),
    .I1(_0192_),
    .I2(_0385_),
    .I3(_0290_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1661_ (.I0(N1END[0]),
    .I1(W1END[0]),
    .I2(E1END[0]),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1662_ (.I0(_0607_),
    .I1(_0606_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.SS4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1663_ (.I0(H),
    .I1(_0018_),
    .I2(_0142_),
    .I3(_0215_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1664_ (.I0(N1END[3]),
    .I1(E1END[3]),
    .I2(W1END[3]),
    .I3(A),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1665_ (.I0(_0609_),
    .I1(_0608_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.SS4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1666_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_0409_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1667_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_0110_),
    .B(_0610_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1668_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_0799_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1669_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(G),
    .B(_0612_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1670_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .A2(_0613_),
    .B(_0611_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1671_ (.I0(N1END[2]),
    .I1(W1END[2]),
    .I2(E1END[2]),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1672_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ),
    .A2(_0615_),
    .B(_0614_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1673_ (.I(_0616_),
    .ZN(\Inst_LUT4AB_switch_matrix.SS4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1674_ (.I0(E1END[2]),
    .I1(W1END[2]),
    .I2(A),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1675_ (.I0(C),
    .I1(D),
    .I2(E),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1676_ (.I0(_0617_),
    .I1(_0618_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1677_ (.I0(G),
    .I1(H),
    .I2(\Inst_LUT4AB_switch_matrix.M_AD ),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1678_ (.I0(_0018_),
    .I1(_0142_),
    .I2(_0204_),
    .I3(_0398_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1679_ (.I0(_0620_),
    .I1(_0621_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1680_ (.I0(_0619_),
    .I1(_0622_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.E6BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1681_ (.I0(E1END[3]),
    .I1(W1END[3]),
    .I2(A),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1682_ (.I0(C),
    .I1(D),
    .I2(E),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1683_ (.I0(_0800_),
    .I1(_0110_),
    .I2(_0192_),
    .I3(_0385_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1684_ (.I0(G),
    .I1(H),
    .I2(\Inst_LUT4AB_switch_matrix.M_AB ),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1685_ (.I0(_0623_),
    .I1(_0624_),
    .I2(_0626_),
    .I3(_0625_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.E6BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1686_ (.I0(E),
    .I1(_0204_),
    .I2(_0398_),
    .I3(_0831_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1687_ (.I0(N1END[1]),
    .I1(E1END[1]),
    .I2(S1END[1]),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1688_ (.I0(_0628_),
    .I1(_0627_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.EE4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1689_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .A2(_0266_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1690_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .A2(_0385_),
    .B(_0629_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1691_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .A2(_0191_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1692_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .A2(C),
    .B(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1693_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .A2(_0632_),
    .B(_0630_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1694_ (.I0(N1END[0]),
    .I1(S1END[0]),
    .I2(E1END[0]),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1695_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ),
    .A2(_0634_),
    .B(_0633_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1696_ (.I(_0635_),
    .ZN(\Inst_LUT4AB_switch_matrix.EE4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1697_ (.I0(H),
    .I1(_0018_),
    .I2(_0142_),
    .I3(_0158_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1698_ (.I0(N1END[3]),
    .I1(E1END[3]),
    .I2(S1END[3]),
    .I3(A),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1699_ (.I0(_0637_),
    .I1(_0636_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.EE4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1700_ (.I0(G),
    .I1(_0800_),
    .I2(_0110_),
    .I3(_0366_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1701_ (.I0(N1END[2]),
    .I1(S1END[2]),
    .I2(E1END[2]),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1702_ (.I0(_0639_),
    .I1(_0638_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.EE4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1703_ (.I0(E),
    .I1(_0204_),
    .I2(_0398_),
    .I3(_0810_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1704_ (.I0(N1END[1]),
    .I1(E1END[1]),
    .I2(W1END[1]),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1705_ (.I0(_0641_),
    .I1(_0640_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.NN4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1706_ (.I0(C),
    .I1(_0192_),
    .I2(_0385_),
    .I3(_0121_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1707_ (.I0(N1END[0]),
    .I1(W1END[0]),
    .I2(E1END[0]),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1708_ (.I0(_0643_),
    .I1(_0642_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.NN4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1709_ (.I0(H),
    .I1(_0018_),
    .I2(_0142_),
    .I3(_0178_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1710_ (.I0(N1END[3]),
    .I1(E1END[3]),
    .I2(W1END[3]),
    .I3(A),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1711_ (.I0(_0645_),
    .I1(_0644_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.NN4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1712_ (.I0(G),
    .I1(_0800_),
    .I2(_0110_),
    .I3(_0375_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1713_ (.I0(N1END[2]),
    .I1(W1END[2]),
    .I2(E1END[2]),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1714_ (.I0(_0647_),
    .I1(_0646_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.NN4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1715_ (.I0(A),
    .I1(_0020_),
    .I2(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .I3(_0830_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.W1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1716_ (.I0(H),
    .I1(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .I2(_0385_),
    .I3(_0405_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.W1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1717_ (.I0(G),
    .I1(_0173_),
    .I2(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .I3(_0194_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.W1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1718_ (.I0(F),
    .I1(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .I2(_0301_),
    .I3(_0120_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.W1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1719_ (.I0(S2END[1]),
    .I1(S4END[0]),
    .I2(W6END[0]),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1720_ (.I0(S2END[0]),
    .I1(W6END[1]),
    .I2(S4END[3]),
    .I3(C),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1721_ (.I0(E6END[0]),
    .I1(S4END[2]),
    .I2(S2END[3]),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1722_ (.I0(E6END[1]),
    .I1(S4END[1]),
    .I2(S2END[2]),
    .I3(A),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1723_ (.I0(H),
    .I1(_0020_),
    .I2(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .I3(_0830_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1724_ (.I0(G),
    .I1(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .I2(_0385_),
    .I3(_0405_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1725_ (.I0(F),
    .I1(_0173_),
    .I2(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .I3(_0194_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1726_ (.I0(E),
    .I1(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .I2(_0301_),
    .I3(_0120_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1727_ (.I0(G),
    .I1(_0020_),
    .I2(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .I3(_0830_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.E1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1728_ (.I0(F),
    .I1(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .I2(_0385_),
    .I3(_0405_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.E1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1729_ (.I0(E),
    .I1(_0173_),
    .I2(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .I3(_0194_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.E1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1730_ (.I0(D),
    .I1(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .I2(_0301_),
    .I3(_0120_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.E1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1731_ (.I0(N2END[1]),
    .I1(W6END[0]),
    .I2(N4END[0]),
    .I3(H),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1732_ (.I0(N2END[0]),
    .I1(N4END[3]),
    .I2(W6END[1]),
    .I3(G),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1733_ (.I0(N2END[3]),
    .I1(N4END[2]),
    .I2(E6END[0]),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1734_ (.I0(N2END[2]),
    .I1(N4END[1]),
    .I2(E6END[1]),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1735_ (.I0(F),
    .I1(_0020_),
    .I2(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .I3(_0830_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1736_ (.I0(E),
    .I1(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .I2(_0385_),
    .I3(_0405_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1737_ (.I0(D),
    .I1(_0173_),
    .I2(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .I3(_0194_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1738_ (.I0(C),
    .I1(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .I2(_0301_),
    .I3(_0120_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1739_ (.A1(_0401_),
    .A2(_0430_),
    .B(_0445_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1740_ (.A1(_0444_),
    .A2(_0648_),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1741_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0419_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1742_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0047_),
    .B(_0649_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1743_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0301_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1744_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0227_),
    .B(_0651_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1745_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1746_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0119_),
    .B(_0653_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1747_ (.A1(_0284_),
    .A2(_0288_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1748_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .B(_0655_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1749_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1750_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_0650_),
    .A3(_0652_),
    .B1(_0654_),
    .B2(_0657_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1751_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ),
    .A2(_0658_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1752_ (.A1(_0733_),
    .A2(_0363_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1753_ (.A1(_0733_),
    .A2(_0821_),
    .B(_0660_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1754_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(_0252_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1755_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(_0172_),
    .B(_0662_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1756_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ),
    .A2(_0663_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1757_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1758_ (.A1(_0733_),
    .A2(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .B(_0665_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1759_ (.A1(_0733_),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1760_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_0667_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1761_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .B(_0668_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1762_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ),
    .A2(_0666_),
    .A3(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1763_ (.A1(_0661_),
    .A2(_0664_),
    .B(_0670_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1764_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ),
    .A2(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1765_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ),
    .A2(_0671_),
    .B(_0460_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1766_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0672_),
    .B(_0659_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1767_ (.A1(_0776_),
    .A2(_0659_),
    .B1(_0673_),
    .B2(_0674_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1768_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ),
    .A2(_0671_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1769_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ),
    .A2(_0658_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1770_ (.A1(_0063_),
    .A2(_0675_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1771_ (.A1(\Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0675_),
    .B(_0676_),
    .C(_0677_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1772_ (.A1(_0734_),
    .A2(_0676_),
    .B(_0678_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1773_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ),
    .A2(_0658_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1774_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ),
    .A2(_0671_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1775_ (.I0(\Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ),
    .I1(_0100_),
    .S(_0680_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1776_ (.I0(_0681_),
    .I1(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(_0679_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1777_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ),
    .A2(_0658_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1778_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .A2(_0682_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1779_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ),
    .A2(_0671_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1780_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ),
    .A2(_0671_),
    .B(_0316_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1781_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0684_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1782_ (.A1(_0682_),
    .A2(_0685_),
    .A3(_0686_),
    .B(_0683_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1783_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ),
    .A2(_0658_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1784_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .A2(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1785_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ),
    .A2(_0671_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1786_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ),
    .A2(_0671_),
    .B(_0495_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1787_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0689_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1788_ (.A1(_0687_),
    .A2(_0690_),
    .A3(_0691_),
    .B(_0688_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1789_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ),
    .A2(_0658_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1790_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .A2(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1791_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ),
    .A2(_0671_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1792_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ),
    .A2(_0671_),
    .B(_0238_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1793_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0694_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1794_ (.A1(_0692_),
    .A2(_0695_),
    .A3(_0696_),
    .B(_0693_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1795_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ),
    .A2(_0658_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1796_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .A2(_0697_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1797_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ),
    .A2(_0671_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1798_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ),
    .A2(_0671_),
    .B(_0348_),
    .C(_0340_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1799_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0699_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1800_ (.A1(_0697_),
    .A2(_0700_),
    .A3(_0701_),
    .B(_0698_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1801_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ),
    .A2(_0658_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1802_ (.A1(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .A2(_0702_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1803_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ),
    .A2(_0671_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1804_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ),
    .A2(_0671_),
    .B(_0429_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1805_ (.A1(\Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0704_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1806_ (.A1(_0702_),
    .A2(_0705_),
    .A3(_0706_),
    .B(_0703_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1807_ (.D(FrameData[24]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1808_ (.D(FrameData[25]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1809_ (.D(FrameData[26]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1810_ (.D(FrameData[27]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1811_ (.D(FrameData[28]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1812_ (.D(FrameData[29]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1813_ (.D(FrameData[30]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1814_ (.D(FrameData[31]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1815_ (.D(FrameData[0]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1816_ (.D(FrameData[1]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1817_ (.D(FrameData[2]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1818_ (.D(FrameData[3]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1819_ (.D(FrameData[4]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1820_ (.D(FrameData[5]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1821_ (.D(FrameData[6]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1822_ (.D(FrameData[7]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1823_ (.D(FrameData[8]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1824_ (.D(FrameData[9]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1825_ (.D(FrameData[10]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1826_ (.D(FrameData[11]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1827_ (.D(FrameData[12]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1828_ (.D(FrameData[13]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1829_ (.D(FrameData[14]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1830_ (.D(FrameData[15]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1831_ (.D(FrameData[16]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1832_ (.D(FrameData[17]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1833_ (.D(FrameData[18]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1834_ (.D(FrameData[19]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1835_ (.D(FrameData[20]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1836_ (.D(FrameData[21]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1837_ (.D(FrameData[22]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1838_ (.D(FrameData[23]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1839_ (.D(FrameData[24]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1840_ (.D(FrameData[25]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1841_ (.D(FrameData[26]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1842_ (.D(FrameData[27]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1843_ (.D(FrameData[28]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1844_ (.D(FrameData[29]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1845_ (.D(FrameData[30]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1846_ (.D(FrameData[31]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1847_ (.D(FrameData[0]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1848_ (.D(FrameData[1]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1849_ (.D(FrameData[2]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1850_ (.D(FrameData[3]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1851_ (.D(FrameData[4]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1852_ (.D(FrameData[5]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1853_ (.D(FrameData[6]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1854_ (.D(FrameData[7]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1855_ (.D(FrameData[8]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1856_ (.D(FrameData[9]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1857_ (.D(FrameData[10]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1858_ (.D(FrameData[11]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1859_ (.D(FrameData[12]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1860_ (.D(FrameData[13]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1861_ (.D(FrameData[14]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1862_ (.D(FrameData[15]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1863_ (.D(FrameData[16]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1864_ (.D(FrameData[17]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1865_ (.D(FrameData[18]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1866_ (.D(FrameData[19]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1867_ (.D(FrameData[20]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1868_ (.D(FrameData[21]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1869_ (.D(FrameData[22]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1870_ (.D(FrameData[23]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1871_ (.D(FrameData[24]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1872_ (.D(FrameData[25]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1873_ (.D(FrameData[26]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1874_ (.D(FrameData[27]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1875_ (.D(FrameData[28]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1876_ (.D(FrameData[29]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1877_ (.D(FrameData[30]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1878_ (.D(FrameData[31]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1879_ (.D(FrameData[0]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1880_ (.D(FrameData[1]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1881_ (.D(FrameData[2]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1882_ (.D(FrameData[3]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1883_ (.D(FrameData[4]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1884_ (.D(FrameData[5]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1885_ (.D(FrameData[6]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1886_ (.D(FrameData[7]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1887_ (.D(FrameData[8]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1888_ (.D(FrameData[9]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1889_ (.D(FrameData[10]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1890_ (.D(FrameData[11]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1891_ (.D(FrameData[12]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1892_ (.D(FrameData[13]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1893_ (.D(FrameData[14]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1894_ (.D(FrameData[15]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1895_ (.D(FrameData[16]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1896_ (.D(FrameData[17]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1897_ (.D(FrameData[18]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1898_ (.D(FrameData[19]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1899_ (.D(FrameData[20]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1900_ (.D(FrameData[21]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1901_ (.D(FrameData[22]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1902_ (.D(FrameData[23]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1903_ (.D(FrameData[24]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1904_ (.D(FrameData[25]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1905_ (.D(FrameData[26]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1906_ (.D(FrameData[27]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1907_ (.D(FrameData[28]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1908_ (.D(FrameData[29]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1909_ (.D(FrameData[30]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1910_ (.D(FrameData[31]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1911_ (.D(FrameData[0]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1912_ (.D(FrameData[1]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1913_ (.D(FrameData[2]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1914_ (.D(FrameData[3]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1915_ (.D(FrameData[4]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1916_ (.D(FrameData[5]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1917_ (.D(FrameData[6]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1918_ (.D(FrameData[7]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1919_ (.D(FrameData[8]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1920_ (.D(FrameData[9]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1921_ (.D(FrameData[10]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1922_ (.D(FrameData[11]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1923_ (.D(FrameData[12]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1924_ (.D(FrameData[13]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1925_ (.D(FrameData[14]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1926_ (.D(FrameData[15]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1927_ (.D(FrameData[16]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1928_ (.D(FrameData[17]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1929_ (.D(FrameData[18]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1930_ (.D(FrameData[19]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1931_ (.D(FrameData[20]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1932_ (.D(FrameData[21]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1933_ (.D(FrameData[22]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1934_ (.D(FrameData[23]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1935_ (.D(FrameData[24]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1936_ (.D(FrameData[25]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1937_ (.D(FrameData[26]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1938_ (.D(FrameData[27]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1939_ (.D(FrameData[28]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1940_ (.D(FrameData[29]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1941_ (.D(FrameData[30]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1942_ (.D(FrameData[31]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1943_ (.D(FrameData[0]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1944_ (.D(FrameData[1]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1945_ (.D(FrameData[2]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1946_ (.D(FrameData[3]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1947_ (.D(FrameData[4]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1948_ (.D(FrameData[5]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1949_ (.D(FrameData[6]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1950_ (.D(FrameData[7]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1951_ (.D(FrameData[8]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1952_ (.D(FrameData[9]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1953_ (.D(FrameData[10]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1954_ (.D(FrameData[11]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1955_ (.D(FrameData[12]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1956_ (.D(FrameData[13]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1957_ (.D(FrameData[14]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1958_ (.D(FrameData[15]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1959_ (.D(FrameData[16]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1960_ (.D(FrameData[17]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1961_ (.D(FrameData[18]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1962_ (.D(FrameData[19]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1963_ (.D(FrameData[20]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1964_ (.D(FrameData[21]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1965_ (.D(FrameData[22]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1966_ (.D(FrameData[23]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1967_ (.D(FrameData[24]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1968_ (.D(FrameData[25]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1969_ (.D(FrameData[26]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1970_ (.D(FrameData[27]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1971_ (.D(FrameData[28]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1972_ (.D(FrameData[29]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1973_ (.D(FrameData[30]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1974_ (.D(FrameData[31]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1975_ (.D(FrameData[0]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1976_ (.D(FrameData[1]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1977_ (.D(FrameData[2]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1978_ (.D(FrameData[3]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1979_ (.D(FrameData[4]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1980_ (.D(FrameData[5]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1981_ (.D(FrameData[6]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1982_ (.D(FrameData[7]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1983_ (.D(FrameData[8]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1984_ (.D(FrameData[9]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1985_ (.D(FrameData[10]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1986_ (.D(FrameData[11]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1987_ (.D(FrameData[12]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1988_ (.D(FrameData[13]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1989_ (.D(FrameData[14]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1990_ (.D(FrameData[15]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1991_ (.D(FrameData[16]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1992_ (.D(FrameData[17]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1993_ (.D(FrameData[18]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1994_ (.D(FrameData[19]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1995_ (.D(FrameData[20]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1996_ (.D(FrameData[21]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1997_ (.D(FrameData[22]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1998_ (.D(FrameData[23]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1999_ (.D(FrameData[24]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2000_ (.D(FrameData[25]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2001_ (.D(FrameData[26]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2002_ (.D(FrameData[27]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2003_ (.D(FrameData[28]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2004_ (.D(FrameData[29]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2005_ (.D(FrameData[30]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2006_ (.D(FrameData[31]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2007_ (.D(FrameData[0]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2008_ (.D(FrameData[1]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2009_ (.D(FrameData[2]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2010_ (.D(FrameData[3]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2011_ (.D(FrameData[4]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2012_ (.D(FrameData[5]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2013_ (.D(FrameData[6]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2014_ (.D(FrameData[7]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2015_ (.D(FrameData[8]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2016_ (.D(FrameData[9]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2017_ (.D(FrameData[10]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2018_ (.D(FrameData[11]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2019_ (.D(FrameData[12]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2020_ (.D(FrameData[13]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2021_ (.D(FrameData[14]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2022_ (.D(FrameData[15]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2023_ (.D(FrameData[16]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2024_ (.D(FrameData[17]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2025_ (.D(FrameData[18]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2026_ (.D(FrameData[19]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2027_ (.D(FrameData[20]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2028_ (.D(FrameData[21]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2029_ (.D(FrameData[22]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2030_ (.D(FrameData[23]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2031_ (.D(FrameData[24]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2032_ (.D(FrameData[25]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2033_ (.D(FrameData[26]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2034_ (.D(FrameData[27]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2035_ (.D(FrameData[28]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2036_ (.D(FrameData[29]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2037_ (.D(FrameData[30]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2038_ (.D(FrameData[31]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2039_ (.D(FrameData[0]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2040_ (.D(FrameData[1]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2041_ (.D(FrameData[2]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2042_ (.D(FrameData[3]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2043_ (.D(FrameData[4]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2044_ (.D(FrameData[5]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2045_ (.D(FrameData[6]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2046_ (.D(FrameData[7]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2047_ (.D(FrameData[8]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2048_ (.D(FrameData[9]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2049_ (.D(FrameData[10]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2050_ (.D(FrameData[11]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2051_ (.D(FrameData[12]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2052_ (.D(FrameData[13]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2053_ (.D(FrameData[14]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2054_ (.D(FrameData[15]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2055_ (.D(FrameData[16]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2056_ (.D(FrameData[17]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2057_ (.D(FrameData[18]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2058_ (.D(FrameData[19]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2059_ (.D(FrameData[20]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2060_ (.D(FrameData[21]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2061_ (.D(FrameData[22]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2062_ (.D(FrameData[23]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2063_ (.D(FrameData[24]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2064_ (.D(FrameData[25]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2065_ (.D(FrameData[26]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2066_ (.D(FrameData[27]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2067_ (.D(FrameData[28]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2068_ (.D(FrameData[29]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2069_ (.D(FrameData[30]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2070_ (.D(FrameData[31]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2071_ (.D(FrameData[0]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2072_ (.D(FrameData[1]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2073_ (.D(FrameData[2]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2074_ (.D(FrameData[3]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2075_ (.D(FrameData[4]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2076_ (.D(FrameData[5]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2077_ (.D(FrameData[6]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2078_ (.D(FrameData[7]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2079_ (.D(FrameData[8]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2080_ (.D(FrameData[9]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2081_ (.D(FrameData[10]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2082_ (.D(FrameData[11]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2083_ (.D(FrameData[12]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2084_ (.D(FrameData[13]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2085_ (.D(FrameData[14]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2086_ (.D(FrameData[15]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2087_ (.D(FrameData[16]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2088_ (.D(FrameData[17]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2089_ (.D(FrameData[18]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2090_ (.D(FrameData[19]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2091_ (.D(FrameData[20]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2092_ (.D(FrameData[21]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2093_ (.D(FrameData[22]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2094_ (.D(FrameData[23]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2095_ (.D(FrameData[24]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2096_ (.D(FrameData[25]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2097_ (.D(FrameData[26]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2098_ (.D(FrameData[27]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2099_ (.D(FrameData[28]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2100_ (.D(FrameData[29]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2101_ (.D(FrameData[30]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2102_ (.D(FrameData[31]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2103_ (.D(FrameData[0]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2104_ (.D(FrameData[1]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2105_ (.D(FrameData[2]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2106_ (.D(FrameData[3]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2107_ (.D(FrameData[4]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2108_ (.D(FrameData[5]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2109_ (.D(FrameData[6]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2110_ (.D(FrameData[7]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2111_ (.D(FrameData[8]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2112_ (.D(FrameData[9]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2113_ (.D(FrameData[10]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2114_ (.D(FrameData[11]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2115_ (.D(FrameData[12]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2116_ (.D(FrameData[13]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2117_ (.D(FrameData[14]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2118_ (.D(FrameData[15]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2119_ (.D(FrameData[16]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2120_ (.D(FrameData[17]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2121_ (.D(FrameData[18]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2122_ (.D(FrameData[19]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2123_ (.D(FrameData[20]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2124_ (.D(FrameData[21]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2125_ (.D(FrameData[22]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2126_ (.D(FrameData[23]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2127_ (.D(FrameData[24]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2128_ (.D(FrameData[25]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2129_ (.D(FrameData[26]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2130_ (.D(FrameData[27]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2131_ (.D(FrameData[28]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2132_ (.D(FrameData[29]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2133_ (.D(FrameData[30]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2134_ (.D(FrameData[31]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2135_ (.D(FrameData[0]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2136_ (.D(FrameData[1]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2137_ (.D(FrameData[2]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2138_ (.D(FrameData[3]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2139_ (.D(FrameData[4]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2140_ (.D(FrameData[5]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2141_ (.D(FrameData[6]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2142_ (.D(FrameData[7]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2143_ (.D(FrameData[8]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2144_ (.D(FrameData[9]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2145_ (.D(FrameData[10]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2146_ (.D(FrameData[11]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2147_ (.D(FrameData[12]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2148_ (.D(FrameData[13]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2149_ (.D(FrameData[14]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2150_ (.D(FrameData[15]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2151_ (.D(FrameData[16]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2152_ (.D(FrameData[17]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2153_ (.D(FrameData[18]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2154_ (.D(FrameData[19]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2155_ (.D(FrameData[20]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2156_ (.D(FrameData[21]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2157_ (.D(FrameData[22]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2158_ (.D(FrameData[23]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2159_ (.D(FrameData[24]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2160_ (.D(FrameData[25]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2161_ (.D(FrameData[26]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2162_ (.D(FrameData[27]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2163_ (.D(FrameData[28]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2164_ (.D(FrameData[29]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2165_ (.D(FrameData[30]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2166_ (.D(FrameData[31]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2167_ (.D(FrameData[0]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2168_ (.D(FrameData[1]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2169_ (.D(FrameData[2]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2170_ (.D(FrameData[3]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2171_ (.D(FrameData[4]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2172_ (.D(FrameData[5]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2173_ (.D(FrameData[6]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2174_ (.D(FrameData[7]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2175_ (.D(FrameData[8]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2176_ (.D(FrameData[9]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2177_ (.D(FrameData[10]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2178_ (.D(FrameData[11]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2179_ (.D(FrameData[12]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2180_ (.D(FrameData[13]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2181_ (.D(FrameData[14]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2182_ (.D(FrameData[15]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2183_ (.D(FrameData[16]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2184_ (.D(FrameData[17]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2185_ (.D(FrameData[18]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2186_ (.D(FrameData[19]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2187_ (.D(FrameData[20]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2188_ (.D(FrameData[21]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2189_ (.D(FrameData[22]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2190_ (.D(FrameData[23]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2191_ (.D(FrameData[24]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2192_ (.D(FrameData[25]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2193_ (.D(FrameData[26]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2194_ (.D(FrameData[27]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2195_ (.D(FrameData[28]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2196_ (.D(FrameData[29]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2197_ (.D(FrameData[30]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2198_ (.D(FrameData[31]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2199_ (.D(FrameData[0]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2200_ (.D(FrameData[1]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2201_ (.D(FrameData[2]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2202_ (.D(FrameData[3]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2203_ (.D(FrameData[4]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2204_ (.D(FrameData[5]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2205_ (.D(FrameData[6]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2206_ (.D(FrameData[7]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2207_ (.D(FrameData[8]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2208_ (.D(FrameData[9]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2209_ (.D(FrameData[10]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2210_ (.D(FrameData[11]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2211_ (.D(FrameData[12]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2212_ (.D(FrameData[13]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2213_ (.D(FrameData[14]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2214_ (.D(FrameData[15]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2215_ (.D(FrameData[16]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2216_ (.D(FrameData[17]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2217_ (.D(FrameData[18]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2218_ (.D(FrameData[19]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2219_ (.D(FrameData[20]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2220_ (.D(FrameData[21]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2221_ (.D(FrameData[22]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2222_ (.D(FrameData[23]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2223_ (.D(FrameData[24]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2224_ (.D(FrameData[25]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2225_ (.D(FrameData[26]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2226_ (.D(FrameData[27]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2227_ (.D(FrameData[28]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2228_ (.D(FrameData[29]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2229_ (.D(FrameData[30]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2230_ (.D(FrameData[31]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2231_ (.D(FrameData[0]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2232_ (.D(FrameData[1]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2233_ (.D(FrameData[2]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2234_ (.D(FrameData[3]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2235_ (.D(FrameData[4]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2236_ (.D(FrameData[5]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2237_ (.D(FrameData[6]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2238_ (.D(FrameData[7]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2239_ (.D(FrameData[8]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2240_ (.D(FrameData[9]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2241_ (.D(FrameData[10]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2242_ (.D(FrameData[11]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2243_ (.D(FrameData[12]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2244_ (.D(FrameData[13]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2245_ (.D(FrameData[14]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2246_ (.D(FrameData[15]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2247_ (.D(FrameData[16]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2248_ (.D(FrameData[17]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2249_ (.D(FrameData[18]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2250_ (.D(FrameData[19]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2251_ (.D(FrameData[20]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2252_ (.D(FrameData[21]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2253_ (.D(FrameData[22]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2254_ (.D(FrameData[23]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2255_ (.D(FrameData[24]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2256_ (.D(FrameData[25]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2257_ (.D(FrameData[26]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2258_ (.D(FrameData[27]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2259_ (.D(FrameData[28]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2260_ (.D(FrameData[29]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2261_ (.D(FrameData[30]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2262_ (.D(FrameData[31]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2263_ (.D(FrameData[0]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2264_ (.D(FrameData[1]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2265_ (.D(FrameData[2]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2266_ (.D(FrameData[3]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2267_ (.D(FrameData[4]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2268_ (.D(FrameData[5]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2269_ (.D(FrameData[6]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2270_ (.D(FrameData[7]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2271_ (.D(FrameData[8]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2272_ (.D(FrameData[9]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2273_ (.D(FrameData[10]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2274_ (.D(FrameData[11]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2275_ (.D(FrameData[12]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2276_ (.D(FrameData[13]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2277_ (.D(FrameData[14]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2278_ (.D(FrameData[15]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2279_ (.D(FrameData[16]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2280_ (.D(FrameData[17]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2281_ (.D(FrameData[18]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2282_ (.D(FrameData[19]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2283_ (.D(FrameData[20]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2284_ (.D(FrameData[21]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2285_ (.D(FrameData[22]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2286_ (.D(FrameData[23]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2287_ (.D(FrameData[24]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2288_ (.D(FrameData[25]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2289_ (.D(FrameData[26]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2290_ (.D(FrameData[27]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2291_ (.D(FrameData[28]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2292_ (.D(FrameData[29]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2293_ (.D(FrameData[30]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2294_ (.D(FrameData[31]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2295_ (.D(FrameData[0]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2296_ (.D(FrameData[1]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2297_ (.D(FrameData[2]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2298_ (.D(FrameData[3]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2299_ (.D(FrameData[4]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2300_ (.D(FrameData[5]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2301_ (.D(FrameData[6]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2302_ (.D(FrameData[7]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2303_ (.D(FrameData[8]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2304_ (.D(FrameData[9]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2305_ (.D(FrameData[10]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2306_ (.D(FrameData[11]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2307_ (.D(FrameData[12]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2308_ (.D(FrameData[13]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2309_ (.D(FrameData[14]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2310_ (.D(FrameData[15]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2311_ (.D(FrameData[16]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2312_ (.D(FrameData[17]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2313_ (.D(FrameData[18]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2314_ (.D(FrameData[19]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2315_ (.D(FrameData[20]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2316_ (.D(FrameData[21]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2317_ (.D(FrameData[22]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2318_ (.D(FrameData[23]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2319_ (.D(FrameData[24]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2320_ (.D(FrameData[25]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2321_ (.D(FrameData[26]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2322_ (.D(FrameData[27]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2323_ (.D(FrameData[28]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2324_ (.D(FrameData[29]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2325_ (.D(FrameData[30]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2326_ (.D(FrameData[31]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2327_ (.D(FrameData[0]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2328_ (.D(FrameData[1]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2329_ (.D(FrameData[2]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2330_ (.D(FrameData[3]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2331_ (.D(FrameData[4]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2332_ (.D(FrameData[5]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2333_ (.D(FrameData[6]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2334_ (.D(FrameData[7]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2335_ (.D(FrameData[8]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2336_ (.D(FrameData[9]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2337_ (.D(FrameData[10]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2338_ (.D(FrameData[11]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2339_ (.D(FrameData[12]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2340_ (.D(FrameData[13]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2341_ (.D(FrameData[14]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2342_ (.D(FrameData[15]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2343_ (.D(FrameData[16]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2344_ (.D(FrameData[17]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2345_ (.D(FrameData[18]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2346_ (.D(FrameData[19]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2347_ (.D(FrameData[20]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2348_ (.D(FrameData[21]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2349_ (.D(FrameData[22]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2350_ (.D(FrameData[23]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2351_ (.D(FrameData[24]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2352_ (.D(FrameData[25]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2353_ (.D(FrameData[26]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2354_ (.D(FrameData[27]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2355_ (.D(FrameData[28]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2356_ (.D(FrameData[29]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2357_ (.D(FrameData[30]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2358_ (.D(FrameData[31]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2359_ (.D(FrameData[0]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2360_ (.D(FrameData[1]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2361_ (.D(FrameData[2]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2362_ (.D(FrameData[3]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2363_ (.D(FrameData[4]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2364_ (.D(FrameData[5]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2365_ (.D(FrameData[6]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2366_ (.D(FrameData[7]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2367_ (.D(FrameData[8]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2368_ (.D(FrameData[9]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2369_ (.D(FrameData[10]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2370_ (.D(FrameData[11]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2371_ (.D(FrameData[12]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2372_ (.D(FrameData[13]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2373_ (.D(FrameData[14]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2374_ (.D(FrameData[15]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2375_ (.D(FrameData[16]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2376_ (.D(FrameData[17]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2377_ (.D(FrameData[18]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2378_ (.D(FrameData[19]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2379_ (.D(FrameData[20]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2380_ (.D(FrameData[21]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2381_ (.D(FrameData[22]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2382_ (.D(FrameData[23]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2383_ (.D(FrameData[24]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2384_ (.D(FrameData[25]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2385_ (.D(FrameData[26]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2386_ (.D(FrameData[27]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2387_ (.D(FrameData[28]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2388_ (.D(FrameData[29]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2389_ (.D(FrameData[30]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2390_ (.D(FrameData[31]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2391_ (.D(FrameData[0]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2392_ (.D(FrameData[1]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2393_ (.D(FrameData[2]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2394_ (.D(FrameData[3]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2395_ (.D(FrameData[4]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2396_ (.D(FrameData[5]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2397_ (.D(FrameData[6]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2398_ (.D(FrameData[7]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2399_ (.D(FrameData[8]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2400_ (.D(FrameData[9]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2401_ (.D(FrameData[10]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2402_ (.D(FrameData[11]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2403_ (.D(FrameData[12]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2404_ (.D(FrameData[13]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2405_ (.D(FrameData[14]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2406_ (.D(FrameData[15]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2407_ (.D(FrameData[16]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2408_ (.D(FrameData[17]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2409_ (.D(FrameData[18]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2410_ (.D(FrameData[19]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2411_ (.D(FrameData[20]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2412_ (.D(FrameData[21]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2413_ (.D(FrameData[22]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2414_ (.D(FrameData[23]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2415_ (.D(FrameData[24]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2416_ (.D(FrameData[25]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2417_ (.D(FrameData[26]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2418_ (.D(FrameData[27]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2419_ (.D(FrameData[28]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2420_ (.D(FrameData[29]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2421_ (.D(FrameData[30]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2422_ (.D(FrameData[31]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2423_ (.D(_0000_),
    .CLK(clknet_1_1__leaf_UserCLK_regs),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2424_ (.D(_0001_),
    .CLK(clknet_1_0__leaf_UserCLK_regs),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2425_ (.D(_0002_),
    .CLK(clknet_1_0__leaf_UserCLK_regs),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2426_ (.D(_0003_),
    .CLK(clknet_1_0__leaf_UserCLK_regs),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2427_ (.D(_0004_),
    .CLK(clknet_1_0__leaf_UserCLK_regs),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2428_ (.D(_0005_),
    .CLK(clknet_1_1__leaf_UserCLK_regs),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2429_ (.D(_0006_),
    .CLK(clknet_1_1__leaf_UserCLK_regs),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2430_ (.D(_0007_),
    .CLK(clknet_1_1__leaf_UserCLK_regs),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2431_ (.I(\Inst_LUT4AB_switch_matrix.E1BEG0 ),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2432_ (.I(\Inst_LUT4AB_switch_matrix.E1BEG1 ),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2433_ (.I(\Inst_LUT4AB_switch_matrix.E1BEG2 ),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2434_ (.I(\Inst_LUT4AB_switch_matrix.E1BEG3 ),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2435_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2436_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2437_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2438_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2439_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2440_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2441_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2442_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2443_ (.I(E2MID[0]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2444_ (.I(E2MID[1]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2445_ (.I(E2MID[2]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2446_ (.I(E2MID[3]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2447_ (.I(E2MID[4]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2448_ (.I(E2MID[5]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2449_ (.I(E2MID[6]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2450_ (.I(E2MID[7]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2451_ (.I(E6END[2]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2452_ (.I(E6END[3]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2453_ (.I(E6END[4]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2454_ (.I(E6END[5]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2455_ (.I(E6END[6]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2456_ (.I(E6END[7]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2457_ (.I(E6END[8]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2458_ (.I(E6END[9]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2459_ (.I(E6END[10]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2460_ (.I(E6END[11]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2461_ (.I(\Inst_LUT4AB_switch_matrix.E6BEG0 ),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2462_ (.I(\Inst_LUT4AB_switch_matrix.E6BEG1 ),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2463_ (.I(EE4END[4]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2464_ (.I(EE4END[5]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2465_ (.I(EE4END[6]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2466_ (.I(EE4END[7]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2467_ (.I(EE4END[8]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2468_ (.I(EE4END[9]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2469_ (.I(EE4END[10]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2470_ (.I(EE4END[11]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2471_ (.I(EE4END[12]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2472_ (.I(EE4END[13]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2473_ (.I(EE4END[14]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2474_ (.I(EE4END[15]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2475_ (.I(\Inst_LUT4AB_switch_matrix.EE4BEG0 ),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2476_ (.I(\Inst_LUT4AB_switch_matrix.EE4BEG1 ),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2477_ (.I(\Inst_LUT4AB_switch_matrix.EE4BEG2 ),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2478_ (.I(\Inst_LUT4AB_switch_matrix.EE4BEG3 ),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2479_ (.I(FrameData[0]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2480_ (.I(FrameData[1]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2481_ (.I(FrameData[2]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2482_ (.I(FrameData[3]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2483_ (.I(FrameData[4]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2484_ (.I(FrameData[5]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2485_ (.I(FrameData[6]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2486_ (.I(FrameData[7]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2487_ (.I(FrameData[8]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2488_ (.I(FrameData[9]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2489_ (.I(FrameData[10]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2490_ (.I(FrameData[11]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2491_ (.I(FrameData[12]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2492_ (.I(FrameData[13]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2493_ (.I(FrameData[14]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2494_ (.I(FrameData[15]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2495_ (.I(FrameData[16]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2496_ (.I(FrameData[17]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2497_ (.I(FrameData[18]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2498_ (.I(FrameData[19]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2499_ (.I(FrameData[20]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2500_ (.I(FrameData[21]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2501_ (.I(FrameData[22]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2502_ (.I(FrameData[23]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2503_ (.I(FrameData[24]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2504_ (.I(FrameData[25]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2505_ (.I(FrameData[26]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2506_ (.I(FrameData[27]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2507_ (.I(FrameData[28]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2508_ (.I(FrameData[29]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2509_ (.I(FrameData[30]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2510_ (.I(FrameData[31]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2511_ (.I(FrameStrobe[0]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2512_ (.I(FrameStrobe[1]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2513_ (.I(FrameStrobe[2]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2514_ (.I(FrameStrobe[3]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2515_ (.I(FrameStrobe[4]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2516_ (.I(FrameStrobe[5]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2517_ (.I(FrameStrobe[6]),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2518_ (.I(FrameStrobe[7]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2519_ (.I(FrameStrobe[8]),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2520_ (.I(FrameStrobe[9]),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2521_ (.I(FrameStrobe[10]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2522_ (.I(FrameStrobe[11]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2523_ (.I(FrameStrobe[12]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2524_ (.I(FrameStrobe[13]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2525_ (.I(FrameStrobe[14]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2526_ (.I(FrameStrobe[15]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2527_ (.I(FrameStrobe[16]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2528_ (.I(FrameStrobe[17]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2529_ (.I(FrameStrobe[18]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2530_ (.I(FrameStrobe[19]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2531_ (.I(\Inst_LUT4AB_switch_matrix.N1BEG0 ),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2532_ (.I(\Inst_LUT4AB_switch_matrix.N1BEG1 ),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2533_ (.I(\Inst_LUT4AB_switch_matrix.N1BEG2 ),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2534_ (.I(\Inst_LUT4AB_switch_matrix.N1BEG3 ),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2535_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2536_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2537_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2538_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2539_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2540_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2541_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2542_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2543_ (.I(N2MID[0]),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2544_ (.I(N2MID[1]),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2545_ (.I(N2MID[2]),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2546_ (.I(N2MID[3]),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2547_ (.I(N2MID[4]),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2548_ (.I(N2MID[5]),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2549_ (.I(N2MID[6]),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2550_ (.I(N2MID[7]),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2551_ (.I(N4END[4]),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2552_ (.I(N4END[5]),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2553_ (.I(N4END[6]),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2554_ (.I(N4END[7]),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2555_ (.I(N4END[8]),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2556_ (.I(N4END[9]),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2557_ (.I(N4END[10]),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2558_ (.I(N4END[11]),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2559_ (.I(N4END[12]),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2560_ (.I(N4END[13]),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2561_ (.I(N4END[14]),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2562_ (.I(N4END[15]),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2563_ (.I(\Inst_LUT4AB_switch_matrix.N4BEG0 ),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2564_ (.I(\Inst_LUT4AB_switch_matrix.N4BEG1 ),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2565_ (.I(\Inst_LUT4AB_switch_matrix.N4BEG2 ),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2566_ (.I(\Inst_LUT4AB_switch_matrix.N4BEG3 ),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2567_ (.I(NN4END[4]),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2568_ (.I(NN4END[5]),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2569_ (.I(NN4END[6]),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2570_ (.I(NN4END[7]),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2571_ (.I(NN4END[8]),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2572_ (.I(NN4END[9]),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2573_ (.I(NN4END[10]),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2574_ (.I(NN4END[11]),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2575_ (.I(NN4END[12]),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2576_ (.I(NN4END[13]),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2577_ (.I(NN4END[14]),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2578_ (.I(NN4END[15]),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2579_ (.I(\Inst_LUT4AB_switch_matrix.NN4BEG0 ),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2580_ (.I(\Inst_LUT4AB_switch_matrix.NN4BEG1 ),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2581_ (.I(\Inst_LUT4AB_switch_matrix.NN4BEG2 ),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2582_ (.I(\Inst_LUT4AB_switch_matrix.NN4BEG3 ),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2583_ (.I(\Inst_LUT4AB_switch_matrix.S1BEG0 ),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2584_ (.I(\Inst_LUT4AB_switch_matrix.S1BEG1 ),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2585_ (.I(\Inst_LUT4AB_switch_matrix.S1BEG2 ),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2586_ (.I(\Inst_LUT4AB_switch_matrix.S1BEG3 ),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2587_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2588_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2589_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2590_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2591_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2592_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2593_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2594_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2595_ (.I(S2MID[0]),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2596_ (.I(S2MID[1]),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2597_ (.I(S2MID[2]),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2598_ (.I(S2MID[3]),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2599_ (.I(S2MID[4]),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2600_ (.I(S2MID[5]),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2601_ (.I(S2MID[6]),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2602_ (.I(S2MID[7]),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2603_ (.I(S4END[4]),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2604_ (.I(S4END[5]),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2605_ (.I(S4END[6]),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2606_ (.I(S4END[7]),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2607_ (.I(S4END[8]),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2608_ (.I(S4END[9]),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2609_ (.I(S4END[10]),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2610_ (.I(S4END[11]),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2611_ (.I(S4END[12]),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2612_ (.I(S4END[13]),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2613_ (.I(S4END[14]),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2614_ (.I(S4END[15]),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2615_ (.I(\Inst_LUT4AB_switch_matrix.S4BEG0 ),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2616_ (.I(\Inst_LUT4AB_switch_matrix.S4BEG1 ),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2617_ (.I(\Inst_LUT4AB_switch_matrix.S4BEG2 ),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2618_ (.I(\Inst_LUT4AB_switch_matrix.S4BEG3 ),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2619_ (.I(SS4END[4]),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2620_ (.I(SS4END[5]),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2621_ (.I(SS4END[6]),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2622_ (.I(SS4END[7]),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2623_ (.I(SS4END[8]),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2624_ (.I(SS4END[9]),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2625_ (.I(SS4END[10]),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2626_ (.I(SS4END[11]),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2627_ (.I(SS4END[12]),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2628_ (.I(SS4END[13]),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2629_ (.I(SS4END[14]),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2630_ (.I(SS4END[15]),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2631_ (.I(\Inst_LUT4AB_switch_matrix.SS4BEG0 ),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2632_ (.I(\Inst_LUT4AB_switch_matrix.SS4BEG1 ),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2633_ (.I(\Inst_LUT4AB_switch_matrix.SS4BEG2 ),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2634_ (.I(\Inst_LUT4AB_switch_matrix.SS4BEG3 ),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2635_ (.I(clknet_1_0__leaf_UserCLK),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2636_ (.I(\Inst_LUT4AB_switch_matrix.W1BEG0 ),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2637_ (.I(\Inst_LUT4AB_switch_matrix.W1BEG1 ),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2638_ (.I(\Inst_LUT4AB_switch_matrix.W1BEG2 ),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2639_ (.I(\Inst_LUT4AB_switch_matrix.W1BEG3 ),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2640_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2641_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2642_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2643_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2644_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2645_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2646_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2647_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG7 ),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2648_ (.I(W2MID[0]),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2649_ (.I(W2MID[1]),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2650_ (.I(W2MID[2]),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2651_ (.I(W2MID[3]),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2652_ (.I(W2MID[4]),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2653_ (.I(W2MID[5]),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2654_ (.I(W2MID[6]),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2655_ (.I(W2MID[7]),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2656_ (.I(W6END[2]),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2657_ (.I(W6END[3]),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2658_ (.I(W6END[4]),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2659_ (.I(W6END[5]),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2660_ (.I(W6END[6]),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2661_ (.I(W6END[7]),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2662_ (.I(W6END[8]),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2663_ (.I(W6END[9]),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2664_ (.I(W6END[10]),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2665_ (.I(W6END[11]),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2666_ (.I(\Inst_LUT4AB_switch_matrix.W6BEG0 ),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2667_ (.I(\Inst_LUT4AB_switch_matrix.W6BEG1 ),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2668_ (.I(WW4END[4]),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2669_ (.I(WW4END[5]),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2670_ (.I(WW4END[6]),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2671_ (.I(WW4END[7]),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2672_ (.I(WW4END[8]),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2673_ (.I(WW4END[9]),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2674_ (.I(WW4END[10]),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2675_ (.I(WW4END[11]),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2676_ (.I(WW4END[12]),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2677_ (.I(WW4END[13]),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2678_ (.I(WW4END[14]),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2679_ (.I(WW4END[15]),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2680_ (.I(\Inst_LUT4AB_switch_matrix.WW4BEG0 ),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2681_ (.I(\Inst_LUT4AB_switch_matrix.WW4BEG1 ),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2682_ (.I(\Inst_LUT4AB_switch_matrix.WW4BEG2 ),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2683_ (.I(\Inst_LUT4AB_switch_matrix.WW4BEG3 ),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_652 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output1 (.I(net1),
    .Z(Co));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output2 (.I(net2),
    .Z(E1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output3 (.I(net3),
    .Z(E1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output4 (.I(net4),
    .Z(E1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output5 (.I(net5),
    .Z(E1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output6 (.I(net6),
    .Z(E2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output7 (.I(net7),
    .Z(E2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output8 (.I(net8),
    .Z(E2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output9 (.I(net9),
    .Z(E2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output10 (.I(net10),
    .Z(E2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output11 (.I(net11),
    .Z(E2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output12 (.I(net12),
    .Z(E2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output13 (.I(net13),
    .Z(E2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output14 (.I(net14),
    .Z(E2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output15 (.I(net15),
    .Z(E2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output16 (.I(net16),
    .Z(E2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output17 (.I(net17),
    .Z(E2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output18 (.I(net18),
    .Z(E2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output19 (.I(net19),
    .Z(E2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output20 (.I(net20),
    .Z(E2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output21 (.I(net21),
    .Z(E2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output22 (.I(net22),
    .Z(E6BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output23 (.I(net23),
    .Z(E6BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output24 (.I(net24),
    .Z(E6BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output25 (.I(net25),
    .Z(E6BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output26 (.I(net26),
    .Z(E6BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output27 (.I(net27),
    .Z(E6BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output28 (.I(net28),
    .Z(E6BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output29 (.I(net29),
    .Z(E6BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output30 (.I(net30),
    .Z(E6BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output31 (.I(net31),
    .Z(E6BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output32 (.I(net32),
    .Z(E6BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output33 (.I(net33),
    .Z(E6BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output34 (.I(net34),
    .Z(EE4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output35 (.I(net35),
    .Z(EE4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output36 (.I(net36),
    .Z(EE4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output37 (.I(net37),
    .Z(EE4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output38 (.I(net38),
    .Z(EE4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output39 (.I(net39),
    .Z(EE4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output40 (.I(net40),
    .Z(EE4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output41 (.I(net41),
    .Z(EE4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output42 (.I(net42),
    .Z(EE4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output43 (.I(net43),
    .Z(EE4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output44 (.I(net44),
    .Z(EE4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output45 (.I(net45),
    .Z(EE4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output46 (.I(net46),
    .Z(EE4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output47 (.I(net47),
    .Z(EE4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output48 (.I(net48),
    .Z(EE4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output49 (.I(net49),
    .Z(EE4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output50 (.I(net50),
    .Z(FrameData_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output51 (.I(net51),
    .Z(FrameData_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output52 (.I(net52),
    .Z(FrameData_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output53 (.I(net53),
    .Z(FrameData_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output54 (.I(net54),
    .Z(FrameData_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output55 (.I(net55),
    .Z(FrameData_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output56 (.I(net56),
    .Z(FrameData_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output57 (.I(net57),
    .Z(FrameData_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output58 (.I(net58),
    .Z(FrameData_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output59 (.I(net59),
    .Z(FrameData_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output60 (.I(net60),
    .Z(FrameData_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output61 (.I(net61),
    .Z(FrameData_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output62 (.I(net62),
    .Z(FrameData_O[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output63 (.I(net63),
    .Z(FrameData_O[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output64 (.I(net64),
    .Z(FrameData_O[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output65 (.I(net65),
    .Z(FrameData_O[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output66 (.I(net66),
    .Z(FrameData_O[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output67 (.I(net67),
    .Z(FrameData_O[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output68 (.I(net68),
    .Z(FrameData_O[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output69 (.I(net69),
    .Z(FrameData_O[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output70 (.I(net70),
    .Z(FrameData_O[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output71 (.I(net71),
    .Z(FrameData_O[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output72 (.I(net72),
    .Z(FrameData_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output73 (.I(net73),
    .Z(FrameData_O[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output74 (.I(net74),
    .Z(FrameData_O[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output75 (.I(net75),
    .Z(FrameData_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output76 (.I(net76),
    .Z(FrameData_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output77 (.I(net77),
    .Z(FrameData_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output78 (.I(net78),
    .Z(FrameData_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output79 (.I(net79),
    .Z(FrameData_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output80 (.I(net80),
    .Z(FrameData_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output81 (.I(net81),
    .Z(FrameData_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output82 (.I(net82),
    .Z(FrameStrobe_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output83 (.I(net83),
    .Z(FrameStrobe_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output84 (.I(net84),
    .Z(FrameStrobe_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output85 (.I(net85),
    .Z(FrameStrobe_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output86 (.I(net86),
    .Z(FrameStrobe_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output87 (.I(net87),
    .Z(FrameStrobe_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output88 (.I(net88),
    .Z(FrameStrobe_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output89 (.I(net89),
    .Z(FrameStrobe_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output90 (.I(net90),
    .Z(FrameStrobe_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output91 (.I(net91),
    .Z(FrameStrobe_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output92 (.I(net92),
    .Z(FrameStrobe_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output93 (.I(net93),
    .Z(FrameStrobe_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output94 (.I(net94),
    .Z(FrameStrobe_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output95 (.I(net95),
    .Z(FrameStrobe_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output96 (.I(net96),
    .Z(FrameStrobe_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output97 (.I(net97),
    .Z(FrameStrobe_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output98 (.I(net98),
    .Z(FrameStrobe_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output99 (.I(net99),
    .Z(FrameStrobe_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output100 (.I(net100),
    .Z(FrameStrobe_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output101 (.I(net101),
    .Z(FrameStrobe_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output102 (.I(net102),
    .Z(N1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output103 (.I(net103),
    .Z(N1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output104 (.I(net104),
    .Z(N1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output105 (.I(net105),
    .Z(N1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output106 (.I(net106),
    .Z(N2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output107 (.I(net107),
    .Z(N2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output108 (.I(net108),
    .Z(N2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output109 (.I(net109),
    .Z(N2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output110 (.I(net110),
    .Z(N2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output111 (.I(net111),
    .Z(N2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output112 (.I(net112),
    .Z(N2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output113 (.I(net113),
    .Z(N2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output114 (.I(net114),
    .Z(N2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output115 (.I(net115),
    .Z(N2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output116 (.I(net116),
    .Z(N2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output117 (.I(net117),
    .Z(N2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output118 (.I(net118),
    .Z(N2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output119 (.I(net119),
    .Z(N2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output120 (.I(net120),
    .Z(N2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output121 (.I(net121),
    .Z(N2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output122 (.I(net122),
    .Z(N4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output123 (.I(net123),
    .Z(N4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output124 (.I(net124),
    .Z(N4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output125 (.I(net125),
    .Z(N4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output126 (.I(net126),
    .Z(N4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output127 (.I(net127),
    .Z(N4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output128 (.I(net128),
    .Z(N4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output129 (.I(net129),
    .Z(N4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output130 (.I(net130),
    .Z(N4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output131 (.I(net131),
    .Z(N4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output132 (.I(net132),
    .Z(N4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output133 (.I(net133),
    .Z(N4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output134 (.I(net134),
    .Z(N4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output135 (.I(net135),
    .Z(N4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output136 (.I(net136),
    .Z(N4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output137 (.I(net137),
    .Z(N4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output138 (.I(net138),
    .Z(NN4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output139 (.I(net139),
    .Z(NN4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output140 (.I(net140),
    .Z(NN4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output141 (.I(net141),
    .Z(NN4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output142 (.I(net142),
    .Z(NN4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output143 (.I(net143),
    .Z(NN4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output144 (.I(net144),
    .Z(NN4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output145 (.I(net145),
    .Z(NN4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output146 (.I(net146),
    .Z(NN4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output147 (.I(net147),
    .Z(NN4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output148 (.I(net148),
    .Z(NN4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output149 (.I(net149),
    .Z(NN4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output150 (.I(net150),
    .Z(NN4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output151 (.I(net151),
    .Z(NN4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output152 (.I(net152),
    .Z(NN4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output153 (.I(net153),
    .Z(NN4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output154 (.I(net154),
    .Z(S1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output155 (.I(net155),
    .Z(S1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output156 (.I(net156),
    .Z(S1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output157 (.I(net157),
    .Z(S1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output158 (.I(net158),
    .Z(S2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output159 (.I(net159),
    .Z(S2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output160 (.I(net160),
    .Z(S2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output161 (.I(net161),
    .Z(S2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output162 (.I(net162),
    .Z(S2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output163 (.I(net163),
    .Z(S2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output164 (.I(net164),
    .Z(S2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output165 (.I(net165),
    .Z(S2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output166 (.I(net166),
    .Z(S2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output167 (.I(net167),
    .Z(S2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output168 (.I(net168),
    .Z(S2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output169 (.I(net169),
    .Z(S2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output170 (.I(net170),
    .Z(S2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output171 (.I(net171),
    .Z(S2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output172 (.I(net172),
    .Z(S2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output173 (.I(net173),
    .Z(S2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output174 (.I(net174),
    .Z(S4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output175 (.I(net175),
    .Z(S4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output176 (.I(net176),
    .Z(S4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output177 (.I(net177),
    .Z(S4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output178 (.I(net178),
    .Z(S4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output179 (.I(net179),
    .Z(S4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output180 (.I(net180),
    .Z(S4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output181 (.I(net181),
    .Z(S4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output182 (.I(net182),
    .Z(S4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output183 (.I(net183),
    .Z(S4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output184 (.I(net184),
    .Z(S4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output185 (.I(net185),
    .Z(S4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output186 (.I(net186),
    .Z(S4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output187 (.I(net187),
    .Z(S4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output188 (.I(net188),
    .Z(S4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output189 (.I(net189),
    .Z(S4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output190 (.I(net190),
    .Z(SS4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output191 (.I(net191),
    .Z(SS4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output192 (.I(net192),
    .Z(SS4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output193 (.I(net193),
    .Z(SS4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output194 (.I(net194),
    .Z(SS4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output195 (.I(net195),
    .Z(SS4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output196 (.I(net196),
    .Z(SS4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output197 (.I(net197),
    .Z(SS4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output198 (.I(net198),
    .Z(SS4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output199 (.I(net199),
    .Z(SS4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output200 (.I(net200),
    .Z(SS4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output201 (.I(net201),
    .Z(SS4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output202 (.I(net202),
    .Z(SS4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output203 (.I(net203),
    .Z(SS4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output204 (.I(net204),
    .Z(SS4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output205 (.I(net205),
    .Z(SS4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output206 (.I(net206),
    .Z(UserCLKo));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output207 (.I(net207),
    .Z(W1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output208 (.I(net208),
    .Z(W1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output209 (.I(net209),
    .Z(W1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output210 (.I(net210),
    .Z(W1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output211 (.I(net211),
    .Z(W2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output212 (.I(net212),
    .Z(W2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output213 (.I(net213),
    .Z(W2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output214 (.I(net214),
    .Z(W2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output215 (.I(net215),
    .Z(W2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output216 (.I(net216),
    .Z(W2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output217 (.I(net217),
    .Z(W2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output218 (.I(net218),
    .Z(W2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output219 (.I(net219),
    .Z(W2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output220 (.I(net220),
    .Z(W2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output221 (.I(net221),
    .Z(W2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output222 (.I(net222),
    .Z(W2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output223 (.I(net223),
    .Z(W2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output224 (.I(net224),
    .Z(W2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output225 (.I(net225),
    .Z(W2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output226 (.I(net226),
    .Z(W2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output227 (.I(net227),
    .Z(W6BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output228 (.I(net228),
    .Z(W6BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output229 (.I(net229),
    .Z(W6BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output230 (.I(net230),
    .Z(W6BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output231 (.I(net231),
    .Z(W6BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output232 (.I(net232),
    .Z(W6BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output233 (.I(net233),
    .Z(W6BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output234 (.I(net234),
    .Z(W6BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output235 (.I(net235),
    .Z(W6BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output236 (.I(net236),
    .Z(W6BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output237 (.I(net237),
    .Z(W6BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output238 (.I(net238),
    .Z(W6BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output239 (.I(net239),
    .Z(WW4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output240 (.I(net240),
    .Z(WW4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output241 (.I(net241),
    .Z(WW4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output242 (.I(net242),
    .Z(WW4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output243 (.I(net243),
    .Z(WW4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output244 (.I(net244),
    .Z(WW4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output245 (.I(net245),
    .Z(WW4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output246 (.I(net246),
    .Z(WW4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output247 (.I(net247),
    .Z(WW4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output248 (.I(net248),
    .Z(WW4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output249 (.I(net249),
    .Z(WW4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output250 (.I(net250),
    .Z(WW4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output251 (.I(net251),
    .Z(WW4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output252 (.I(net252),
    .Z(WW4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output253 (.I(net253),
    .Z(WW4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output254 (.I(net254),
    .Z(WW4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_regs_0_UserCLK (.I(UserCLK),
    .Z(UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_UserCLK (.I(UserCLK),
    .Z(clknet_0_UserCLK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_UserCLK (.I(clknet_0_UserCLK),
    .Z(clknet_1_0__leaf_UserCLK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_UserCLK_regs (.I(UserCLK_regs),
    .Z(clknet_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_1_0__leaf_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_1_1__leaf_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(E6END[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(E6END[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_3 (.I(E6END[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_4 (.I(EE4END[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_5 (.I(EE4END[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_6 (.I(EE4END[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_7 (.I(EE4END[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_8 (.I(EE4END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_9 (.I(EE4END[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_10 (.I(\Inst_LUT4AB_switch_matrix.JW2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_11 (.I(N4END[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_12 (.I(N4END[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_13 (.I(N4END[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_14 (.I(N4END[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_15 (.I(N4END[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_16 (.I(N4END[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_17 (.I(N4END[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_18 (.I(N4END[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_19 (.I(N4END[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_20 (.I(N4END[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_21 (.I(N4END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_22 (.I(N4END[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_23 (.I(NN4END[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_24 (.I(NN4END[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_25 (.I(NN4END[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_26 (.I(NN4END[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_27 (.I(NN4END[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_28 (.I(NN4END[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_29 (.I(NN4END[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_30 (.I(NN4END[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_31 (.I(NN4END[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_32 (.I(NN4END[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_33 (.I(NN4END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_34 (.I(NN4END[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_35 (.I(SS4END[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_36 (.I(SS4END[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_37 (.I(SS4END[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_38 (.I(SS4END[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_39 (.I(SS4END[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_40 (.I(SS4END[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_41 (.I(SS4END[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_42 (.I(SS4END[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_43 (.I(SS4END[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_44 (.I(SS4END[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_45 (.I(SS4END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_46 (.I(SS4END[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_47 (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_48 (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_49 (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_50 (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_51 (.I(B));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_52 (.I(EE4END[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_53 (.I(N4END[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_54 (.I(SS4END[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_55 (.I(W2MID[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_56 (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_57 (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_58 (.I(W6END[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_59 (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_60 (.I(N4END[13]));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_478 ();
endmodule
