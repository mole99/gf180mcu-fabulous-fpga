magic
tech gf180mcuD
magscale 1 5
timestamp 1764324520
<< metal1 >>
rect 336 6677 15512 6694
rect 336 6651 2233 6677
rect 2259 6651 2285 6677
rect 2311 6651 2337 6677
rect 2363 6651 12233 6677
rect 12259 6651 12285 6677
rect 12311 6651 12337 6677
rect 12363 6651 15512 6677
rect 336 6634 15512 6651
rect 1079 6593 1105 6599
rect 1079 6561 1105 6567
rect 1863 6593 1889 6599
rect 1863 6561 1889 6567
rect 2983 6593 3009 6599
rect 2983 6561 3009 6567
rect 3767 6593 3793 6599
rect 3767 6561 3793 6567
rect 4887 6593 4913 6599
rect 4887 6561 4913 6567
rect 5671 6593 5697 6599
rect 5671 6561 5697 6567
rect 6567 6593 6593 6599
rect 6567 6561 6593 6567
rect 7015 6593 7041 6599
rect 7015 6561 7041 6567
rect 7855 6593 7881 6599
rect 7855 6561 7881 6567
rect 9479 6593 9505 6599
rect 9479 6561 9505 6567
rect 11271 6593 11297 6599
rect 11271 6561 11297 6567
rect 12223 6593 12249 6599
rect 12223 6561 12249 6567
rect 13007 6593 13033 6599
rect 13007 6561 13033 6567
rect 14127 6593 14153 6599
rect 14127 6561 14153 6567
rect 14911 6593 14937 6599
rect 14911 6561 14937 6567
rect 7575 6537 7601 6543
rect 3257 6511 3263 6537
rect 3289 6511 3295 6537
rect 7575 6505 7601 6511
rect 1353 6455 1359 6481
rect 1385 6455 1391 6481
rect 2137 6455 2143 6481
rect 2169 6455 2175 6481
rect 3929 6455 3935 6481
rect 3961 6455 3967 6481
rect 5161 6455 5167 6481
rect 5193 6455 5199 6481
rect 5945 6455 5951 6481
rect 5977 6455 5983 6481
rect 6729 6455 6735 6481
rect 6761 6455 6767 6481
rect 9081 6455 9087 6481
rect 9113 6455 9119 6481
rect 10817 6455 10823 6481
rect 10849 6455 10855 6481
rect 10985 6455 10991 6481
rect 11017 6455 11023 6481
rect 11937 6455 11943 6481
rect 11969 6455 11975 6481
rect 12833 6455 12839 6481
rect 12865 6455 12871 6481
rect 13953 6455 13959 6481
rect 13985 6455 13991 6481
rect 14625 6455 14631 6481
rect 14657 6455 14663 6481
rect 6287 6425 6313 6431
rect 6287 6393 6313 6399
rect 8863 6425 8889 6431
rect 9697 6399 9703 6425
rect 9729 6399 9735 6425
rect 10481 6399 10487 6425
rect 10513 6399 10519 6425
rect 8863 6393 8889 6399
rect 336 6285 15512 6302
rect 336 6259 1903 6285
rect 1929 6259 1955 6285
rect 1981 6259 2007 6285
rect 2033 6259 11903 6285
rect 11929 6259 11955 6285
rect 11981 6259 12007 6285
rect 12033 6259 15512 6285
rect 336 6242 15512 6259
rect 3655 6201 3681 6207
rect 3655 6169 3681 6175
rect 5055 6201 5081 6207
rect 5055 6169 5081 6175
rect 6007 6201 6033 6207
rect 6007 6169 6033 6175
rect 6735 6201 6761 6207
rect 6735 6169 6761 6175
rect 11383 6201 11409 6207
rect 11383 6169 11409 6175
rect 11999 6201 12025 6207
rect 11999 6169 12025 6175
rect 12951 6201 12977 6207
rect 12951 6169 12977 6175
rect 14519 6201 14545 6207
rect 14519 6169 14545 6175
rect 1919 6145 1945 6151
rect 10039 6145 10065 6151
rect 2753 6119 2759 6145
rect 2785 6119 2791 6145
rect 4153 6119 4159 6145
rect 4185 6119 4191 6145
rect 9249 6119 9255 6145
rect 9281 6119 9287 6145
rect 10593 6119 10599 6145
rect 10625 6119 10631 6145
rect 1919 6113 1945 6119
rect 10039 6113 10065 6119
rect 7687 6089 7713 6095
rect 3145 6063 3151 6089
rect 3177 6063 3183 6089
rect 7233 6063 7239 6089
rect 7265 6063 7271 6089
rect 7687 6057 7713 6063
rect 8135 6089 8161 6095
rect 8135 6057 8161 6063
rect 8583 6089 8609 6095
rect 9479 6089 9505 6095
rect 8969 6063 8975 6089
rect 9001 6063 9007 6089
rect 8583 6057 8609 6063
rect 9479 6057 9505 6063
rect 9759 6089 9785 6095
rect 14289 6063 14295 6089
rect 14321 6063 14327 6089
rect 9759 6057 9785 6063
rect 7407 6033 7433 6039
rect 2193 6007 2199 6033
rect 2225 6007 2231 6033
rect 4545 6007 4551 6033
rect 4577 6007 4583 6033
rect 5329 6007 5335 6033
rect 5361 6007 5367 6033
rect 5497 6007 5503 6033
rect 5529 6007 5535 6033
rect 7407 6001 7433 6007
rect 7855 6033 7881 6039
rect 7855 6001 7881 6007
rect 8303 6033 8329 6039
rect 8303 6001 8329 6007
rect 8751 6033 8777 6039
rect 13735 6033 13761 6039
rect 10929 6007 10935 6033
rect 10961 6007 10967 6033
rect 11097 6007 11103 6033
rect 11129 6007 11135 6033
rect 12497 6007 12503 6033
rect 12529 6007 12535 6033
rect 12665 6007 12671 6033
rect 12697 6007 12703 6033
rect 8751 6001 8777 6007
rect 13735 6001 13761 6007
rect 15303 6033 15329 6039
rect 15303 6001 15329 6007
rect 2983 5977 3009 5983
rect 2983 5945 3009 5951
rect 13455 5977 13481 5983
rect 13455 5945 13481 5951
rect 15023 5977 15049 5983
rect 15023 5945 15049 5951
rect 336 5893 15512 5910
rect 336 5867 2233 5893
rect 2259 5867 2285 5893
rect 2311 5867 2337 5893
rect 2363 5867 12233 5893
rect 12259 5867 12285 5893
rect 12311 5867 12337 5893
rect 12363 5867 15512 5893
rect 336 5850 15512 5867
rect 2311 5809 2337 5815
rect 2311 5777 2337 5783
rect 3879 5809 3905 5815
rect 3879 5777 3905 5783
rect 4775 5809 4801 5815
rect 4775 5777 4801 5783
rect 11607 5809 11633 5815
rect 11607 5777 11633 5783
rect 14127 5809 14153 5815
rect 14127 5777 14153 5783
rect 1527 5753 1553 5759
rect 1527 5721 1553 5727
rect 4495 5753 4521 5759
rect 5161 5727 5167 5753
rect 5193 5727 5199 5753
rect 7121 5727 7127 5753
rect 7153 5727 7159 5753
rect 4495 5721 4521 5727
rect 7631 5697 7657 5703
rect 1745 5671 1751 5697
rect 1777 5671 1783 5697
rect 2585 5671 2591 5697
rect 2617 5671 2623 5697
rect 2977 5671 2983 5697
rect 3009 5671 3015 5697
rect 3257 5671 3263 5697
rect 3289 5671 3295 5697
rect 4153 5671 4159 5697
rect 4185 5671 4191 5697
rect 5553 5671 5559 5697
rect 5585 5671 5591 5697
rect 5721 5671 5727 5697
rect 5753 5671 5759 5697
rect 7631 5665 7657 5671
rect 9759 5697 9785 5703
rect 10711 5697 10737 5703
rect 10257 5671 10263 5697
rect 10289 5671 10295 5697
rect 11321 5671 11327 5697
rect 11353 5671 11359 5697
rect 12273 5671 12279 5697
rect 12305 5671 12311 5697
rect 13057 5671 13063 5697
rect 13089 5671 13095 5697
rect 13841 5671 13847 5697
rect 13873 5671 13879 5697
rect 14681 5671 14687 5697
rect 14713 5671 14719 5697
rect 9759 5665 9785 5671
rect 10711 5665 10737 5671
rect 6623 5641 6649 5647
rect 6057 5615 6063 5641
rect 6089 5615 6095 5641
rect 6623 5609 6649 5615
rect 7911 5641 7937 5647
rect 7911 5609 7937 5615
rect 10039 5641 10065 5647
rect 10039 5609 10065 5615
rect 10487 5641 10513 5647
rect 12559 5641 12585 5647
rect 10929 5615 10935 5641
rect 10961 5615 10967 5641
rect 10487 5609 10513 5615
rect 12559 5609 12585 5615
rect 13567 5641 13593 5647
rect 13567 5609 13593 5615
rect 15191 5585 15217 5591
rect 15191 5553 15217 5559
rect 336 5501 15512 5518
rect 336 5475 1903 5501
rect 1929 5475 1955 5501
rect 1981 5475 2007 5501
rect 2033 5475 11903 5501
rect 11929 5475 11955 5501
rect 11981 5475 12007 5501
rect 12033 5475 15512 5501
rect 336 5458 15512 5475
rect 1919 5417 1945 5423
rect 1919 5385 1945 5391
rect 3487 5417 3513 5423
rect 3487 5385 3513 5391
rect 4271 5417 4297 5423
rect 4271 5385 4297 5391
rect 5055 5417 5081 5423
rect 5055 5385 5081 5391
rect 11831 5417 11857 5423
rect 11831 5385 11857 5391
rect 12615 5417 12641 5423
rect 12615 5385 12641 5391
rect 7183 5361 7209 5367
rect 8807 5361 8833 5367
rect 11383 5361 11409 5367
rect 5777 5335 5783 5361
rect 5809 5335 5815 5361
rect 6561 5335 6567 5361
rect 6593 5335 6599 5361
rect 8353 5335 8359 5361
rect 8385 5335 8391 5361
rect 9809 5335 9815 5361
rect 9841 5335 9847 5361
rect 13505 5335 13511 5361
rect 13537 5335 13543 5361
rect 14457 5335 14463 5361
rect 14489 5335 14495 5361
rect 7183 5329 7209 5335
rect 8807 5329 8833 5335
rect 11383 5329 11409 5335
rect 2703 5305 2729 5311
rect 2081 5279 2087 5305
rect 2113 5279 2119 5305
rect 2703 5273 2729 5279
rect 2983 5305 3009 5311
rect 7463 5305 7489 5311
rect 3761 5279 3767 5305
rect 3793 5279 3799 5305
rect 4545 5279 4551 5305
rect 4577 5279 4583 5305
rect 5329 5279 5335 5305
rect 5361 5279 5367 5305
rect 7009 5279 7015 5305
rect 7041 5279 7047 5305
rect 2983 5273 3009 5279
rect 7463 5273 7489 5279
rect 9087 5305 9113 5311
rect 9087 5273 9113 5279
rect 9535 5305 9561 5311
rect 11103 5305 11129 5311
rect 9977 5279 9983 5305
rect 10009 5279 10015 5305
rect 11545 5279 11551 5305
rect 11577 5279 11583 5305
rect 14289 5279 14295 5305
rect 14321 5279 14327 5305
rect 9535 5273 9561 5279
rect 11103 5273 11129 5279
rect 7967 5249 7993 5255
rect 6113 5223 6119 5249
rect 6145 5223 6151 5249
rect 7967 5217 7993 5223
rect 9255 5249 9281 5255
rect 10655 5249 10681 5255
rect 10481 5223 10487 5249
rect 10513 5223 10519 5249
rect 9255 5217 9281 5223
rect 10655 5217 10681 5223
rect 10935 5249 10961 5255
rect 12329 5223 12335 5249
rect 12361 5223 12367 5249
rect 13113 5223 13119 5249
rect 13145 5223 13151 5249
rect 14681 5223 14687 5249
rect 14713 5223 14719 5249
rect 15073 5223 15079 5249
rect 15105 5223 15111 5249
rect 10935 5217 10961 5223
rect 7687 5193 7713 5199
rect 7687 5161 7713 5167
rect 8135 5193 8161 5199
rect 8135 5161 8161 5167
rect 10319 5193 10345 5199
rect 10319 5161 10345 5167
rect 336 5109 15512 5126
rect 336 5083 2233 5109
rect 2259 5083 2285 5109
rect 2311 5083 2337 5109
rect 2363 5083 12233 5109
rect 12259 5083 12285 5109
rect 12311 5083 12337 5109
rect 12363 5083 15512 5109
rect 336 5066 15512 5083
rect 3095 5025 3121 5031
rect 3095 4993 3121 4999
rect 3879 5025 3905 5031
rect 3879 4993 3905 4999
rect 7183 5025 7209 5031
rect 7183 4993 7209 4999
rect 10543 5025 10569 5031
rect 10543 4993 10569 4999
rect 11551 5025 11577 5031
rect 11551 4993 11577 4999
rect 12559 5025 12585 5031
rect 12559 4993 12585 4999
rect 10823 4969 10849 4975
rect 4937 4943 4943 4969
rect 4969 4943 4975 4969
rect 5329 4943 5335 4969
rect 5361 4943 5367 4969
rect 14289 4943 14295 4969
rect 14321 4943 14327 4969
rect 10823 4937 10849 4943
rect 11383 4913 11409 4919
rect 2025 4887 2031 4913
rect 2057 4887 2063 4913
rect 3313 4887 3319 4913
rect 3345 4887 3351 4913
rect 4153 4887 4159 4913
rect 4185 4887 4191 4913
rect 6113 4887 6119 4913
rect 6145 4887 6151 4913
rect 6673 4887 6679 4913
rect 6705 4887 6711 4913
rect 12273 4887 12279 4913
rect 12305 4887 12311 4913
rect 13561 4887 13567 4913
rect 13593 4887 13599 4913
rect 14009 4887 14015 4913
rect 14041 4887 14047 4913
rect 14737 4887 14743 4913
rect 14769 4887 14775 4913
rect 11383 4881 11409 4887
rect 2479 4857 2505 4863
rect 6903 4857 6929 4863
rect 11831 4857 11857 4863
rect 6505 4831 6511 4857
rect 6537 4831 6543 4857
rect 11153 4831 11159 4857
rect 11185 4831 11191 4857
rect 2479 4825 2505 4831
rect 6903 4825 6929 4831
rect 11831 4825 11857 4831
rect 13175 4857 13201 4863
rect 13175 4825 13201 4831
rect 5615 4801 5641 4807
rect 5615 4769 5641 4775
rect 15191 4801 15217 4807
rect 15191 4769 15217 4775
rect 336 4717 15512 4734
rect 336 4691 1903 4717
rect 1929 4691 1955 4717
rect 1981 4691 2007 4717
rect 2033 4691 11903 4717
rect 11929 4691 11955 4717
rect 11981 4691 12007 4717
rect 12033 4691 15512 4717
rect 336 4674 15512 4691
rect 3711 4633 3737 4639
rect 3711 4601 3737 4607
rect 5223 4633 5249 4639
rect 5223 4601 5249 4607
rect 12671 4633 12697 4639
rect 12671 4601 12697 4607
rect 13455 4633 13481 4639
rect 13455 4601 13481 4607
rect 7855 4577 7881 4583
rect 14519 4577 14545 4583
rect 3033 4551 3039 4577
rect 3065 4551 3071 4577
rect 4321 4551 4327 4577
rect 4353 4551 4359 4577
rect 11713 4551 11719 4577
rect 11745 4551 11751 4577
rect 7855 4545 7881 4551
rect 14519 4545 14545 4551
rect 2143 4521 2169 4527
rect 6007 4521 6033 4527
rect 12223 4521 12249 4527
rect 4769 4495 4775 4521
rect 4801 4495 4807 4521
rect 11993 4495 11999 4521
rect 12025 4495 12031 4521
rect 13057 4495 13063 4521
rect 13089 4495 13095 4521
rect 14289 4495 14295 4521
rect 14321 4495 14327 4521
rect 14681 4495 14687 4521
rect 14713 4495 14719 4521
rect 2143 4489 2169 4495
rect 6007 4489 6033 4495
rect 12223 4489 12249 4495
rect 1863 4465 1889 4471
rect 5727 4465 5753 4471
rect 2585 4439 2591 4465
rect 2617 4439 2623 4465
rect 3985 4439 3991 4465
rect 4017 4439 4023 4465
rect 4937 4439 4943 4465
rect 4969 4439 4975 4465
rect 1863 4433 1889 4439
rect 5727 4433 5753 4439
rect 8471 4465 8497 4471
rect 13953 4439 13959 4465
rect 13985 4439 13991 4465
rect 15073 4439 15079 4465
rect 15105 4439 15111 4465
rect 8471 4433 8497 4439
rect 7575 4409 7601 4415
rect 7575 4377 7601 4383
rect 8191 4409 8217 4415
rect 8191 4377 8217 4383
rect 11495 4409 11521 4415
rect 11495 4377 11521 4383
rect 336 4325 15512 4342
rect 336 4299 2233 4325
rect 2259 4299 2285 4325
rect 2311 4299 2337 4325
rect 2363 4299 12233 4325
rect 12259 4299 12285 4325
rect 12311 4299 12337 4325
rect 12363 4299 15512 4325
rect 336 4282 15512 4299
rect 5783 4241 5809 4247
rect 5783 4209 5809 4215
rect 6231 4241 6257 4247
rect 6231 4209 6257 4215
rect 2311 4185 2337 4191
rect 4439 4185 4465 4191
rect 4153 4159 4159 4185
rect 4185 4159 4191 4185
rect 2311 4153 2337 4159
rect 4439 4153 4465 4159
rect 5279 4185 5305 4191
rect 5279 4153 5305 4159
rect 5503 4185 5529 4191
rect 12329 4159 12335 4185
rect 12361 4159 12367 4185
rect 12721 4159 12727 4185
rect 12753 4159 12759 4185
rect 5503 4153 5529 4159
rect 2591 4129 2617 4135
rect 4719 4129 4745 4135
rect 3369 4103 3375 4129
rect 3401 4103 3407 4129
rect 7849 4103 7855 4129
rect 7881 4103 7887 4129
rect 13225 4103 13231 4129
rect 13257 4103 13263 4129
rect 13897 4103 13903 4129
rect 13929 4103 13935 4129
rect 14681 4103 14687 4129
rect 14713 4103 14719 4129
rect 2591 4097 2617 4103
rect 4719 4097 4745 4103
rect 3655 4073 3681 4079
rect 5951 4073 5977 4079
rect 13623 4073 13649 4079
rect 2921 4047 2927 4073
rect 2953 4047 2959 4073
rect 5049 4047 5055 4073
rect 5081 4047 5087 4073
rect 8017 4047 8023 4073
rect 8049 4047 8055 4073
rect 3655 4041 3681 4047
rect 5951 4041 5977 4047
rect 13623 4041 13649 4047
rect 14407 4073 14433 4079
rect 14407 4041 14433 4047
rect 15191 4017 15217 4023
rect 15191 3985 15217 3991
rect 336 3933 15512 3950
rect 336 3907 1903 3933
rect 1929 3907 1955 3933
rect 1981 3907 2007 3933
rect 2033 3907 11903 3933
rect 11929 3907 11955 3933
rect 11981 3907 12007 3933
rect 12033 3907 15512 3933
rect 336 3890 15512 3907
rect 12895 3849 12921 3855
rect 12895 3817 12921 3823
rect 13847 3849 13873 3855
rect 13847 3817 13873 3823
rect 3431 3793 3457 3799
rect 5167 3793 5193 3799
rect 4097 3767 4103 3793
rect 4129 3767 4135 3793
rect 3431 3761 3457 3767
rect 5167 3761 5193 3767
rect 8079 3793 8105 3799
rect 15129 3767 15135 3793
rect 15161 3767 15167 3793
rect 8079 3761 8105 3767
rect 7799 3737 7825 3743
rect 5385 3711 5391 3737
rect 5417 3711 5423 3737
rect 13169 3711 13175 3737
rect 13201 3711 13207 3737
rect 7799 3705 7825 3711
rect 3711 3681 3737 3687
rect 3711 3649 3737 3655
rect 7631 3681 7657 3687
rect 13337 3655 13343 3681
rect 13369 3655 13375 3681
rect 14681 3655 14687 3681
rect 14713 3655 14719 3681
rect 7631 3649 7657 3655
rect 4327 3625 4353 3631
rect 4327 3593 4353 3599
rect 7351 3625 7377 3631
rect 7351 3593 7377 3599
rect 336 3541 15512 3558
rect 336 3515 2233 3541
rect 2259 3515 2285 3541
rect 2311 3515 2337 3541
rect 2363 3515 12233 3541
rect 12259 3515 12285 3541
rect 12311 3515 12337 3541
rect 12363 3515 15512 3541
rect 336 3498 15512 3515
rect 13113 3375 13119 3401
rect 13145 3375 13151 3401
rect 3879 3345 3905 3351
rect 7183 3345 7209 3351
rect 4097 3319 4103 3345
rect 4129 3319 4135 3345
rect 8409 3319 8415 3345
rect 8441 3319 8447 3345
rect 13897 3319 13903 3345
rect 13929 3319 13935 3345
rect 14681 3319 14687 3345
rect 14713 3319 14719 3345
rect 3879 3313 3905 3319
rect 7183 3313 7209 3319
rect 7463 3289 7489 3295
rect 7463 3257 7489 3263
rect 8639 3289 8665 3295
rect 8639 3257 8665 3263
rect 13623 3289 13649 3295
rect 13623 3257 13649 3263
rect 15191 3289 15217 3295
rect 15191 3257 15217 3263
rect 14407 3233 14433 3239
rect 14407 3201 14433 3207
rect 336 3149 15512 3166
rect 336 3123 1903 3149
rect 1929 3123 1955 3149
rect 1981 3123 2007 3149
rect 2033 3123 11903 3149
rect 11929 3123 11955 3149
rect 11981 3123 12007 3149
rect 12033 3123 15512 3149
rect 336 3106 15512 3123
rect 7519 3009 7545 3015
rect 15129 2983 15135 3009
rect 15161 2983 15167 3009
rect 7519 2977 7545 2983
rect 7239 2953 7265 2959
rect 7239 2921 7265 2927
rect 14681 2871 14687 2897
rect 14713 2871 14719 2897
rect 336 2757 15512 2774
rect 336 2731 2233 2757
rect 2259 2731 2285 2757
rect 2311 2731 2337 2757
rect 2363 2731 12233 2757
rect 12259 2731 12285 2757
rect 12311 2731 12337 2757
rect 12363 2731 15512 2757
rect 336 2714 15512 2731
rect 7239 2673 7265 2679
rect 7239 2641 7265 2647
rect 8863 2673 8889 2679
rect 8863 2641 8889 2647
rect 7519 2617 7545 2623
rect 7519 2585 7545 2591
rect 8695 2617 8721 2623
rect 8695 2585 8721 2591
rect 9143 2617 9169 2623
rect 13897 2591 13903 2617
rect 13929 2591 13935 2617
rect 14681 2591 14687 2617
rect 14713 2591 14719 2617
rect 15073 2591 15079 2617
rect 15105 2591 15111 2617
rect 9143 2585 9169 2591
rect 6791 2561 6817 2567
rect 6791 2529 6817 2535
rect 7799 2561 7825 2567
rect 7799 2529 7825 2535
rect 8079 2561 8105 2567
rect 8079 2529 8105 2535
rect 8415 2561 8441 2567
rect 8415 2529 8441 2535
rect 7071 2505 7097 2511
rect 7071 2473 7097 2479
rect 14407 2505 14433 2511
rect 14407 2473 14433 2479
rect 336 2365 15512 2382
rect 336 2339 1903 2365
rect 1929 2339 1955 2365
rect 1981 2339 2007 2365
rect 2033 2339 11903 2365
rect 11929 2339 11955 2365
rect 11981 2339 12007 2365
rect 12033 2339 15512 2365
rect 336 2322 15512 2339
rect 8135 2225 8161 2231
rect 7513 2199 7519 2225
rect 7545 2199 7551 2225
rect 15129 2199 15135 2225
rect 15161 2199 15167 2225
rect 8135 2193 8161 2199
rect 14681 2143 14687 2169
rect 14713 2143 14719 2169
rect 7295 2057 7321 2063
rect 7295 2025 7321 2031
rect 7855 2057 7881 2063
rect 7855 2025 7881 2031
rect 336 1973 15512 1990
rect 336 1947 2233 1973
rect 2259 1947 2285 1973
rect 2311 1947 2337 1973
rect 2363 1947 12233 1973
rect 12259 1947 12285 1973
rect 12311 1947 12337 1973
rect 12363 1947 15512 1973
rect 336 1930 15512 1947
rect 13567 1833 13593 1839
rect 13897 1807 13903 1833
rect 13929 1807 13935 1833
rect 14289 1807 14295 1833
rect 14321 1807 14327 1833
rect 13567 1801 13593 1807
rect 6959 1777 6985 1783
rect 6959 1745 6985 1751
rect 13287 1777 13313 1783
rect 14737 1751 14743 1777
rect 14769 1751 14775 1777
rect 13287 1745 13313 1751
rect 7239 1721 7265 1727
rect 7239 1689 7265 1695
rect 15191 1721 15217 1727
rect 15191 1689 15217 1695
rect 336 1581 15512 1598
rect 336 1555 1903 1581
rect 1929 1555 1955 1581
rect 1981 1555 2007 1581
rect 2033 1555 11903 1581
rect 11929 1555 11955 1581
rect 11981 1555 12007 1581
rect 12033 1555 15512 1581
rect 336 1538 15512 1555
rect 8919 1441 8945 1447
rect 8353 1415 8359 1441
rect 8385 1415 8391 1441
rect 8919 1409 8945 1415
rect 12055 1441 12081 1447
rect 12055 1409 12081 1415
rect 13007 1441 13033 1447
rect 14289 1415 14295 1441
rect 14321 1415 14327 1441
rect 15129 1415 15135 1441
rect 15161 1415 15167 1441
rect 13007 1409 13033 1415
rect 7015 1385 7041 1391
rect 7015 1353 7041 1359
rect 7687 1385 7713 1391
rect 7687 1353 7713 1359
rect 8639 1385 8665 1391
rect 13337 1359 13343 1385
rect 13369 1359 13375 1385
rect 14681 1359 14687 1385
rect 14713 1359 14719 1385
rect 8639 1353 8665 1359
rect 7295 1329 7321 1335
rect 7295 1297 7321 1303
rect 7967 1329 7993 1335
rect 13729 1303 13735 1329
rect 13761 1303 13767 1329
rect 7967 1297 7993 1303
rect 8135 1273 8161 1279
rect 8135 1241 8161 1247
rect 11775 1273 11801 1279
rect 11775 1241 11801 1247
rect 12727 1273 12753 1279
rect 12727 1241 12753 1247
rect 14519 1273 14545 1279
rect 14519 1241 14545 1247
rect 336 1189 15512 1206
rect 336 1163 2233 1189
rect 2259 1163 2285 1189
rect 2311 1163 2337 1189
rect 2363 1163 12233 1189
rect 12259 1163 12285 1189
rect 12311 1163 12337 1189
rect 12363 1163 15512 1189
rect 336 1146 15512 1163
rect 9311 1105 9337 1111
rect 9311 1073 9337 1079
rect 7407 1049 7433 1055
rect 7407 1017 7433 1023
rect 8079 1049 8105 1055
rect 8079 1017 8105 1023
rect 9591 1049 9617 1055
rect 9591 1017 9617 1023
rect 10655 1049 10681 1055
rect 10655 1017 10681 1023
rect 11103 1049 11129 1055
rect 11103 1017 11129 1023
rect 11607 1049 11633 1055
rect 11607 1017 11633 1023
rect 12839 1049 12865 1055
rect 13897 1023 13903 1049
rect 13929 1023 13935 1049
rect 14681 1023 14687 1049
rect 14713 1023 14719 1049
rect 15073 1023 15079 1049
rect 15105 1023 15111 1049
rect 12839 1017 12865 1023
rect 6959 993 6985 999
rect 6959 961 6985 967
rect 7127 993 7153 999
rect 7127 961 7153 967
rect 7799 993 7825 999
rect 7799 961 7825 967
rect 9815 993 9841 999
rect 9815 961 9841 967
rect 10375 993 10401 999
rect 10375 961 10401 967
rect 10823 993 10849 999
rect 10823 961 10849 967
rect 11327 993 11353 999
rect 11327 961 11353 967
rect 12559 993 12585 999
rect 13113 967 13119 993
rect 13145 967 13151 993
rect 12559 961 12585 967
rect 14407 937 14433 943
rect 6729 911 6735 937
rect 6761 911 6767 937
rect 10033 911 10039 937
rect 10065 911 10071 937
rect 14407 905 14433 911
rect 13623 881 13649 887
rect 13623 849 13649 855
rect 336 797 15512 814
rect 336 771 1903 797
rect 1929 771 1955 797
rect 1981 771 2007 797
rect 2033 771 11903 797
rect 11929 771 11955 797
rect 11981 771 12007 797
rect 12033 771 15512 797
rect 336 754 15512 771
rect 15191 713 15217 719
rect 15191 681 15217 687
rect 6567 657 6593 663
rect 11663 657 11689 663
rect 5553 631 5559 657
rect 5585 631 5591 657
rect 8353 631 8359 657
rect 8385 631 8391 657
rect 9137 631 9143 657
rect 9169 631 9175 657
rect 10761 631 10767 657
rect 10793 631 10799 657
rect 14345 631 14351 657
rect 14377 631 14383 657
rect 6567 625 6593 631
rect 11663 625 11689 631
rect 7855 601 7881 607
rect 6337 575 6343 601
rect 6369 575 6375 601
rect 10089 575 10095 601
rect 10121 575 10127 601
rect 12161 575 12167 601
rect 12193 575 12199 601
rect 13897 575 13903 601
rect 13929 575 13935 601
rect 14737 575 14743 601
rect 14769 575 14775 601
rect 7855 569 7881 575
rect 10201 519 10207 545
rect 10233 519 10239 545
rect 12945 519 12951 545
rect 12977 519 12983 545
rect 13337 519 13343 545
rect 13369 519 13375 545
rect 5783 489 5809 495
rect 5783 457 5809 463
rect 7575 489 7601 495
rect 7575 457 7601 463
rect 8135 489 8161 495
rect 8135 457 8161 463
rect 8919 489 8945 495
rect 8919 457 8945 463
rect 10543 489 10569 495
rect 10543 457 10569 463
rect 11383 489 11409 495
rect 11383 457 11409 463
rect 12447 489 12473 495
rect 12447 457 12473 463
rect 336 405 15512 422
rect 336 379 2233 405
rect 2259 379 2285 405
rect 2311 379 2337 405
rect 2363 379 12233 405
rect 12259 379 12285 405
rect 12311 379 12337 405
rect 12363 379 15512 405
rect 336 362 15512 379
<< via1 >>
rect 2233 6651 2259 6677
rect 2285 6651 2311 6677
rect 2337 6651 2363 6677
rect 12233 6651 12259 6677
rect 12285 6651 12311 6677
rect 12337 6651 12363 6677
rect 1079 6567 1105 6593
rect 1863 6567 1889 6593
rect 2983 6567 3009 6593
rect 3767 6567 3793 6593
rect 4887 6567 4913 6593
rect 5671 6567 5697 6593
rect 6567 6567 6593 6593
rect 7015 6567 7041 6593
rect 7855 6567 7881 6593
rect 9479 6567 9505 6593
rect 11271 6567 11297 6593
rect 12223 6567 12249 6593
rect 13007 6567 13033 6593
rect 14127 6567 14153 6593
rect 14911 6567 14937 6593
rect 3263 6511 3289 6537
rect 7575 6511 7601 6537
rect 1359 6455 1385 6481
rect 2143 6455 2169 6481
rect 3935 6455 3961 6481
rect 5167 6455 5193 6481
rect 5951 6455 5977 6481
rect 6735 6455 6761 6481
rect 9087 6455 9113 6481
rect 10823 6455 10849 6481
rect 10991 6455 11017 6481
rect 11943 6455 11969 6481
rect 12839 6455 12865 6481
rect 13959 6455 13985 6481
rect 14631 6455 14657 6481
rect 6287 6399 6313 6425
rect 8863 6399 8889 6425
rect 9703 6399 9729 6425
rect 10487 6399 10513 6425
rect 1903 6259 1929 6285
rect 1955 6259 1981 6285
rect 2007 6259 2033 6285
rect 11903 6259 11929 6285
rect 11955 6259 11981 6285
rect 12007 6259 12033 6285
rect 3655 6175 3681 6201
rect 5055 6175 5081 6201
rect 6007 6175 6033 6201
rect 6735 6175 6761 6201
rect 11383 6175 11409 6201
rect 11999 6175 12025 6201
rect 12951 6175 12977 6201
rect 14519 6175 14545 6201
rect 1919 6119 1945 6145
rect 2759 6119 2785 6145
rect 4159 6119 4185 6145
rect 9255 6119 9281 6145
rect 10039 6119 10065 6145
rect 10599 6119 10625 6145
rect 3151 6063 3177 6089
rect 7239 6063 7265 6089
rect 7687 6063 7713 6089
rect 8135 6063 8161 6089
rect 8583 6063 8609 6089
rect 8975 6063 9001 6089
rect 9479 6063 9505 6089
rect 9759 6063 9785 6089
rect 14295 6063 14321 6089
rect 2199 6007 2225 6033
rect 4551 6007 4577 6033
rect 5335 6007 5361 6033
rect 5503 6007 5529 6033
rect 7407 6007 7433 6033
rect 7855 6007 7881 6033
rect 8303 6007 8329 6033
rect 8751 6007 8777 6033
rect 10935 6007 10961 6033
rect 11103 6007 11129 6033
rect 12503 6007 12529 6033
rect 12671 6007 12697 6033
rect 13735 6007 13761 6033
rect 15303 6007 15329 6033
rect 2983 5951 3009 5977
rect 13455 5951 13481 5977
rect 15023 5951 15049 5977
rect 2233 5867 2259 5893
rect 2285 5867 2311 5893
rect 2337 5867 2363 5893
rect 12233 5867 12259 5893
rect 12285 5867 12311 5893
rect 12337 5867 12363 5893
rect 2311 5783 2337 5809
rect 3879 5783 3905 5809
rect 4775 5783 4801 5809
rect 11607 5783 11633 5809
rect 14127 5783 14153 5809
rect 1527 5727 1553 5753
rect 4495 5727 4521 5753
rect 5167 5727 5193 5753
rect 7127 5727 7153 5753
rect 1751 5671 1777 5697
rect 2591 5671 2617 5697
rect 2983 5671 3009 5697
rect 3263 5671 3289 5697
rect 4159 5671 4185 5697
rect 5559 5671 5585 5697
rect 5727 5671 5753 5697
rect 7631 5671 7657 5697
rect 9759 5671 9785 5697
rect 10263 5671 10289 5697
rect 10711 5671 10737 5697
rect 11327 5671 11353 5697
rect 12279 5671 12305 5697
rect 13063 5671 13089 5697
rect 13847 5671 13873 5697
rect 14687 5671 14713 5697
rect 6063 5615 6089 5641
rect 6623 5615 6649 5641
rect 7911 5615 7937 5641
rect 10039 5615 10065 5641
rect 10487 5615 10513 5641
rect 10935 5615 10961 5641
rect 12559 5615 12585 5641
rect 13567 5615 13593 5641
rect 15191 5559 15217 5585
rect 1903 5475 1929 5501
rect 1955 5475 1981 5501
rect 2007 5475 2033 5501
rect 11903 5475 11929 5501
rect 11955 5475 11981 5501
rect 12007 5475 12033 5501
rect 1919 5391 1945 5417
rect 3487 5391 3513 5417
rect 4271 5391 4297 5417
rect 5055 5391 5081 5417
rect 11831 5391 11857 5417
rect 12615 5391 12641 5417
rect 5783 5335 5809 5361
rect 6567 5335 6593 5361
rect 7183 5335 7209 5361
rect 8359 5335 8385 5361
rect 8807 5335 8833 5361
rect 9815 5335 9841 5361
rect 11383 5335 11409 5361
rect 13511 5335 13537 5361
rect 14463 5335 14489 5361
rect 2087 5279 2113 5305
rect 2703 5279 2729 5305
rect 2983 5279 3009 5305
rect 3767 5279 3793 5305
rect 4551 5279 4577 5305
rect 5335 5279 5361 5305
rect 7015 5279 7041 5305
rect 7463 5279 7489 5305
rect 9087 5279 9113 5305
rect 9535 5279 9561 5305
rect 9983 5279 10009 5305
rect 11103 5279 11129 5305
rect 11551 5279 11577 5305
rect 14295 5279 14321 5305
rect 6119 5223 6145 5249
rect 7967 5223 7993 5249
rect 9255 5223 9281 5249
rect 10487 5223 10513 5249
rect 10655 5223 10681 5249
rect 10935 5223 10961 5249
rect 12335 5223 12361 5249
rect 13119 5223 13145 5249
rect 14687 5223 14713 5249
rect 15079 5223 15105 5249
rect 7687 5167 7713 5193
rect 8135 5167 8161 5193
rect 10319 5167 10345 5193
rect 2233 5083 2259 5109
rect 2285 5083 2311 5109
rect 2337 5083 2363 5109
rect 12233 5083 12259 5109
rect 12285 5083 12311 5109
rect 12337 5083 12363 5109
rect 3095 4999 3121 5025
rect 3879 4999 3905 5025
rect 7183 4999 7209 5025
rect 10543 4999 10569 5025
rect 11551 4999 11577 5025
rect 12559 4999 12585 5025
rect 4943 4943 4969 4969
rect 5335 4943 5361 4969
rect 10823 4943 10849 4969
rect 14295 4943 14321 4969
rect 2031 4887 2057 4913
rect 3319 4887 3345 4913
rect 4159 4887 4185 4913
rect 6119 4887 6145 4913
rect 6679 4887 6705 4913
rect 11383 4887 11409 4913
rect 12279 4887 12305 4913
rect 13567 4887 13593 4913
rect 14015 4887 14041 4913
rect 14743 4887 14769 4913
rect 2479 4831 2505 4857
rect 6511 4831 6537 4857
rect 6903 4831 6929 4857
rect 11159 4831 11185 4857
rect 11831 4831 11857 4857
rect 13175 4831 13201 4857
rect 5615 4775 5641 4801
rect 15191 4775 15217 4801
rect 1903 4691 1929 4717
rect 1955 4691 1981 4717
rect 2007 4691 2033 4717
rect 11903 4691 11929 4717
rect 11955 4691 11981 4717
rect 12007 4691 12033 4717
rect 3711 4607 3737 4633
rect 5223 4607 5249 4633
rect 12671 4607 12697 4633
rect 13455 4607 13481 4633
rect 3039 4551 3065 4577
rect 4327 4551 4353 4577
rect 7855 4551 7881 4577
rect 11719 4551 11745 4577
rect 14519 4551 14545 4577
rect 2143 4495 2169 4521
rect 4775 4495 4801 4521
rect 6007 4495 6033 4521
rect 11999 4495 12025 4521
rect 12223 4495 12249 4521
rect 13063 4495 13089 4521
rect 14295 4495 14321 4521
rect 14687 4495 14713 4521
rect 1863 4439 1889 4465
rect 2591 4439 2617 4465
rect 3991 4439 4017 4465
rect 4943 4439 4969 4465
rect 5727 4439 5753 4465
rect 8471 4439 8497 4465
rect 13959 4439 13985 4465
rect 15079 4439 15105 4465
rect 7575 4383 7601 4409
rect 8191 4383 8217 4409
rect 11495 4383 11521 4409
rect 2233 4299 2259 4325
rect 2285 4299 2311 4325
rect 2337 4299 2363 4325
rect 12233 4299 12259 4325
rect 12285 4299 12311 4325
rect 12337 4299 12363 4325
rect 5783 4215 5809 4241
rect 6231 4215 6257 4241
rect 2311 4159 2337 4185
rect 4159 4159 4185 4185
rect 4439 4159 4465 4185
rect 5279 4159 5305 4185
rect 5503 4159 5529 4185
rect 12335 4159 12361 4185
rect 12727 4159 12753 4185
rect 2591 4103 2617 4129
rect 3375 4103 3401 4129
rect 4719 4103 4745 4129
rect 7855 4103 7881 4129
rect 13231 4103 13257 4129
rect 13903 4103 13929 4129
rect 14687 4103 14713 4129
rect 2927 4047 2953 4073
rect 3655 4047 3681 4073
rect 5055 4047 5081 4073
rect 5951 4047 5977 4073
rect 8023 4047 8049 4073
rect 13623 4047 13649 4073
rect 14407 4047 14433 4073
rect 15191 3991 15217 4017
rect 1903 3907 1929 3933
rect 1955 3907 1981 3933
rect 2007 3907 2033 3933
rect 11903 3907 11929 3933
rect 11955 3907 11981 3933
rect 12007 3907 12033 3933
rect 12895 3823 12921 3849
rect 13847 3823 13873 3849
rect 3431 3767 3457 3793
rect 4103 3767 4129 3793
rect 5167 3767 5193 3793
rect 8079 3767 8105 3793
rect 15135 3767 15161 3793
rect 5391 3711 5417 3737
rect 7799 3711 7825 3737
rect 13175 3711 13201 3737
rect 3711 3655 3737 3681
rect 7631 3655 7657 3681
rect 13343 3655 13369 3681
rect 14687 3655 14713 3681
rect 4327 3599 4353 3625
rect 7351 3599 7377 3625
rect 2233 3515 2259 3541
rect 2285 3515 2311 3541
rect 2337 3515 2363 3541
rect 12233 3515 12259 3541
rect 12285 3515 12311 3541
rect 12337 3515 12363 3541
rect 13119 3375 13145 3401
rect 3879 3319 3905 3345
rect 4103 3319 4129 3345
rect 7183 3319 7209 3345
rect 8415 3319 8441 3345
rect 13903 3319 13929 3345
rect 14687 3319 14713 3345
rect 7463 3263 7489 3289
rect 8639 3263 8665 3289
rect 13623 3263 13649 3289
rect 15191 3263 15217 3289
rect 14407 3207 14433 3233
rect 1903 3123 1929 3149
rect 1955 3123 1981 3149
rect 2007 3123 2033 3149
rect 11903 3123 11929 3149
rect 11955 3123 11981 3149
rect 12007 3123 12033 3149
rect 7519 2983 7545 3009
rect 15135 2983 15161 3009
rect 7239 2927 7265 2953
rect 14687 2871 14713 2897
rect 2233 2731 2259 2757
rect 2285 2731 2311 2757
rect 2337 2731 2363 2757
rect 12233 2731 12259 2757
rect 12285 2731 12311 2757
rect 12337 2731 12363 2757
rect 7239 2647 7265 2673
rect 8863 2647 8889 2673
rect 7519 2591 7545 2617
rect 8695 2591 8721 2617
rect 9143 2591 9169 2617
rect 13903 2591 13929 2617
rect 14687 2591 14713 2617
rect 15079 2591 15105 2617
rect 6791 2535 6817 2561
rect 7799 2535 7825 2561
rect 8079 2535 8105 2561
rect 8415 2535 8441 2561
rect 7071 2479 7097 2505
rect 14407 2479 14433 2505
rect 1903 2339 1929 2365
rect 1955 2339 1981 2365
rect 2007 2339 2033 2365
rect 11903 2339 11929 2365
rect 11955 2339 11981 2365
rect 12007 2339 12033 2365
rect 7519 2199 7545 2225
rect 8135 2199 8161 2225
rect 15135 2199 15161 2225
rect 14687 2143 14713 2169
rect 7295 2031 7321 2057
rect 7855 2031 7881 2057
rect 2233 1947 2259 1973
rect 2285 1947 2311 1973
rect 2337 1947 2363 1973
rect 12233 1947 12259 1973
rect 12285 1947 12311 1973
rect 12337 1947 12363 1973
rect 13567 1807 13593 1833
rect 13903 1807 13929 1833
rect 14295 1807 14321 1833
rect 6959 1751 6985 1777
rect 13287 1751 13313 1777
rect 14743 1751 14769 1777
rect 7239 1695 7265 1721
rect 15191 1695 15217 1721
rect 1903 1555 1929 1581
rect 1955 1555 1981 1581
rect 2007 1555 2033 1581
rect 11903 1555 11929 1581
rect 11955 1555 11981 1581
rect 12007 1555 12033 1581
rect 8359 1415 8385 1441
rect 8919 1415 8945 1441
rect 12055 1415 12081 1441
rect 13007 1415 13033 1441
rect 14295 1415 14321 1441
rect 15135 1415 15161 1441
rect 7015 1359 7041 1385
rect 7687 1359 7713 1385
rect 8639 1359 8665 1385
rect 13343 1359 13369 1385
rect 14687 1359 14713 1385
rect 7295 1303 7321 1329
rect 7967 1303 7993 1329
rect 13735 1303 13761 1329
rect 8135 1247 8161 1273
rect 11775 1247 11801 1273
rect 12727 1247 12753 1273
rect 14519 1247 14545 1273
rect 2233 1163 2259 1189
rect 2285 1163 2311 1189
rect 2337 1163 2363 1189
rect 12233 1163 12259 1189
rect 12285 1163 12311 1189
rect 12337 1163 12363 1189
rect 9311 1079 9337 1105
rect 7407 1023 7433 1049
rect 8079 1023 8105 1049
rect 9591 1023 9617 1049
rect 10655 1023 10681 1049
rect 11103 1023 11129 1049
rect 11607 1023 11633 1049
rect 12839 1023 12865 1049
rect 13903 1023 13929 1049
rect 14687 1023 14713 1049
rect 15079 1023 15105 1049
rect 6959 967 6985 993
rect 7127 967 7153 993
rect 7799 967 7825 993
rect 9815 967 9841 993
rect 10375 967 10401 993
rect 10823 967 10849 993
rect 11327 967 11353 993
rect 12559 967 12585 993
rect 13119 967 13145 993
rect 6735 911 6761 937
rect 10039 911 10065 937
rect 14407 911 14433 937
rect 13623 855 13649 881
rect 1903 771 1929 797
rect 1955 771 1981 797
rect 2007 771 2033 797
rect 11903 771 11929 797
rect 11955 771 11981 797
rect 12007 771 12033 797
rect 15191 687 15217 713
rect 5559 631 5585 657
rect 6567 631 6593 657
rect 8359 631 8385 657
rect 9143 631 9169 657
rect 10767 631 10793 657
rect 11663 631 11689 657
rect 14351 631 14377 657
rect 6343 575 6369 601
rect 7855 575 7881 601
rect 10095 575 10121 601
rect 12167 575 12193 601
rect 13903 575 13929 601
rect 14743 575 14769 601
rect 10207 519 10233 545
rect 12951 519 12977 545
rect 13343 519 13369 545
rect 5783 463 5809 489
rect 7575 463 7601 489
rect 8135 463 8161 489
rect 8919 463 8945 489
rect 10543 463 10569 489
rect 11383 463 11409 489
rect 12447 463 12473 489
rect 2233 379 2259 405
rect 2285 379 2311 405
rect 2337 379 2363 405
rect 12233 379 12259 405
rect 12285 379 12311 405
rect 12337 379 12363 405
<< metal2 >>
rect 2688 7056 2744 7112
rect 2800 7056 2856 7112
rect 2912 7056 2968 7112
rect 3024 7056 3080 7112
rect 3136 7056 3192 7112
rect 3248 7056 3304 7112
rect 3360 7056 3416 7112
rect 3472 7056 3528 7112
rect 3584 7056 3640 7112
rect 3696 7056 3752 7112
rect 3808 7056 3864 7112
rect 3920 7056 3976 7112
rect 4032 7056 4088 7112
rect 4144 7056 4200 7112
rect 4256 7056 4312 7112
rect 4368 7056 4424 7112
rect 4480 7056 4536 7112
rect 4592 7056 4648 7112
rect 4704 7056 4760 7112
rect 4816 7056 4872 7112
rect 4928 7056 4984 7112
rect 5040 7056 5096 7112
rect 5152 7056 5208 7112
rect 5264 7056 5320 7112
rect 5376 7056 5432 7112
rect 5488 7056 5544 7112
rect 5600 7056 5656 7112
rect 5712 7056 5768 7112
rect 5824 7056 5880 7112
rect 5936 7056 5992 7112
rect 6048 7056 6104 7112
rect 6160 7056 6216 7112
rect 6272 7056 6328 7112
rect 6384 7056 6440 7112
rect 6496 7056 6552 7112
rect 6608 7056 6664 7112
rect 6720 7056 6776 7112
rect 6832 7056 6888 7112
rect 6944 7056 7000 7112
rect 7056 7056 7112 7112
rect 7168 7056 7224 7112
rect 7280 7056 7336 7112
rect 7392 7056 7448 7112
rect 7504 7056 7560 7112
rect 7616 7056 7672 7112
rect 7728 7056 7784 7112
rect 7840 7056 7896 7112
rect 7952 7056 8008 7112
rect 8064 7056 8120 7112
rect 8176 7056 8232 7112
rect 8288 7056 8344 7112
rect 8400 7056 8456 7112
rect 8512 7056 8568 7112
rect 8624 7056 8680 7112
rect 8736 7056 8792 7112
rect 8848 7056 8904 7112
rect 8960 7056 9016 7112
rect 9072 7056 9128 7112
rect 9184 7056 9240 7112
rect 9296 7056 9352 7112
rect 9408 7056 9464 7112
rect 9520 7056 9576 7112
rect 9632 7056 9688 7112
rect 9744 7056 9800 7112
rect 9856 7056 9912 7112
rect 9968 7056 10024 7112
rect 10080 7056 10136 7112
rect 10192 7056 10248 7112
rect 10304 7056 10360 7112
rect 10416 7056 10472 7112
rect 10528 7056 10584 7112
rect 10640 7056 10696 7112
rect 10752 7056 10808 7112
rect 10864 7056 10920 7112
rect 10976 7056 11032 7112
rect 11088 7056 11144 7112
rect 11200 7056 11256 7112
rect 11312 7056 11368 7112
rect 11424 7056 11480 7112
rect 11536 7056 11592 7112
rect 11648 7056 11704 7112
rect 11760 7056 11816 7112
rect 11872 7056 11928 7112
rect 11984 7056 12040 7112
rect 12096 7056 12152 7112
rect 12208 7056 12264 7112
rect 12320 7056 12376 7112
rect 12432 7056 12488 7112
rect 12544 7056 12600 7112
rect 12656 7056 12712 7112
rect 12768 7056 12824 7112
rect 12880 7056 12936 7112
rect 12992 7056 13048 7112
rect 70 6986 98 6991
rect 70 826 98 6958
rect 2422 6874 2450 6879
rect 1862 6818 1890 6823
rect 294 6762 322 6767
rect 126 6538 154 6543
rect 126 1666 154 6510
rect 182 6090 210 6095
rect 182 4130 210 6062
rect 182 4102 266 4130
rect 238 3234 266 4102
rect 238 3201 266 3206
rect 294 2450 322 6734
rect 1078 6594 1106 6599
rect 1078 6547 1106 6566
rect 1862 6593 1890 6790
rect 2232 6678 2364 6683
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2232 6645 2364 6650
rect 1862 6567 1863 6593
rect 1889 6567 1890 6593
rect 1862 6561 1890 6567
rect 1358 6481 1386 6487
rect 1358 6455 1359 6481
rect 1385 6455 1386 6481
rect 1246 6314 1274 6319
rect 910 5866 938 5871
rect 406 5642 434 5647
rect 406 3682 434 5614
rect 406 3649 434 3654
rect 686 4074 714 4079
rect 686 3066 714 4046
rect 686 3033 714 3038
rect 294 2417 322 2422
rect 910 1890 938 5838
rect 1078 5418 1106 5423
rect 1078 3010 1106 5390
rect 1078 2977 1106 2982
rect 910 1857 938 1862
rect 1246 1778 1274 6286
rect 1358 5362 1386 6455
rect 2142 6481 2170 6487
rect 2142 6455 2143 6481
rect 2169 6455 2170 6481
rect 1902 6286 2034 6291
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 1902 6253 2034 6258
rect 1918 6146 1946 6151
rect 1918 6099 1946 6118
rect 1526 5810 1554 5815
rect 1526 5753 1554 5782
rect 1526 5727 1527 5753
rect 1553 5727 1554 5753
rect 1526 5721 1554 5727
rect 1358 5329 1386 5334
rect 1750 5697 1778 5703
rect 1750 5671 1751 5697
rect 1777 5671 1778 5697
rect 1246 1745 1274 1750
rect 126 1633 154 1638
rect 70 793 98 798
rect 1750 658 1778 5671
rect 1902 5502 2034 5507
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 1902 5469 2034 5474
rect 1918 5418 1946 5423
rect 1918 5371 1946 5390
rect 2086 5305 2114 5311
rect 2086 5279 2087 5305
rect 2113 5279 2114 5305
rect 2030 4914 2058 4919
rect 2030 4867 2058 4886
rect 1902 4718 2034 4723
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 1902 4685 2034 4690
rect 1862 4466 1890 4471
rect 1862 4419 1890 4438
rect 2086 4214 2114 5279
rect 2142 5250 2170 6455
rect 2198 6034 2226 6039
rect 2198 5987 2226 6006
rect 2232 5894 2364 5899
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2232 5861 2364 5866
rect 2310 5809 2338 5815
rect 2310 5783 2311 5809
rect 2337 5783 2338 5809
rect 2310 5754 2338 5783
rect 2310 5721 2338 5726
rect 2142 5217 2170 5222
rect 2232 5110 2364 5115
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2232 5077 2364 5082
rect 2422 5026 2450 6846
rect 2534 6202 2562 6207
rect 2534 5866 2562 6174
rect 2142 4998 2450 5026
rect 2478 5838 2562 5866
rect 2646 6090 2674 6095
rect 2142 4521 2170 4998
rect 2142 4495 2143 4521
rect 2169 4495 2170 4521
rect 2142 4489 2170 4495
rect 2422 4914 2450 4919
rect 2232 4326 2364 4331
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2232 4293 2364 4298
rect 2422 4214 2450 4886
rect 2478 4857 2506 5838
rect 2478 4831 2479 4857
rect 2505 4831 2506 4857
rect 2478 4825 2506 4831
rect 2590 5697 2618 5703
rect 2590 5671 2591 5697
rect 2617 5671 2618 5697
rect 2590 4690 2618 5671
rect 2646 5306 2674 6062
rect 2702 5418 2730 7056
rect 2758 6258 2786 6263
rect 2758 6145 2786 6230
rect 2758 6119 2759 6145
rect 2785 6119 2786 6145
rect 2758 6113 2786 6119
rect 2814 6034 2842 7056
rect 2926 6202 2954 7056
rect 2982 6650 3010 6655
rect 2982 6593 3010 6622
rect 2982 6567 2983 6593
rect 3009 6567 3010 6593
rect 2982 6561 3010 6567
rect 2926 6169 2954 6174
rect 2814 6006 2954 6034
rect 2702 5385 2730 5390
rect 2702 5306 2730 5311
rect 2646 5305 2730 5306
rect 2646 5279 2703 5305
rect 2729 5279 2730 5305
rect 2646 5278 2730 5279
rect 2702 5273 2730 5278
rect 2590 4657 2618 4662
rect 2590 4466 2618 4471
rect 2590 4419 2618 4438
rect 2030 4186 2114 4214
rect 2310 4186 2450 4214
rect 2030 4153 2058 4158
rect 2310 4185 2338 4186
rect 2310 4159 2311 4185
rect 2337 4159 2338 4185
rect 2310 4153 2338 4159
rect 2590 4129 2618 4135
rect 2590 4103 2591 4129
rect 2617 4103 2618 4129
rect 2590 3962 2618 4103
rect 2926 4073 2954 6006
rect 2982 5977 3010 5983
rect 2982 5951 2983 5977
rect 3009 5951 3010 5977
rect 2982 5922 3010 5951
rect 2982 5889 3010 5894
rect 2982 5698 3010 5703
rect 2982 5651 3010 5670
rect 2982 5306 3010 5311
rect 2982 5259 3010 5278
rect 3038 4577 3066 7056
rect 3150 6594 3178 7056
rect 3262 6706 3290 7056
rect 3150 6561 3178 6566
rect 3206 6678 3290 6706
rect 3318 6930 3346 6935
rect 3150 6258 3178 6263
rect 3150 6089 3178 6230
rect 3150 6063 3151 6089
rect 3177 6063 3178 6089
rect 3150 6057 3178 6063
rect 3094 5978 3122 5983
rect 3094 5025 3122 5950
rect 3206 5754 3234 6678
rect 3262 6594 3290 6599
rect 3262 6537 3290 6566
rect 3262 6511 3263 6537
rect 3289 6511 3290 6537
rect 3262 6505 3290 6511
rect 3206 5721 3234 5726
rect 3094 4999 3095 5025
rect 3121 4999 3122 5025
rect 3094 4993 3122 4999
rect 3262 5697 3290 5703
rect 3262 5671 3263 5697
rect 3289 5671 3290 5697
rect 3038 4551 3039 4577
rect 3065 4551 3066 4577
rect 3038 4545 3066 4551
rect 3262 4242 3290 5671
rect 3318 5306 3346 6902
rect 3374 6146 3402 7056
rect 3374 6113 3402 6118
rect 3486 5978 3514 7056
rect 3486 5945 3514 5950
rect 3486 5418 3514 5423
rect 3486 5371 3514 5390
rect 3318 5273 3346 5278
rect 3262 4209 3290 4214
rect 3318 4913 3346 4919
rect 3318 4887 3319 4913
rect 3345 4887 3346 4913
rect 2926 4047 2927 4073
rect 2953 4047 2954 4073
rect 2926 4041 2954 4047
rect 3318 4018 3346 4887
rect 3598 4214 3626 7056
rect 3654 6202 3682 6207
rect 3654 6155 3682 6174
rect 3710 4633 3738 7056
rect 3822 6818 3850 7056
rect 3822 6785 3850 6790
rect 3766 6762 3794 6767
rect 3766 6593 3794 6734
rect 3934 6594 3962 7056
rect 3766 6567 3767 6593
rect 3793 6567 3794 6593
rect 3766 6561 3794 6567
rect 3822 6566 3962 6594
rect 3822 5698 3850 6566
rect 3934 6481 3962 6487
rect 3934 6455 3935 6481
rect 3961 6455 3962 6481
rect 3878 5866 3906 5871
rect 3878 5809 3906 5838
rect 3878 5783 3879 5809
rect 3905 5783 3906 5809
rect 3878 5777 3906 5783
rect 3822 5665 3850 5670
rect 3934 5362 3962 6455
rect 4046 5418 4074 7056
rect 4158 6818 4186 7056
rect 4046 5385 4074 5390
rect 4102 6790 4186 6818
rect 3822 5334 3962 5362
rect 3766 5306 3794 5311
rect 3766 5259 3794 5278
rect 3710 4607 3711 4633
rect 3737 4607 3738 4633
rect 3710 4601 3738 4607
rect 3598 4186 3682 4214
rect 3318 3985 3346 3990
rect 3374 4129 3402 4135
rect 3374 4103 3375 4129
rect 3401 4103 3402 4129
rect 1902 3934 2034 3939
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2590 3929 2618 3934
rect 1902 3901 2034 3906
rect 3374 3794 3402 4103
rect 3654 4073 3682 4186
rect 3654 4047 3655 4073
rect 3681 4047 3682 4073
rect 3654 4041 3682 4047
rect 3430 3794 3458 3799
rect 3374 3793 3458 3794
rect 3374 3767 3431 3793
rect 3457 3767 3458 3793
rect 3374 3766 3458 3767
rect 3430 3761 3458 3766
rect 3374 3682 3402 3687
rect 2232 3542 2364 3547
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2232 3509 2364 3514
rect 1902 3150 2034 3155
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 1902 3117 2034 3122
rect 2232 2758 2364 2763
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2232 2725 2364 2730
rect 1902 2366 2034 2371
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 1902 2333 2034 2338
rect 3374 2002 3402 3654
rect 3710 3682 3738 3687
rect 3710 3635 3738 3654
rect 3822 3346 3850 5334
rect 4102 5306 4130 6790
rect 4158 6706 4186 6711
rect 4158 6145 4186 6678
rect 4158 6119 4159 6145
rect 4185 6119 4186 6145
rect 4158 6113 4186 6119
rect 4270 5754 4298 7056
rect 4382 6650 4410 7056
rect 4382 6617 4410 6622
rect 4494 6482 4522 7056
rect 4438 6454 4522 6482
rect 4438 5866 4466 6454
rect 4606 6202 4634 7056
rect 4718 6202 4746 7056
rect 4606 6174 4690 6202
rect 4662 6090 4690 6174
rect 4718 6169 4746 6174
rect 4774 6370 4802 6375
rect 4662 6062 4746 6090
rect 4438 5833 4466 5838
rect 4494 6034 4522 6039
rect 4270 5726 4354 5754
rect 4158 5698 4186 5703
rect 4158 5651 4186 5670
rect 3878 5278 4130 5306
rect 4158 5474 4186 5479
rect 3878 5025 3906 5278
rect 4158 5026 4186 5446
rect 4270 5418 4298 5423
rect 4270 5371 4298 5390
rect 3878 4999 3879 5025
rect 3905 4999 3906 5025
rect 3878 4993 3906 4999
rect 4046 4998 4186 5026
rect 4270 5026 4298 5031
rect 3990 4465 4018 4471
rect 3990 4439 3991 4465
rect 4017 4439 4018 4465
rect 3990 4074 4018 4439
rect 3990 4041 4018 4046
rect 3822 3313 3850 3318
rect 3878 3514 3906 3519
rect 3878 3345 3906 3486
rect 3878 3319 3879 3345
rect 3905 3319 3906 3345
rect 3878 3313 3906 3319
rect 4046 3346 4074 4998
rect 4214 4970 4242 4975
rect 4158 4914 4186 4919
rect 4158 4867 4186 4886
rect 4102 4578 4130 4583
rect 4102 3793 4130 4550
rect 4158 4298 4186 4303
rect 4158 4185 4186 4270
rect 4158 4159 4159 4185
rect 4185 4159 4186 4185
rect 4158 4153 4186 4159
rect 4102 3767 4103 3793
rect 4129 3767 4130 3793
rect 4102 3761 4130 3767
rect 4214 3738 4242 4942
rect 4214 3705 4242 3710
rect 4102 3346 4130 3351
rect 4046 3345 4130 3346
rect 4046 3319 4103 3345
rect 4129 3319 4130 3345
rect 4046 3318 4130 3319
rect 4102 3313 4130 3318
rect 4270 3066 4298 4998
rect 4326 4577 4354 5726
rect 4494 5753 4522 6006
rect 4550 6034 4578 6039
rect 4550 6033 4690 6034
rect 4550 6007 4551 6033
rect 4577 6007 4690 6033
rect 4550 6006 4690 6007
rect 4550 6001 4578 6006
rect 4494 5727 4495 5753
rect 4521 5727 4522 5753
rect 4494 5721 4522 5727
rect 4550 5922 4578 5927
rect 4550 5305 4578 5894
rect 4550 5279 4551 5305
rect 4577 5279 4578 5305
rect 4550 5273 4578 5279
rect 4326 4551 4327 4577
rect 4353 4551 4354 4577
rect 4326 4545 4354 4551
rect 4662 4466 4690 6006
rect 4718 5418 4746 6062
rect 4774 5809 4802 6342
rect 4774 5783 4775 5809
rect 4801 5783 4802 5809
rect 4774 5777 4802 5783
rect 4718 5385 4746 5390
rect 4830 5306 4858 7056
rect 4886 6818 4914 6823
rect 4886 6593 4914 6790
rect 4886 6567 4887 6593
rect 4913 6567 4914 6593
rect 4886 6561 4914 6567
rect 4830 5273 4858 5278
rect 4942 4969 4970 7056
rect 5054 6762 5082 7056
rect 5054 6729 5082 6734
rect 5166 6706 5194 7056
rect 5166 6673 5194 6678
rect 5278 6594 5306 7056
rect 5110 6566 5306 6594
rect 5054 6202 5082 6207
rect 5054 6155 5082 6174
rect 5054 5418 5082 5423
rect 5110 5418 5138 6566
rect 5166 6481 5194 6487
rect 5166 6455 5167 6481
rect 5193 6455 5194 6481
rect 5166 6258 5194 6455
rect 5166 6225 5194 6230
rect 5222 6314 5250 6319
rect 5166 6146 5194 6151
rect 5166 5753 5194 6118
rect 5166 5727 5167 5753
rect 5193 5727 5194 5753
rect 5166 5721 5194 5727
rect 5222 5586 5250 6286
rect 5334 6034 5362 6039
rect 5334 5987 5362 6006
rect 5390 5922 5418 7056
rect 5502 6146 5530 7056
rect 5614 6202 5642 7056
rect 5670 6594 5698 6599
rect 5670 6547 5698 6566
rect 5614 6169 5642 6174
rect 5502 6113 5530 6118
rect 5502 6033 5530 6039
rect 5502 6007 5503 6033
rect 5529 6007 5530 6033
rect 5502 5978 5530 6007
rect 5502 5945 5530 5950
rect 5334 5894 5418 5922
rect 5334 5642 5362 5894
rect 5726 5866 5754 7056
rect 5838 6818 5866 7056
rect 5838 6785 5866 6790
rect 5950 6594 5978 7056
rect 5894 6566 5978 6594
rect 5726 5838 5810 5866
rect 5558 5697 5586 5703
rect 5558 5671 5559 5697
rect 5585 5671 5586 5697
rect 5334 5614 5530 5642
rect 5222 5558 5418 5586
rect 5054 5417 5138 5418
rect 5054 5391 5055 5417
rect 5081 5391 5138 5417
rect 5054 5390 5138 5391
rect 5334 5474 5362 5479
rect 5054 5385 5082 5390
rect 5222 5306 5250 5311
rect 4942 4943 4943 4969
rect 4969 4943 4970 4969
rect 4942 4937 4970 4943
rect 5166 5250 5194 5255
rect 4774 4634 4802 4639
rect 4774 4521 4802 4606
rect 4774 4495 4775 4521
rect 4801 4495 4802 4521
rect 4774 4489 4802 4495
rect 4662 4433 4690 4438
rect 4942 4465 4970 4471
rect 4942 4439 4943 4465
rect 4969 4439 4970 4465
rect 4438 4186 4466 4191
rect 4438 4139 4466 4158
rect 4718 4130 4746 4135
rect 4718 4083 4746 4102
rect 4326 3626 4354 3631
rect 4326 3579 4354 3598
rect 4942 3514 4970 4439
rect 5054 4074 5082 4079
rect 5054 4027 5082 4046
rect 5166 3793 5194 5222
rect 5222 4633 5250 5278
rect 5334 5305 5362 5446
rect 5334 5279 5335 5305
rect 5361 5279 5362 5305
rect 5334 5273 5362 5279
rect 5334 5026 5362 5031
rect 5334 4969 5362 4998
rect 5334 4943 5335 4969
rect 5361 4943 5362 4969
rect 5334 4937 5362 4943
rect 5222 4607 5223 4633
rect 5249 4607 5250 4633
rect 5222 4601 5250 4607
rect 5278 4186 5306 4191
rect 5278 4139 5306 4158
rect 5166 3767 5167 3793
rect 5193 3767 5194 3793
rect 5166 3761 5194 3767
rect 5390 3737 5418 5558
rect 5502 4802 5530 5614
rect 5558 4970 5586 5671
rect 5726 5697 5754 5703
rect 5726 5671 5727 5697
rect 5753 5671 5754 5697
rect 5558 4937 5586 4942
rect 5670 5642 5698 5647
rect 5614 4802 5642 4807
rect 5502 4801 5642 4802
rect 5502 4775 5615 4801
rect 5641 4775 5642 4801
rect 5502 4774 5642 4775
rect 5614 4769 5642 4774
rect 5502 4242 5530 4247
rect 5502 4185 5530 4214
rect 5670 4214 5698 5614
rect 5726 4578 5754 5671
rect 5782 5361 5810 5838
rect 5894 5418 5922 6566
rect 5950 6482 5978 6487
rect 5950 6435 5978 6454
rect 6006 6202 6034 6207
rect 6006 6155 6034 6174
rect 5894 5385 5922 5390
rect 6006 5978 6034 5983
rect 5782 5335 5783 5361
rect 5809 5335 5810 5361
rect 5782 5329 5810 5335
rect 5726 4545 5754 4550
rect 5782 5138 5810 5143
rect 5726 4465 5754 4471
rect 5726 4439 5727 4465
rect 5753 4439 5754 4465
rect 5726 4298 5754 4439
rect 5782 4354 5810 5110
rect 5838 5082 5866 5087
rect 5838 4522 5866 5054
rect 5838 4489 5866 4494
rect 6006 4521 6034 5950
rect 6062 5641 6090 7056
rect 6174 6202 6202 7056
rect 6286 6594 6314 7056
rect 6286 6561 6314 6566
rect 6174 6169 6202 6174
rect 6286 6425 6314 6431
rect 6286 6399 6287 6425
rect 6313 6399 6314 6425
rect 6286 5698 6314 6399
rect 6286 5665 6314 5670
rect 6062 5615 6063 5641
rect 6089 5615 6090 5641
rect 6062 5609 6090 5615
rect 6398 5642 6426 7056
rect 6510 6202 6538 7056
rect 6566 6818 6594 6823
rect 6566 6593 6594 6790
rect 6566 6567 6567 6593
rect 6593 6567 6594 6593
rect 6566 6561 6594 6567
rect 6622 6594 6650 7056
rect 6734 6874 6762 7056
rect 6734 6841 6762 6846
rect 6622 6561 6650 6566
rect 6734 6482 6762 6487
rect 6510 6169 6538 6174
rect 6678 6481 6762 6482
rect 6678 6455 6735 6481
rect 6761 6455 6762 6481
rect 6678 6454 6762 6455
rect 6622 5642 6650 5647
rect 6398 5641 6650 5642
rect 6398 5615 6623 5641
rect 6649 5615 6650 5641
rect 6398 5614 6650 5615
rect 6622 5609 6650 5614
rect 6678 5530 6706 6454
rect 6734 6449 6762 6454
rect 6734 6202 6762 6207
rect 6734 6155 6762 6174
rect 6510 5502 6706 5530
rect 6118 5250 6146 5255
rect 6118 5203 6146 5222
rect 6118 4914 6146 4919
rect 6118 4867 6146 4886
rect 6510 4857 6538 5502
rect 6566 5418 6594 5423
rect 6566 5361 6594 5390
rect 6566 5335 6567 5361
rect 6593 5335 6594 5361
rect 6566 5329 6594 5335
rect 6510 4831 6511 4857
rect 6537 4831 6538 4857
rect 6510 4825 6538 4831
rect 6678 4913 6706 4919
rect 6678 4887 6679 4913
rect 6705 4887 6706 4913
rect 6678 4858 6706 4887
rect 6678 4825 6706 4830
rect 6006 4495 6007 4521
rect 6033 4495 6034 4521
rect 6006 4489 6034 4495
rect 6230 4522 6258 4527
rect 5782 4321 5810 4326
rect 5726 4265 5754 4270
rect 5782 4241 5810 4247
rect 5782 4215 5783 4241
rect 5809 4215 5810 4241
rect 5782 4214 5810 4215
rect 5670 4186 5810 4214
rect 6230 4241 6258 4494
rect 6230 4215 6231 4241
rect 6257 4215 6258 4241
rect 6230 4209 6258 4215
rect 5502 4159 5503 4185
rect 5529 4159 5530 4185
rect 5502 4153 5530 4159
rect 5950 4073 5978 4079
rect 5950 4047 5951 4073
rect 5977 4047 5978 4073
rect 5950 4018 5978 4047
rect 5950 3985 5978 3990
rect 6846 3962 6874 7056
rect 6958 6090 6986 7056
rect 7014 6594 7042 6599
rect 7014 6547 7042 6566
rect 6902 6062 6986 6090
rect 6902 5586 6930 6062
rect 6902 5558 6986 5586
rect 6902 4857 6930 4863
rect 6902 4831 6903 4857
rect 6929 4831 6930 4857
rect 6902 4690 6930 4831
rect 6902 4657 6930 4662
rect 6846 3929 6874 3934
rect 5390 3711 5391 3737
rect 5417 3711 5418 3737
rect 5390 3705 5418 3711
rect 6958 3682 6986 5558
rect 7014 5530 7042 5535
rect 7014 5305 7042 5502
rect 7014 5279 7015 5305
rect 7041 5279 7042 5305
rect 7014 5273 7042 5279
rect 7070 4130 7098 7056
rect 7126 6426 7154 6431
rect 7126 5753 7154 6398
rect 7126 5727 7127 5753
rect 7153 5727 7154 5753
rect 7126 5721 7154 5727
rect 7182 5642 7210 7056
rect 7294 6314 7322 7056
rect 7294 6281 7322 6286
rect 7406 6146 7434 7056
rect 7350 6118 7434 6146
rect 7238 6090 7266 6095
rect 7238 6043 7266 6062
rect 7182 5609 7210 5614
rect 7182 5362 7210 5367
rect 7182 5315 7210 5334
rect 7182 5194 7210 5199
rect 7182 5025 7210 5166
rect 7182 4999 7183 5025
rect 7209 4999 7210 5025
rect 7182 4993 7210 4999
rect 7350 4186 7378 6118
rect 7406 6033 7434 6039
rect 7406 6007 7407 6033
rect 7433 6007 7434 6033
rect 7406 5922 7434 6007
rect 7518 5978 7546 7056
rect 7574 6538 7602 6543
rect 7574 6491 7602 6510
rect 7518 5945 7546 5950
rect 7406 5889 7434 5894
rect 7630 5810 7658 7056
rect 7742 6370 7770 7056
rect 7854 6706 7882 7056
rect 7742 6337 7770 6342
rect 7798 6678 7882 6706
rect 7686 6146 7714 6151
rect 7686 6089 7714 6118
rect 7798 6090 7826 6678
rect 7854 6594 7882 6599
rect 7854 6547 7882 6566
rect 7686 6063 7687 6089
rect 7713 6063 7714 6089
rect 7686 6057 7714 6063
rect 7742 6062 7826 6090
rect 7574 5782 7658 5810
rect 7462 5362 7490 5367
rect 7462 5305 7490 5334
rect 7462 5279 7463 5305
rect 7489 5279 7490 5305
rect 7462 5273 7490 5279
rect 7574 4522 7602 5782
rect 7574 4489 7602 4494
rect 7630 5697 7658 5703
rect 7630 5671 7631 5697
rect 7657 5671 7658 5697
rect 7574 4410 7602 4415
rect 7574 4363 7602 4382
rect 7630 4298 7658 5671
rect 7686 5193 7714 5199
rect 7686 5167 7687 5193
rect 7713 5167 7714 5193
rect 7686 5082 7714 5167
rect 7742 5194 7770 6062
rect 7854 6034 7882 6039
rect 7742 5161 7770 5166
rect 7798 6033 7882 6034
rect 7798 6007 7855 6033
rect 7881 6007 7882 6033
rect 7798 6006 7882 6007
rect 7686 5049 7714 5054
rect 7798 4634 7826 6006
rect 7854 6001 7882 6006
rect 7910 5642 7938 5647
rect 7910 5595 7938 5614
rect 7966 5362 7994 7056
rect 8078 5754 8106 7056
rect 8134 6650 8162 6655
rect 8134 6089 8162 6622
rect 8190 6202 8218 7056
rect 8190 6169 8218 6174
rect 8302 6146 8330 7056
rect 8414 6818 8442 7056
rect 8414 6785 8442 6790
rect 8526 6594 8554 7056
rect 8638 6650 8666 7056
rect 8638 6617 8666 6622
rect 8526 6561 8554 6566
rect 8750 6538 8778 7056
rect 8302 6113 8330 6118
rect 8582 6510 8778 6538
rect 8862 6538 8890 7056
rect 8974 6594 9002 7056
rect 8974 6566 9058 6594
rect 8862 6510 9002 6538
rect 8134 6063 8135 6089
rect 8161 6063 8162 6089
rect 8134 6057 8162 6063
rect 8582 6089 8610 6510
rect 8862 6425 8890 6431
rect 8862 6399 8863 6425
rect 8889 6399 8890 6425
rect 8582 6063 8583 6089
rect 8609 6063 8610 6089
rect 8582 6057 8610 6063
rect 8806 6258 8834 6263
rect 8078 5721 8106 5726
rect 8302 6033 8330 6039
rect 8302 6007 8303 6033
rect 8329 6007 8330 6033
rect 7966 5329 7994 5334
rect 7966 5249 7994 5255
rect 7966 5223 7967 5249
rect 7993 5223 7994 5249
rect 7966 4858 7994 5223
rect 8134 5193 8162 5199
rect 8134 5167 8135 5193
rect 8161 5167 8162 5193
rect 8134 5138 8162 5167
rect 8134 5105 8162 5110
rect 7966 4825 7994 4830
rect 7798 4601 7826 4606
rect 7854 4690 7882 4695
rect 7854 4577 7882 4662
rect 7854 4551 7855 4577
rect 7881 4551 7882 4577
rect 7854 4545 7882 4551
rect 8302 4578 8330 6007
rect 8750 6033 8778 6039
rect 8750 6007 8751 6033
rect 8777 6007 8778 6033
rect 8694 5698 8722 5703
rect 8358 5361 8386 5367
rect 8358 5335 8359 5361
rect 8385 5335 8386 5361
rect 8358 4634 8386 5335
rect 8694 5026 8722 5670
rect 8750 5586 8778 6007
rect 8750 5553 8778 5558
rect 8806 5361 8834 6230
rect 8862 6090 8890 6399
rect 8862 6057 8890 6062
rect 8974 6089 9002 6510
rect 8974 6063 8975 6089
rect 9001 6063 9002 6089
rect 8974 6057 9002 6063
rect 8806 5335 8807 5361
rect 8833 5335 8834 5361
rect 8806 5329 8834 5335
rect 8974 5642 9002 5647
rect 8694 4993 8722 4998
rect 8358 4601 8386 4606
rect 8302 4545 8330 4550
rect 7350 4153 7378 4158
rect 7574 4270 7658 4298
rect 7910 4522 7938 4527
rect 7070 4097 7098 4102
rect 6958 3649 6986 3654
rect 7518 3794 7546 3799
rect 7350 3625 7378 3631
rect 7350 3599 7351 3625
rect 7377 3599 7378 3625
rect 4942 3481 4970 3486
rect 6734 3514 6762 3519
rect 4270 3033 4298 3038
rect 2232 1974 2364 1979
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 3374 1969 3402 1974
rect 2232 1941 2364 1946
rect 1902 1582 2034 1587
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 1902 1549 2034 1554
rect 1918 1498 1946 1503
rect 1750 625 1778 630
rect 1806 1470 1918 1498
rect 1134 98 1162 103
rect 1134 56 1162 70
rect 1806 56 1834 1470
rect 1918 1465 1946 1470
rect 2232 1190 2364 1195
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2232 1157 2364 1162
rect 2478 994 2506 999
rect 1902 798 2034 803
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 1902 765 2034 770
rect 2232 406 2364 411
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2232 373 2364 378
rect 2478 56 2506 966
rect 6734 937 6762 3486
rect 7350 3402 7378 3599
rect 7350 3369 7378 3374
rect 7182 3345 7210 3351
rect 7182 3319 7183 3345
rect 7209 3319 7210 3345
rect 7182 3290 7210 3319
rect 7182 3257 7210 3262
rect 7462 3290 7490 3295
rect 7462 3243 7490 3262
rect 7238 3066 7266 3071
rect 7182 2954 7210 2959
rect 7182 2674 7210 2926
rect 7238 2953 7266 3038
rect 7518 3009 7546 3766
rect 7574 3122 7602 4270
rect 7854 4129 7882 4135
rect 7854 4103 7855 4129
rect 7881 4103 7882 4129
rect 7742 4018 7770 4023
rect 7574 3089 7602 3094
rect 7630 3681 7658 3687
rect 7630 3655 7631 3681
rect 7657 3655 7658 3681
rect 7518 2983 7519 3009
rect 7545 2983 7546 3009
rect 7518 2977 7546 2983
rect 7238 2927 7239 2953
rect 7265 2927 7266 2953
rect 7238 2921 7266 2927
rect 7630 2898 7658 3655
rect 7630 2865 7658 2870
rect 7238 2674 7266 2679
rect 7182 2673 7266 2674
rect 7182 2647 7239 2673
rect 7265 2647 7266 2673
rect 7182 2646 7266 2647
rect 7238 2641 7266 2646
rect 7518 2618 7546 2623
rect 7518 2571 7546 2590
rect 6790 2561 6818 2567
rect 6790 2535 6791 2561
rect 6817 2535 6818 2561
rect 6790 2058 6818 2535
rect 6790 2025 6818 2030
rect 7070 2505 7098 2511
rect 7070 2479 7071 2505
rect 7097 2479 7098 2505
rect 7070 1890 7098 2479
rect 7518 2225 7546 2231
rect 7518 2199 7519 2225
rect 7545 2199 7546 2225
rect 7518 2114 7546 2199
rect 7518 2081 7546 2086
rect 7070 1857 7098 1862
rect 7294 2057 7322 2063
rect 7294 2031 7295 2057
rect 7321 2031 7322 2057
rect 7294 1834 7322 2031
rect 7294 1801 7322 1806
rect 6958 1777 6986 1783
rect 6958 1751 6959 1777
rect 6985 1751 6986 1777
rect 6958 1106 6986 1751
rect 7238 1722 7266 1727
rect 7238 1675 7266 1694
rect 7014 1442 7042 1447
rect 7014 1385 7042 1414
rect 7014 1359 7015 1385
rect 7041 1359 7042 1385
rect 7014 1353 7042 1359
rect 7406 1442 7434 1447
rect 7294 1329 7322 1335
rect 7294 1303 7295 1329
rect 7321 1303 7322 1329
rect 7294 1218 7322 1303
rect 7294 1185 7322 1190
rect 6958 1073 6986 1078
rect 7070 1078 7210 1106
rect 6958 994 6986 999
rect 7070 994 7098 1078
rect 6958 993 7098 994
rect 6958 967 6959 993
rect 6985 967 7098 993
rect 6958 966 7098 967
rect 7126 993 7154 999
rect 7126 967 7127 993
rect 7153 967 7154 993
rect 6958 961 6986 966
rect 6734 911 6735 937
rect 6761 911 6762 937
rect 6734 905 6762 911
rect 3822 882 3850 887
rect 3150 98 3178 103
rect 3150 56 3178 70
rect 3822 56 3850 854
rect 5558 770 5586 775
rect 5166 658 5194 663
rect 4494 434 4522 439
rect 4494 56 4522 406
rect 5166 56 5194 630
rect 5558 657 5586 742
rect 5558 631 5559 657
rect 5585 631 5586 657
rect 5558 625 5586 631
rect 6566 658 6594 663
rect 6566 611 6594 630
rect 6342 602 6370 607
rect 6342 601 6538 602
rect 6342 575 6343 601
rect 6369 575 6538 601
rect 6342 574 6538 575
rect 6342 569 6370 574
rect 5782 490 5810 495
rect 5782 489 5866 490
rect 5782 463 5783 489
rect 5809 463 5866 489
rect 5782 462 5866 463
rect 5782 457 5810 462
rect 5838 56 5866 462
rect 6510 56 6538 574
rect 7126 210 7154 967
rect 7126 177 7154 182
rect 7182 56 7210 1078
rect 7406 1049 7434 1414
rect 7686 1386 7714 1391
rect 7686 1339 7714 1358
rect 7406 1023 7407 1049
rect 7433 1023 7434 1049
rect 7406 1017 7434 1023
rect 7742 770 7770 3990
rect 7798 3738 7826 3743
rect 7798 3691 7826 3710
rect 7854 3458 7882 4103
rect 7854 3425 7882 3430
rect 7910 3346 7938 4494
rect 8470 4465 8498 4471
rect 8470 4439 8471 4465
rect 8497 4439 8498 4465
rect 8190 4409 8218 4415
rect 8190 4383 8191 4409
rect 8217 4383 8218 4409
rect 7910 3313 7938 3318
rect 8022 4073 8050 4079
rect 8022 4047 8023 4073
rect 8049 4047 8050 4073
rect 8022 3346 8050 4047
rect 8078 3906 8106 3911
rect 8078 3793 8106 3878
rect 8190 3850 8218 4383
rect 8470 4130 8498 4439
rect 8470 4097 8498 4102
rect 8190 3817 8218 3822
rect 8078 3767 8079 3793
rect 8105 3767 8106 3793
rect 8078 3761 8106 3767
rect 8974 3738 9002 5614
rect 9030 4746 9058 6566
rect 9086 6481 9114 7056
rect 9198 6594 9226 7056
rect 9198 6561 9226 6566
rect 9086 6455 9087 6481
rect 9113 6455 9114 6481
rect 9086 6449 9114 6455
rect 9254 6145 9282 6151
rect 9254 6119 9255 6145
rect 9281 6119 9282 6145
rect 9254 5530 9282 6119
rect 9310 6090 9338 7056
rect 9422 6930 9450 7056
rect 9422 6897 9450 6902
rect 9534 6706 9562 7056
rect 9310 6057 9338 6062
rect 9422 6678 9562 6706
rect 9254 5497 9282 5502
rect 9086 5306 9114 5311
rect 9086 5259 9114 5278
rect 9254 5250 9282 5255
rect 9254 5203 9282 5222
rect 9030 4713 9058 4718
rect 9086 5194 9114 5199
rect 8974 3705 9002 3710
rect 8918 3402 8946 3407
rect 8022 3313 8050 3318
rect 8414 3345 8442 3351
rect 8414 3319 8415 3345
rect 8441 3319 8442 3345
rect 8302 3066 8330 3071
rect 7798 2561 7826 2567
rect 7798 2535 7799 2561
rect 7825 2535 7826 2561
rect 7798 2282 7826 2535
rect 8078 2562 8106 2567
rect 8078 2515 8106 2534
rect 7798 2249 7826 2254
rect 8134 2226 8162 2231
rect 8134 2179 8162 2198
rect 7854 2057 7882 2063
rect 7854 2031 7855 2057
rect 7881 2031 7882 2057
rect 7854 2002 7882 2031
rect 7854 1969 7882 1974
rect 7966 1329 7994 1335
rect 7966 1303 7967 1329
rect 7993 1303 7994 1329
rect 7966 1106 7994 1303
rect 8134 1274 8162 1279
rect 8134 1227 8162 1246
rect 7966 1073 7994 1078
rect 8078 1050 8106 1055
rect 8078 1003 8106 1022
rect 7798 993 7826 999
rect 7798 967 7799 993
rect 7825 967 7826 993
rect 7798 938 7826 967
rect 7798 905 7826 910
rect 7742 737 7770 742
rect 8302 658 8330 3038
rect 8414 2674 8442 3319
rect 8414 2641 8442 2646
rect 8638 3289 8666 3295
rect 8638 3263 8639 3289
rect 8665 3263 8666 3289
rect 8414 2561 8442 2567
rect 8414 2535 8415 2561
rect 8441 2535 8442 2561
rect 8414 2506 8442 2535
rect 8414 2473 8442 2478
rect 8638 2170 8666 3263
rect 8862 3010 8890 3015
rect 8694 2674 8722 2679
rect 8694 2617 8722 2646
rect 8862 2673 8890 2982
rect 8862 2647 8863 2673
rect 8889 2647 8890 2673
rect 8862 2641 8890 2647
rect 8694 2591 8695 2617
rect 8721 2591 8722 2617
rect 8694 2585 8722 2591
rect 8638 2137 8666 2142
rect 8638 1946 8666 1951
rect 8358 1441 8386 1447
rect 8358 1415 8359 1441
rect 8385 1415 8386 1441
rect 8358 1330 8386 1415
rect 8638 1385 8666 1918
rect 8918 1441 8946 3374
rect 8918 1415 8919 1441
rect 8945 1415 8946 1441
rect 8918 1409 8946 1415
rect 8638 1359 8639 1385
rect 8665 1359 8666 1385
rect 8638 1353 8666 1359
rect 8358 1297 8386 1302
rect 8526 938 8554 943
rect 8302 625 8330 630
rect 8358 657 8386 663
rect 8358 631 8359 657
rect 8385 631 8386 657
rect 7854 602 7882 607
rect 7854 555 7882 574
rect 8358 546 8386 631
rect 8358 513 8386 518
rect 7574 489 7602 495
rect 7574 463 7575 489
rect 7601 463 7602 489
rect 7574 266 7602 463
rect 8134 490 8162 495
rect 8134 443 8162 462
rect 7574 233 7602 238
rect 7854 210 7882 215
rect 7854 56 7882 182
rect 8526 56 8554 910
rect 9086 658 9114 5166
rect 9198 4410 9226 4415
rect 9142 4074 9170 4079
rect 9142 2617 9170 4046
rect 9198 3234 9226 4382
rect 9198 3201 9226 3206
rect 9366 4298 9394 4303
rect 9142 2591 9143 2617
rect 9169 2591 9170 2617
rect 9142 2585 9170 2591
rect 9310 1498 9338 1503
rect 9310 1105 9338 1470
rect 9310 1079 9311 1105
rect 9337 1079 9338 1105
rect 9310 1073 9338 1079
rect 9142 658 9170 663
rect 9086 657 9170 658
rect 9086 631 9143 657
rect 9169 631 9170 657
rect 9086 630 9170 631
rect 9142 625 9170 630
rect 8918 489 8946 495
rect 8918 463 8919 489
rect 8945 463 8946 489
rect 8918 210 8946 463
rect 9366 434 9394 4270
rect 9422 3626 9450 6678
rect 9478 6594 9506 6599
rect 9478 6547 9506 6566
rect 9646 6482 9674 7056
rect 9478 6454 9674 6482
rect 9478 6089 9506 6454
rect 9702 6426 9730 6431
rect 9702 6379 9730 6398
rect 9758 6258 9786 7056
rect 9478 6063 9479 6089
rect 9505 6063 9506 6089
rect 9478 6057 9506 6063
rect 9702 6230 9786 6258
rect 9590 5922 9618 5927
rect 9534 5642 9562 5647
rect 9534 5305 9562 5614
rect 9534 5279 9535 5305
rect 9561 5279 9562 5305
rect 9534 5273 9562 5279
rect 9422 3593 9450 3598
rect 9590 1049 9618 5894
rect 9702 5306 9730 6230
rect 9758 6090 9786 6095
rect 9758 6043 9786 6062
rect 9814 6034 9842 6039
rect 9702 5273 9730 5278
rect 9758 5697 9786 5703
rect 9758 5671 9759 5697
rect 9785 5671 9786 5697
rect 9758 1778 9786 5671
rect 9814 5361 9842 6006
rect 9870 5642 9898 7056
rect 9870 5609 9898 5614
rect 9926 6034 9954 6039
rect 9814 5335 9815 5361
rect 9841 5335 9842 5361
rect 9814 5329 9842 5335
rect 9870 5418 9898 5423
rect 9870 3514 9898 5390
rect 9870 3481 9898 3486
rect 9758 1745 9786 1750
rect 9926 1694 9954 6006
rect 9982 5305 10010 7056
rect 10038 6482 10066 6487
rect 10038 6145 10066 6454
rect 10038 6119 10039 6145
rect 10065 6119 10066 6145
rect 10038 6113 10066 6119
rect 9982 5279 9983 5305
rect 10009 5279 10010 5305
rect 9982 5273 10010 5279
rect 10038 5641 10066 5647
rect 10038 5615 10039 5641
rect 10065 5615 10066 5641
rect 10038 4242 10066 5615
rect 10094 5026 10122 7056
rect 10206 5866 10234 7056
rect 10150 5838 10234 5866
rect 10150 5250 10178 5838
rect 10262 5697 10290 5703
rect 10262 5671 10263 5697
rect 10289 5671 10290 5697
rect 10150 5217 10178 5222
rect 10206 5530 10234 5535
rect 10094 4993 10122 4998
rect 10038 4209 10066 4214
rect 10206 2450 10234 5502
rect 10206 2417 10234 2422
rect 9926 1666 10066 1694
rect 9590 1023 9591 1049
rect 9617 1023 9618 1049
rect 9590 1017 9618 1023
rect 9814 994 9842 999
rect 9814 947 9842 966
rect 10038 937 10066 1666
rect 10262 1666 10290 5671
rect 10318 5362 10346 7056
rect 10430 6930 10458 7056
rect 10318 5329 10346 5334
rect 10374 6902 10458 6930
rect 10262 1633 10290 1638
rect 10318 5193 10346 5199
rect 10318 5167 10319 5193
rect 10345 5167 10346 5193
rect 10318 1274 10346 5167
rect 10374 5138 10402 6902
rect 10486 6425 10514 6431
rect 10486 6399 10487 6425
rect 10513 6399 10514 6425
rect 10486 6090 10514 6399
rect 10486 6057 10514 6062
rect 10542 5978 10570 7056
rect 10654 6986 10682 7056
rect 10654 6953 10682 6958
rect 10598 6930 10626 6935
rect 10598 6145 10626 6902
rect 10598 6119 10599 6145
rect 10625 6119 10626 6145
rect 10598 6113 10626 6119
rect 10766 5978 10794 7056
rect 10878 6594 10906 7056
rect 10990 6650 11018 7056
rect 10990 6617 11018 6622
rect 10878 6561 10906 6566
rect 11102 6538 11130 7056
rect 11102 6505 11130 6510
rect 10822 6482 10850 6487
rect 10822 6481 10906 6482
rect 10822 6455 10823 6481
rect 10849 6455 10906 6481
rect 10822 6454 10906 6455
rect 10822 6449 10850 6454
rect 10542 5945 10570 5950
rect 10654 5950 10794 5978
rect 10654 5754 10682 5950
rect 10430 5726 10682 5754
rect 10430 5250 10458 5726
rect 10710 5697 10738 5703
rect 10710 5671 10711 5697
rect 10737 5671 10738 5697
rect 10486 5641 10514 5647
rect 10486 5615 10487 5641
rect 10513 5615 10514 5641
rect 10486 5362 10514 5615
rect 10710 5530 10738 5671
rect 10710 5497 10738 5502
rect 10766 5586 10794 5591
rect 10486 5334 10738 5362
rect 10486 5250 10514 5255
rect 10430 5249 10514 5250
rect 10430 5223 10487 5249
rect 10513 5223 10514 5249
rect 10430 5222 10514 5223
rect 10486 5217 10514 5222
rect 10654 5250 10682 5255
rect 10654 5203 10682 5222
rect 10374 5105 10402 5110
rect 10542 5026 10570 5031
rect 10542 4979 10570 4998
rect 10710 4354 10738 5334
rect 10710 4321 10738 4326
rect 10766 3906 10794 5558
rect 10822 4970 10850 4975
rect 10822 4923 10850 4942
rect 10878 4578 10906 6454
rect 10990 6481 11018 6487
rect 10990 6455 10991 6481
rect 11017 6455 11018 6481
rect 10934 6033 10962 6039
rect 10934 6007 10935 6033
rect 10961 6007 10962 6033
rect 10934 5641 10962 6007
rect 10990 5922 11018 6455
rect 11102 6034 11130 6039
rect 11102 5987 11130 6006
rect 10990 5889 11018 5894
rect 11214 5810 11242 7056
rect 11270 6594 11298 6599
rect 11270 6547 11298 6566
rect 11326 6202 11354 7056
rect 11326 6169 11354 6174
rect 11382 6650 11410 6655
rect 11382 6201 11410 6622
rect 11382 6175 11383 6201
rect 11409 6175 11410 6201
rect 11382 6169 11410 6175
rect 11214 5777 11242 5782
rect 10934 5615 10935 5641
rect 10961 5615 10962 5641
rect 10934 5609 10962 5615
rect 11326 5697 11354 5703
rect 11326 5671 11327 5697
rect 11353 5671 11354 5697
rect 11102 5362 11130 5367
rect 11102 5305 11130 5334
rect 11102 5279 11103 5305
rect 11129 5279 11130 5305
rect 11102 5273 11130 5279
rect 11158 5306 11186 5311
rect 10934 5249 10962 5255
rect 10934 5223 10935 5249
rect 10961 5223 10962 5249
rect 10934 4914 10962 5223
rect 10934 4881 10962 4886
rect 11158 4857 11186 5278
rect 11158 4831 11159 4857
rect 11185 4831 11186 4857
rect 11158 4825 11186 4831
rect 10878 4545 10906 4550
rect 10766 3873 10794 3878
rect 10766 2058 10794 2063
rect 10038 911 10039 937
rect 10065 911 10066 937
rect 10038 905 10066 911
rect 10206 1246 10346 1274
rect 10654 1666 10682 1671
rect 10094 601 10122 607
rect 10094 575 10095 601
rect 10121 575 10122 601
rect 9366 401 9394 406
rect 9870 490 9898 495
rect 8918 177 8946 182
rect 9198 266 9226 271
rect 9198 56 9226 238
rect 9870 56 9898 462
rect 1120 0 1176 56
rect 1792 0 1848 56
rect 2464 0 2520 56
rect 3136 0 3192 56
rect 3808 0 3864 56
rect 4480 0 4536 56
rect 5152 0 5208 56
rect 5824 0 5880 56
rect 6496 0 6552 56
rect 7168 0 7224 56
rect 7840 0 7896 56
rect 8512 0 8568 56
rect 9184 0 9240 56
rect 9856 0 9912 56
rect 10094 42 10122 575
rect 10206 545 10234 1246
rect 10654 1049 10682 1638
rect 10654 1023 10655 1049
rect 10681 1023 10682 1049
rect 10654 1017 10682 1023
rect 10206 519 10207 545
rect 10233 519 10234 545
rect 10206 513 10234 519
rect 10374 993 10402 999
rect 10374 967 10375 993
rect 10401 967 10402 993
rect 10374 98 10402 967
rect 10766 657 10794 2030
rect 11326 1694 11354 5671
rect 11382 5474 11410 5479
rect 11382 5361 11410 5446
rect 11438 5418 11466 7056
rect 11550 6818 11578 7056
rect 11550 6785 11578 6790
rect 11662 6482 11690 7056
rect 11774 7042 11802 7056
rect 11774 7009 11802 7014
rect 11886 6594 11914 7056
rect 11886 6561 11914 6566
rect 11662 6449 11690 6454
rect 11942 6481 11970 6487
rect 11942 6455 11943 6481
rect 11969 6455 11970 6481
rect 11942 6370 11970 6455
rect 11998 6426 12026 7056
rect 11998 6393 12026 6398
rect 11942 6337 11970 6342
rect 11902 6286 12034 6291
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 11902 6253 12034 6258
rect 11998 6202 12026 6207
rect 11998 6155 12026 6174
rect 11606 5810 11634 5815
rect 11606 5763 11634 5782
rect 11438 5385 11466 5390
rect 11550 5754 11578 5759
rect 11382 5335 11383 5361
rect 11409 5335 11410 5361
rect 11382 5329 11410 5335
rect 11550 5305 11578 5726
rect 11902 5502 12034 5507
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 11902 5469 12034 5474
rect 12110 5474 12138 7056
rect 12222 6762 12250 7056
rect 12334 6874 12362 7056
rect 12334 6841 12362 6846
rect 12222 6729 12250 6734
rect 12232 6678 12364 6683
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12232 6645 12364 6650
rect 12110 5441 12138 5446
rect 12166 6594 12194 6599
rect 11830 5418 11858 5423
rect 11830 5371 11858 5390
rect 12166 5418 12194 6566
rect 12222 6593 12250 6599
rect 12222 6567 12223 6593
rect 12249 6567 12250 6593
rect 12222 6538 12250 6567
rect 12222 6505 12250 6510
rect 12232 5894 12364 5899
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12232 5861 12364 5866
rect 12166 5385 12194 5390
rect 12222 5810 12250 5815
rect 11550 5279 11551 5305
rect 11577 5279 11578 5305
rect 11550 5273 11578 5279
rect 12222 5194 12250 5782
rect 12446 5754 12474 7056
rect 12558 6370 12586 7056
rect 12558 6337 12586 6342
rect 12670 6202 12698 7056
rect 12670 6169 12698 6174
rect 12726 6314 12754 6319
rect 12502 6034 12530 6039
rect 12502 5987 12530 6006
rect 12670 6033 12698 6039
rect 12670 6007 12671 6033
rect 12697 6007 12698 6033
rect 12670 5866 12698 6007
rect 12670 5833 12698 5838
rect 12446 5726 12698 5754
rect 12278 5697 12306 5703
rect 12278 5671 12279 5697
rect 12305 5671 12306 5697
rect 12278 5362 12306 5671
rect 12558 5642 12586 5647
rect 12558 5595 12586 5614
rect 12278 5329 12306 5334
rect 12558 5474 12586 5479
rect 12166 5166 12250 5194
rect 12334 5249 12362 5255
rect 12334 5223 12335 5249
rect 12361 5223 12362 5249
rect 12334 5194 12362 5223
rect 11550 5138 11578 5143
rect 11550 5025 11578 5110
rect 11550 4999 11551 5025
rect 11577 4999 11578 5025
rect 11550 4993 11578 4999
rect 11774 4970 11802 4975
rect 11102 1666 11354 1694
rect 11382 4913 11410 4919
rect 11382 4887 11383 4913
rect 11409 4887 11410 4913
rect 11102 1049 11130 1666
rect 11382 1498 11410 4887
rect 11662 4914 11690 4919
rect 11494 4410 11522 4415
rect 11494 4363 11522 4382
rect 11382 1465 11410 1470
rect 11606 3682 11634 3687
rect 11102 1023 11103 1049
rect 11129 1023 11130 1049
rect 11102 1017 11130 1023
rect 11606 1049 11634 3654
rect 11606 1023 11607 1049
rect 11633 1023 11634 1049
rect 11606 1017 11634 1023
rect 10822 993 10850 999
rect 10822 967 10823 993
rect 10849 967 10850 993
rect 10822 882 10850 967
rect 11326 994 11354 999
rect 11326 947 11354 966
rect 10822 849 10850 854
rect 10766 631 10767 657
rect 10793 631 10794 657
rect 10766 625 10794 631
rect 11214 714 11242 719
rect 10542 490 10570 495
rect 10542 443 10570 462
rect 10374 65 10402 70
rect 10542 322 10570 327
rect 10542 56 10570 294
rect 11214 56 11242 686
rect 11662 657 11690 4886
rect 11718 4578 11746 4583
rect 11718 4531 11746 4550
rect 11774 1694 11802 4942
rect 11830 4857 11858 4863
rect 11830 4831 11831 4857
rect 11857 4831 11858 4857
rect 11830 4634 11858 4831
rect 11902 4718 12034 4723
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 11902 4685 12034 4690
rect 11942 4634 11970 4639
rect 12166 4634 12194 5166
rect 12334 5161 12362 5166
rect 12446 5250 12474 5255
rect 12232 5110 12364 5115
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12232 5077 12364 5082
rect 12278 4914 12306 4919
rect 12278 4867 12306 4886
rect 11830 4606 11914 4634
rect 11886 4466 11914 4606
rect 11886 4433 11914 4438
rect 11942 4298 11970 4606
rect 11998 4606 12194 4634
rect 12334 4858 12362 4863
rect 11998 4521 12026 4606
rect 11998 4495 11999 4521
rect 12025 4495 12026 4521
rect 11998 4489 12026 4495
rect 12222 4522 12250 4527
rect 12222 4475 12250 4494
rect 12334 4522 12362 4830
rect 12334 4489 12362 4494
rect 12232 4326 12364 4331
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12232 4293 12364 4298
rect 11942 4265 11970 4270
rect 12334 4242 12362 4247
rect 12334 4185 12362 4214
rect 12334 4159 12335 4185
rect 12361 4159 12362 4185
rect 12334 4153 12362 4159
rect 11902 3934 12034 3939
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 11902 3901 12034 3906
rect 12232 3542 12364 3547
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12232 3509 12364 3514
rect 11902 3150 12034 3155
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 11902 3117 12034 3122
rect 12232 2758 12364 2763
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12232 2725 12364 2730
rect 11902 2366 12034 2371
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 11902 2333 12034 2338
rect 12232 1974 12364 1979
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12232 1941 12364 1946
rect 12446 1694 12474 5222
rect 12558 5025 12586 5446
rect 12614 5418 12642 5423
rect 12614 5371 12642 5390
rect 12558 4999 12559 5025
rect 12585 4999 12586 5025
rect 12558 4993 12586 4999
rect 12614 4914 12642 4919
rect 12614 4018 12642 4886
rect 12670 4633 12698 5726
rect 12670 4607 12671 4633
rect 12697 4607 12698 4633
rect 12670 4601 12698 4607
rect 12726 4185 12754 6286
rect 12782 4858 12810 7056
rect 12894 6594 12922 7056
rect 12950 6818 12978 6823
rect 12950 6594 12978 6790
rect 13006 6706 13034 7056
rect 13454 7042 13482 7047
rect 13398 7014 13454 7042
rect 13006 6678 13090 6706
rect 13006 6594 13034 6599
rect 12950 6593 13034 6594
rect 12950 6567 13007 6593
rect 13033 6567 13034 6593
rect 12950 6566 13034 6567
rect 12894 6561 12922 6566
rect 13006 6561 13034 6566
rect 12838 6481 12866 6487
rect 12838 6455 12839 6481
rect 12865 6455 12866 6481
rect 12838 6034 12866 6455
rect 12950 6482 12978 6487
rect 12950 6201 12978 6454
rect 12950 6175 12951 6201
rect 12977 6175 12978 6201
rect 12950 6169 12978 6175
rect 13006 6146 13034 6151
rect 12838 6006 12922 6034
rect 12782 4825 12810 4830
rect 12838 5866 12866 5871
rect 12726 4159 12727 4185
rect 12753 4159 12754 4185
rect 12726 4153 12754 4159
rect 12614 3985 12642 3990
rect 12838 3066 12866 5838
rect 12894 4914 12922 6006
rect 12894 4881 12922 4886
rect 13006 4802 13034 6118
rect 13062 5810 13090 6678
rect 13398 6146 13426 7014
rect 13454 7009 13482 7014
rect 14350 6986 14378 6991
rect 13398 6113 13426 6118
rect 13510 6874 13538 6879
rect 13062 5777 13090 5782
rect 13230 5978 13258 5983
rect 12894 4774 13034 4802
rect 13062 5697 13090 5703
rect 13062 5671 13063 5697
rect 13089 5671 13090 5697
rect 12894 3849 12922 4774
rect 13062 4634 13090 5671
rect 13118 5250 13146 5255
rect 13118 5203 13146 5222
rect 13174 4858 13202 4863
rect 13174 4811 13202 4830
rect 13230 4746 13258 5950
rect 13454 5977 13482 5983
rect 13454 5951 13455 5977
rect 13481 5951 13482 5977
rect 13174 4718 13258 4746
rect 13286 5922 13314 5927
rect 13062 4606 13146 4634
rect 13062 4522 13090 4527
rect 12894 3823 12895 3849
rect 12921 3823 12922 3849
rect 12894 3817 12922 3823
rect 12950 4521 13090 4522
rect 12950 4495 13063 4521
rect 13089 4495 13090 4521
rect 12950 4494 13090 4495
rect 12838 3033 12866 3038
rect 11774 1666 11858 1694
rect 11830 1633 11858 1638
rect 12110 1666 12474 1694
rect 11902 1582 12034 1587
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 11902 1549 12034 1554
rect 11830 1498 11858 1503
rect 11662 631 11663 657
rect 11689 631 11690 657
rect 11662 625 11690 631
rect 11774 1273 11802 1279
rect 11774 1247 11775 1273
rect 11801 1247 11802 1273
rect 11382 489 11410 495
rect 11382 463 11383 489
rect 11409 463 11410 489
rect 11382 266 11410 463
rect 11774 322 11802 1247
rect 11830 714 11858 1470
rect 12054 1442 12082 1447
rect 12110 1442 12138 1666
rect 12054 1441 12138 1442
rect 12054 1415 12055 1441
rect 12081 1415 12138 1441
rect 12054 1414 12138 1415
rect 12054 1409 12082 1414
rect 12726 1274 12754 1279
rect 12614 1273 12754 1274
rect 12614 1247 12727 1273
rect 12753 1247 12754 1273
rect 12614 1246 12754 1247
rect 12232 1190 12364 1195
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12232 1157 12364 1162
rect 12558 994 12586 999
rect 12502 993 12586 994
rect 12502 967 12559 993
rect 12585 967 12586 993
rect 12502 966 12586 967
rect 11902 798 12034 803
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 11902 765 12034 770
rect 12502 714 12530 966
rect 12558 961 12586 966
rect 12614 882 12642 1246
rect 12726 1241 12754 1246
rect 12838 1050 12866 1055
rect 12950 1050 12978 4494
rect 13062 4489 13090 4494
rect 13062 4410 13090 4415
rect 13062 3402 13090 4382
rect 13118 3682 13146 4606
rect 13174 3737 13202 4718
rect 13174 3711 13175 3737
rect 13201 3711 13202 3737
rect 13174 3705 13202 3711
rect 13230 4129 13258 4135
rect 13230 4103 13231 4129
rect 13257 4103 13258 4129
rect 13118 3649 13146 3654
rect 13118 3402 13146 3407
rect 13062 3401 13146 3402
rect 13062 3375 13119 3401
rect 13145 3375 13146 3401
rect 13062 3374 13146 3375
rect 13118 3369 13146 3374
rect 13230 2226 13258 4103
rect 13230 2193 13258 2198
rect 13286 2114 13314 5894
rect 13454 5866 13482 5951
rect 13454 5833 13482 5838
rect 13398 5810 13426 5815
rect 13398 5754 13426 5782
rect 13398 5726 13482 5754
rect 13454 4633 13482 5726
rect 13510 5361 13538 6846
rect 14126 6762 14154 6767
rect 14126 6593 14154 6734
rect 14126 6567 14127 6593
rect 14153 6567 14154 6593
rect 14126 6561 14154 6567
rect 13790 6538 13818 6543
rect 13566 6426 13594 6431
rect 13566 5641 13594 6398
rect 13734 6034 13762 6039
rect 13734 5987 13762 6006
rect 13678 5866 13706 5871
rect 13566 5615 13567 5641
rect 13593 5615 13594 5641
rect 13566 5609 13594 5615
rect 13622 5642 13650 5647
rect 13510 5335 13511 5361
rect 13537 5335 13538 5361
rect 13510 5329 13538 5335
rect 13454 4607 13455 4633
rect 13481 4607 13482 4633
rect 13454 4601 13482 4607
rect 13566 4913 13594 4919
rect 13566 4887 13567 4913
rect 13593 4887 13594 4913
rect 13342 3681 13370 3687
rect 13342 3655 13343 3681
rect 13369 3655 13370 3681
rect 13342 3402 13370 3655
rect 13342 3369 13370 3374
rect 13006 2086 13314 2114
rect 13006 1441 13034 2086
rect 13454 1890 13482 1895
rect 13006 1415 13007 1441
rect 13033 1415 13034 1441
rect 13006 1409 13034 1415
rect 13286 1777 13314 1783
rect 13286 1751 13287 1777
rect 13313 1751 13314 1777
rect 12838 1049 12978 1050
rect 12838 1023 12839 1049
rect 12865 1023 12978 1049
rect 12838 1022 12978 1023
rect 12838 1017 12866 1022
rect 13118 993 13146 999
rect 13118 967 13119 993
rect 13145 967 13146 993
rect 13118 938 13146 967
rect 13118 905 13146 910
rect 11830 686 11914 714
rect 11774 289 11802 294
rect 11382 233 11410 238
rect 11886 56 11914 686
rect 12502 681 12530 686
rect 12558 854 12642 882
rect 12166 602 12194 607
rect 12166 555 12194 574
rect 12446 489 12474 495
rect 12446 463 12447 489
rect 12473 463 12474 489
rect 12232 406 12364 411
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12232 373 12364 378
rect 12446 266 12474 463
rect 12446 233 12474 238
rect 12558 56 12586 854
rect 12950 546 12978 551
rect 12950 499 12978 518
rect 13286 378 13314 1751
rect 13342 1442 13370 1447
rect 13342 1385 13370 1414
rect 13342 1359 13343 1385
rect 13369 1359 13370 1385
rect 13342 1353 13370 1359
rect 13454 1386 13482 1862
rect 13566 1833 13594 4887
rect 13622 4073 13650 5614
rect 13678 4634 13706 5838
rect 13678 4601 13706 4606
rect 13790 4214 13818 6510
rect 13958 6482 13986 6487
rect 13958 6481 14098 6482
rect 13958 6455 13959 6481
rect 13985 6455 14098 6481
rect 13958 6454 14098 6455
rect 13958 6449 13986 6454
rect 13902 5866 13930 5871
rect 13846 5697 13874 5703
rect 13846 5671 13847 5697
rect 13873 5671 13874 5697
rect 13846 5306 13874 5671
rect 13846 5273 13874 5278
rect 13902 4214 13930 5838
rect 14014 4913 14042 4919
rect 14014 4887 14015 4913
rect 14041 4887 14042 4913
rect 13622 4047 13623 4073
rect 13649 4047 13650 4073
rect 13622 4041 13650 4047
rect 13678 4186 13818 4214
rect 13846 4186 13930 4214
rect 13958 4465 13986 4471
rect 13958 4439 13959 4465
rect 13985 4439 13986 4465
rect 13622 3290 13650 3295
rect 13678 3290 13706 4186
rect 13846 3849 13874 4186
rect 13902 4129 13930 4135
rect 13902 4103 13903 4129
rect 13929 4103 13930 4129
rect 13902 4074 13930 4103
rect 13902 4041 13930 4046
rect 13846 3823 13847 3849
rect 13873 3823 13874 3849
rect 13846 3817 13874 3823
rect 13622 3289 13706 3290
rect 13622 3263 13623 3289
rect 13649 3263 13706 3289
rect 13622 3262 13706 3263
rect 13902 3345 13930 3351
rect 13902 3319 13903 3345
rect 13929 3319 13930 3345
rect 13902 3290 13930 3319
rect 13622 3257 13650 3262
rect 13902 3257 13930 3262
rect 13902 2674 13930 2679
rect 13902 2617 13930 2646
rect 13902 2591 13903 2617
rect 13929 2591 13930 2617
rect 13902 2585 13930 2591
rect 13566 1807 13567 1833
rect 13593 1807 13594 1833
rect 13566 1801 13594 1807
rect 13902 2114 13930 2119
rect 13902 1833 13930 2086
rect 13902 1807 13903 1833
rect 13929 1807 13930 1833
rect 13902 1801 13930 1807
rect 13454 1353 13482 1358
rect 13846 1722 13874 1727
rect 13734 1329 13762 1335
rect 13734 1303 13735 1329
rect 13761 1303 13762 1329
rect 13622 881 13650 887
rect 13622 855 13623 881
rect 13649 855 13650 881
rect 13622 714 13650 855
rect 13622 681 13650 686
rect 13342 545 13370 551
rect 13342 519 13343 545
rect 13369 519 13370 545
rect 13342 490 13370 519
rect 13342 457 13370 462
rect 13230 350 13314 378
rect 13230 56 13258 350
rect 13734 98 13762 1303
rect 13846 602 13874 1694
rect 13958 1722 13986 4439
rect 14014 3794 14042 4887
rect 14070 4214 14098 6454
rect 14126 6370 14154 6375
rect 14126 5809 14154 6342
rect 14294 6089 14322 6095
rect 14294 6063 14295 6089
rect 14321 6063 14322 6089
rect 14294 5922 14322 6063
rect 14294 5889 14322 5894
rect 14126 5783 14127 5809
rect 14153 5783 14154 5809
rect 14126 5777 14154 5783
rect 14294 5306 14322 5311
rect 14350 5306 14378 6958
rect 14910 6594 14938 6599
rect 14910 6547 14938 6566
rect 14630 6482 14658 6487
rect 14574 6481 14658 6482
rect 14574 6455 14631 6481
rect 14657 6455 14658 6481
rect 14574 6454 14658 6455
rect 14518 6202 14546 6207
rect 14518 6155 14546 6174
rect 14462 5698 14490 5703
rect 14294 5305 14378 5306
rect 14294 5279 14295 5305
rect 14321 5279 14378 5305
rect 14294 5278 14378 5279
rect 14406 5418 14434 5423
rect 14294 5273 14322 5278
rect 14294 5194 14322 5199
rect 14294 4969 14322 5166
rect 14294 4943 14295 4969
rect 14321 4943 14322 4969
rect 14294 4937 14322 4943
rect 14294 4521 14322 4527
rect 14294 4495 14295 4521
rect 14321 4495 14322 4521
rect 14294 4214 14322 4495
rect 14070 4186 14154 4214
rect 14014 3761 14042 3766
rect 14126 2058 14154 4186
rect 14126 2025 14154 2030
rect 14238 4186 14322 4214
rect 13958 1689 13986 1694
rect 13902 1330 13930 1335
rect 13902 1049 13930 1302
rect 13902 1023 13903 1049
rect 13929 1023 13930 1049
rect 13902 1017 13930 1023
rect 13902 602 13930 607
rect 13846 601 13930 602
rect 13846 575 13903 601
rect 13929 575 13930 601
rect 13846 574 13930 575
rect 13902 569 13930 574
rect 13734 65 13762 70
rect 13902 98 13930 103
rect 13902 56 13930 70
rect 14070 98 14098 103
rect 10094 9 10122 14
rect 10528 0 10584 56
rect 11200 0 11256 56
rect 11872 0 11928 56
rect 12544 0 12600 56
rect 13216 0 13272 56
rect 13888 0 13944 56
rect 14070 42 14098 70
rect 14238 42 14266 4186
rect 14406 4073 14434 5390
rect 14462 5361 14490 5670
rect 14462 5335 14463 5361
rect 14489 5335 14490 5361
rect 14462 5329 14490 5335
rect 14518 4578 14546 4583
rect 14574 4578 14602 6454
rect 14630 6449 14658 6454
rect 15302 6033 15330 6039
rect 15302 6007 15303 6033
rect 15329 6007 15330 6033
rect 15022 5977 15050 5983
rect 15022 5951 15023 5977
rect 15049 5951 15050 5977
rect 14686 5697 14714 5703
rect 14686 5671 14687 5697
rect 14713 5671 14714 5697
rect 14686 5586 14714 5671
rect 14686 5553 14714 5558
rect 14686 5249 14714 5255
rect 14686 5223 14687 5249
rect 14713 5223 14714 5249
rect 14686 4802 14714 5223
rect 14686 4769 14714 4774
rect 14742 4913 14770 4919
rect 14742 4887 14743 4913
rect 14769 4887 14770 4913
rect 14518 4577 14602 4578
rect 14518 4551 14519 4577
rect 14545 4551 14602 4577
rect 14518 4550 14602 4551
rect 14686 4578 14714 4583
rect 14518 4545 14546 4550
rect 14686 4521 14714 4550
rect 14686 4495 14687 4521
rect 14713 4495 14714 4521
rect 14686 4489 14714 4495
rect 14742 4522 14770 4887
rect 14742 4489 14770 4494
rect 14686 4130 14714 4135
rect 14686 4083 14714 4102
rect 14406 4047 14407 4073
rect 14433 4047 14434 4073
rect 14406 4041 14434 4047
rect 14686 3682 14714 3687
rect 14686 3635 14714 3654
rect 14686 3346 14714 3351
rect 14686 3299 14714 3318
rect 14406 3233 14434 3239
rect 14406 3207 14407 3233
rect 14433 3207 14434 3233
rect 14406 3178 14434 3207
rect 14406 3145 14434 3150
rect 14686 2898 14714 2903
rect 14686 2851 14714 2870
rect 14686 2618 14714 2623
rect 14686 2571 14714 2590
rect 14742 2562 14770 2567
rect 14406 2506 14434 2511
rect 14406 2459 14434 2478
rect 14686 2170 14714 2175
rect 14686 2123 14714 2142
rect 14294 1834 14322 1839
rect 14294 1787 14322 1806
rect 14742 1777 14770 2534
rect 14742 1751 14743 1777
rect 14769 1751 14770 1777
rect 14742 1745 14770 1751
rect 14294 1722 14322 1727
rect 14294 1441 14322 1694
rect 14294 1415 14295 1441
rect 14321 1415 14322 1441
rect 14294 1409 14322 1415
rect 14686 1386 14714 1391
rect 14686 1339 14714 1358
rect 14518 1274 14546 1279
rect 14518 1273 14602 1274
rect 14518 1247 14519 1273
rect 14545 1247 14602 1273
rect 14518 1246 14602 1247
rect 14518 1241 14546 1246
rect 14406 1162 14434 1167
rect 14350 938 14378 943
rect 14350 657 14378 910
rect 14406 937 14434 1134
rect 14406 911 14407 937
rect 14433 911 14434 937
rect 14406 905 14434 911
rect 14350 631 14351 657
rect 14377 631 14378 657
rect 14350 625 14378 631
rect 14574 56 14602 1246
rect 14686 1106 14714 1111
rect 14686 1049 14714 1078
rect 14686 1023 14687 1049
rect 14713 1023 14714 1049
rect 14686 1017 14714 1023
rect 14742 994 14770 999
rect 14742 601 14770 966
rect 15022 658 15050 5951
rect 15302 5978 15330 6007
rect 15302 5945 15330 5950
rect 15190 5585 15218 5591
rect 15190 5559 15191 5585
rect 15217 5559 15218 5585
rect 15078 5249 15106 5255
rect 15078 5223 15079 5249
rect 15105 5223 15106 5249
rect 15078 4746 15106 5223
rect 15190 4970 15218 5559
rect 15190 4937 15218 4942
rect 15078 4713 15106 4718
rect 15190 4801 15218 4807
rect 15190 4775 15191 4801
rect 15217 4775 15218 4801
rect 15190 4522 15218 4775
rect 15190 4489 15218 4494
rect 15078 4465 15106 4471
rect 15078 4439 15079 4465
rect 15105 4439 15106 4465
rect 15078 4298 15106 4439
rect 15078 4265 15106 4270
rect 15134 4074 15162 4079
rect 15134 3793 15162 4046
rect 15190 4017 15218 4023
rect 15190 3991 15191 4017
rect 15217 3991 15218 4017
rect 15190 3850 15218 3991
rect 15190 3817 15218 3822
rect 15134 3767 15135 3793
rect 15161 3767 15162 3793
rect 15134 3761 15162 3767
rect 15190 3626 15218 3631
rect 15134 3402 15162 3407
rect 15134 3009 15162 3374
rect 15190 3289 15218 3598
rect 15190 3263 15191 3289
rect 15217 3263 15218 3289
rect 15190 3257 15218 3263
rect 15134 2983 15135 3009
rect 15161 2983 15162 3009
rect 15134 2977 15162 2983
rect 15078 2954 15106 2959
rect 15078 2617 15106 2926
rect 15078 2591 15079 2617
rect 15105 2591 15106 2617
rect 15078 2585 15106 2591
rect 15134 2730 15162 2735
rect 15134 2225 15162 2702
rect 15134 2199 15135 2225
rect 15161 2199 15162 2225
rect 15134 2193 15162 2199
rect 15190 2282 15218 2287
rect 15134 2058 15162 2063
rect 15078 1610 15106 1615
rect 15078 1049 15106 1582
rect 15134 1441 15162 2030
rect 15190 1721 15218 2254
rect 15190 1695 15191 1721
rect 15217 1695 15218 1721
rect 15190 1689 15218 1695
rect 15134 1415 15135 1441
rect 15161 1415 15162 1441
rect 15134 1409 15162 1415
rect 15078 1023 15079 1049
rect 15105 1023 15106 1049
rect 15078 1017 15106 1023
rect 15190 1386 15218 1391
rect 15190 713 15218 1358
rect 15190 687 15191 713
rect 15217 687 15218 713
rect 15190 681 15218 687
rect 15022 625 15050 630
rect 14742 575 14743 601
rect 14769 575 14770 601
rect 14742 569 14770 575
rect 14070 14 14266 42
rect 14560 0 14616 56
<< via2 >>
rect 70 6958 98 6986
rect 2422 6846 2450 6874
rect 1862 6790 1890 6818
rect 294 6734 322 6762
rect 126 6510 154 6538
rect 182 6062 210 6090
rect 238 3206 266 3234
rect 1078 6593 1106 6594
rect 1078 6567 1079 6593
rect 1079 6567 1105 6593
rect 1105 6567 1106 6593
rect 1078 6566 1106 6567
rect 2232 6677 2260 6678
rect 2232 6651 2233 6677
rect 2233 6651 2259 6677
rect 2259 6651 2260 6677
rect 2232 6650 2260 6651
rect 2284 6677 2312 6678
rect 2284 6651 2285 6677
rect 2285 6651 2311 6677
rect 2311 6651 2312 6677
rect 2284 6650 2312 6651
rect 2336 6677 2364 6678
rect 2336 6651 2337 6677
rect 2337 6651 2363 6677
rect 2363 6651 2364 6677
rect 2336 6650 2364 6651
rect 1246 6286 1274 6314
rect 910 5838 938 5866
rect 406 5614 434 5642
rect 406 3654 434 3682
rect 686 4046 714 4074
rect 686 3038 714 3066
rect 294 2422 322 2450
rect 1078 5390 1106 5418
rect 1078 2982 1106 3010
rect 910 1862 938 1890
rect 1902 6285 1930 6286
rect 1902 6259 1903 6285
rect 1903 6259 1929 6285
rect 1929 6259 1930 6285
rect 1902 6258 1930 6259
rect 1954 6285 1982 6286
rect 1954 6259 1955 6285
rect 1955 6259 1981 6285
rect 1981 6259 1982 6285
rect 1954 6258 1982 6259
rect 2006 6285 2034 6286
rect 2006 6259 2007 6285
rect 2007 6259 2033 6285
rect 2033 6259 2034 6285
rect 2006 6258 2034 6259
rect 1918 6145 1946 6146
rect 1918 6119 1919 6145
rect 1919 6119 1945 6145
rect 1945 6119 1946 6145
rect 1918 6118 1946 6119
rect 1526 5782 1554 5810
rect 1358 5334 1386 5362
rect 1246 1750 1274 1778
rect 126 1638 154 1666
rect 70 798 98 826
rect 1902 5501 1930 5502
rect 1902 5475 1903 5501
rect 1903 5475 1929 5501
rect 1929 5475 1930 5501
rect 1902 5474 1930 5475
rect 1954 5501 1982 5502
rect 1954 5475 1955 5501
rect 1955 5475 1981 5501
rect 1981 5475 1982 5501
rect 1954 5474 1982 5475
rect 2006 5501 2034 5502
rect 2006 5475 2007 5501
rect 2007 5475 2033 5501
rect 2033 5475 2034 5501
rect 2006 5474 2034 5475
rect 1918 5417 1946 5418
rect 1918 5391 1919 5417
rect 1919 5391 1945 5417
rect 1945 5391 1946 5417
rect 1918 5390 1946 5391
rect 2030 4913 2058 4914
rect 2030 4887 2031 4913
rect 2031 4887 2057 4913
rect 2057 4887 2058 4913
rect 2030 4886 2058 4887
rect 1902 4717 1930 4718
rect 1902 4691 1903 4717
rect 1903 4691 1929 4717
rect 1929 4691 1930 4717
rect 1902 4690 1930 4691
rect 1954 4717 1982 4718
rect 1954 4691 1955 4717
rect 1955 4691 1981 4717
rect 1981 4691 1982 4717
rect 1954 4690 1982 4691
rect 2006 4717 2034 4718
rect 2006 4691 2007 4717
rect 2007 4691 2033 4717
rect 2033 4691 2034 4717
rect 2006 4690 2034 4691
rect 1862 4465 1890 4466
rect 1862 4439 1863 4465
rect 1863 4439 1889 4465
rect 1889 4439 1890 4465
rect 1862 4438 1890 4439
rect 2198 6033 2226 6034
rect 2198 6007 2199 6033
rect 2199 6007 2225 6033
rect 2225 6007 2226 6033
rect 2198 6006 2226 6007
rect 2232 5893 2260 5894
rect 2232 5867 2233 5893
rect 2233 5867 2259 5893
rect 2259 5867 2260 5893
rect 2232 5866 2260 5867
rect 2284 5893 2312 5894
rect 2284 5867 2285 5893
rect 2285 5867 2311 5893
rect 2311 5867 2312 5893
rect 2284 5866 2312 5867
rect 2336 5893 2364 5894
rect 2336 5867 2337 5893
rect 2337 5867 2363 5893
rect 2363 5867 2364 5893
rect 2336 5866 2364 5867
rect 2310 5726 2338 5754
rect 2142 5222 2170 5250
rect 2232 5109 2260 5110
rect 2232 5083 2233 5109
rect 2233 5083 2259 5109
rect 2259 5083 2260 5109
rect 2232 5082 2260 5083
rect 2284 5109 2312 5110
rect 2284 5083 2285 5109
rect 2285 5083 2311 5109
rect 2311 5083 2312 5109
rect 2284 5082 2312 5083
rect 2336 5109 2364 5110
rect 2336 5083 2337 5109
rect 2337 5083 2363 5109
rect 2363 5083 2364 5109
rect 2336 5082 2364 5083
rect 2534 6174 2562 6202
rect 2646 6062 2674 6090
rect 2422 4886 2450 4914
rect 2232 4325 2260 4326
rect 2232 4299 2233 4325
rect 2233 4299 2259 4325
rect 2259 4299 2260 4325
rect 2232 4298 2260 4299
rect 2284 4325 2312 4326
rect 2284 4299 2285 4325
rect 2285 4299 2311 4325
rect 2311 4299 2312 4325
rect 2284 4298 2312 4299
rect 2336 4325 2364 4326
rect 2336 4299 2337 4325
rect 2337 4299 2363 4325
rect 2363 4299 2364 4325
rect 2336 4298 2364 4299
rect 2758 6230 2786 6258
rect 2982 6622 3010 6650
rect 2926 6174 2954 6202
rect 2702 5390 2730 5418
rect 2590 4662 2618 4690
rect 2590 4465 2618 4466
rect 2590 4439 2591 4465
rect 2591 4439 2617 4465
rect 2617 4439 2618 4465
rect 2590 4438 2618 4439
rect 2030 4158 2058 4186
rect 2982 5894 3010 5922
rect 2982 5697 3010 5698
rect 2982 5671 2983 5697
rect 2983 5671 3009 5697
rect 3009 5671 3010 5697
rect 2982 5670 3010 5671
rect 2982 5305 3010 5306
rect 2982 5279 2983 5305
rect 2983 5279 3009 5305
rect 3009 5279 3010 5305
rect 2982 5278 3010 5279
rect 3150 6566 3178 6594
rect 3318 6902 3346 6930
rect 3150 6230 3178 6258
rect 3094 5950 3122 5978
rect 3262 6566 3290 6594
rect 3206 5726 3234 5754
rect 3374 6118 3402 6146
rect 3486 5950 3514 5978
rect 3486 5417 3514 5418
rect 3486 5391 3487 5417
rect 3487 5391 3513 5417
rect 3513 5391 3514 5417
rect 3486 5390 3514 5391
rect 3318 5278 3346 5306
rect 3262 4214 3290 4242
rect 3654 6201 3682 6202
rect 3654 6175 3655 6201
rect 3655 6175 3681 6201
rect 3681 6175 3682 6201
rect 3654 6174 3682 6175
rect 3822 6790 3850 6818
rect 3766 6734 3794 6762
rect 3878 5838 3906 5866
rect 3822 5670 3850 5698
rect 4046 5390 4074 5418
rect 3766 5305 3794 5306
rect 3766 5279 3767 5305
rect 3767 5279 3793 5305
rect 3793 5279 3794 5305
rect 3766 5278 3794 5279
rect 3318 3990 3346 4018
rect 1902 3933 1930 3934
rect 1902 3907 1903 3933
rect 1903 3907 1929 3933
rect 1929 3907 1930 3933
rect 1902 3906 1930 3907
rect 1954 3933 1982 3934
rect 1954 3907 1955 3933
rect 1955 3907 1981 3933
rect 1981 3907 1982 3933
rect 1954 3906 1982 3907
rect 2006 3933 2034 3934
rect 2006 3907 2007 3933
rect 2007 3907 2033 3933
rect 2033 3907 2034 3933
rect 2590 3934 2618 3962
rect 2006 3906 2034 3907
rect 3374 3654 3402 3682
rect 2232 3541 2260 3542
rect 2232 3515 2233 3541
rect 2233 3515 2259 3541
rect 2259 3515 2260 3541
rect 2232 3514 2260 3515
rect 2284 3541 2312 3542
rect 2284 3515 2285 3541
rect 2285 3515 2311 3541
rect 2311 3515 2312 3541
rect 2284 3514 2312 3515
rect 2336 3541 2364 3542
rect 2336 3515 2337 3541
rect 2337 3515 2363 3541
rect 2363 3515 2364 3541
rect 2336 3514 2364 3515
rect 1902 3149 1930 3150
rect 1902 3123 1903 3149
rect 1903 3123 1929 3149
rect 1929 3123 1930 3149
rect 1902 3122 1930 3123
rect 1954 3149 1982 3150
rect 1954 3123 1955 3149
rect 1955 3123 1981 3149
rect 1981 3123 1982 3149
rect 1954 3122 1982 3123
rect 2006 3149 2034 3150
rect 2006 3123 2007 3149
rect 2007 3123 2033 3149
rect 2033 3123 2034 3149
rect 2006 3122 2034 3123
rect 2232 2757 2260 2758
rect 2232 2731 2233 2757
rect 2233 2731 2259 2757
rect 2259 2731 2260 2757
rect 2232 2730 2260 2731
rect 2284 2757 2312 2758
rect 2284 2731 2285 2757
rect 2285 2731 2311 2757
rect 2311 2731 2312 2757
rect 2284 2730 2312 2731
rect 2336 2757 2364 2758
rect 2336 2731 2337 2757
rect 2337 2731 2363 2757
rect 2363 2731 2364 2757
rect 2336 2730 2364 2731
rect 1902 2365 1930 2366
rect 1902 2339 1903 2365
rect 1903 2339 1929 2365
rect 1929 2339 1930 2365
rect 1902 2338 1930 2339
rect 1954 2365 1982 2366
rect 1954 2339 1955 2365
rect 1955 2339 1981 2365
rect 1981 2339 1982 2365
rect 1954 2338 1982 2339
rect 2006 2365 2034 2366
rect 2006 2339 2007 2365
rect 2007 2339 2033 2365
rect 2033 2339 2034 2365
rect 2006 2338 2034 2339
rect 3710 3681 3738 3682
rect 3710 3655 3711 3681
rect 3711 3655 3737 3681
rect 3737 3655 3738 3681
rect 3710 3654 3738 3655
rect 4158 6678 4186 6706
rect 4382 6622 4410 6650
rect 4718 6174 4746 6202
rect 4774 6342 4802 6370
rect 4438 5838 4466 5866
rect 4494 6006 4522 6034
rect 4158 5697 4186 5698
rect 4158 5671 4159 5697
rect 4159 5671 4185 5697
rect 4185 5671 4186 5697
rect 4158 5670 4186 5671
rect 4158 5446 4186 5474
rect 4270 5417 4298 5418
rect 4270 5391 4271 5417
rect 4271 5391 4297 5417
rect 4297 5391 4298 5417
rect 4270 5390 4298 5391
rect 4270 4998 4298 5026
rect 3990 4046 4018 4074
rect 3822 3318 3850 3346
rect 3878 3486 3906 3514
rect 4214 4942 4242 4970
rect 4158 4913 4186 4914
rect 4158 4887 4159 4913
rect 4159 4887 4185 4913
rect 4185 4887 4186 4913
rect 4158 4886 4186 4887
rect 4102 4550 4130 4578
rect 4158 4270 4186 4298
rect 4214 3710 4242 3738
rect 4550 5894 4578 5922
rect 4718 5390 4746 5418
rect 4886 6790 4914 6818
rect 4830 5278 4858 5306
rect 5054 6734 5082 6762
rect 5166 6678 5194 6706
rect 5054 6201 5082 6202
rect 5054 6175 5055 6201
rect 5055 6175 5081 6201
rect 5081 6175 5082 6201
rect 5054 6174 5082 6175
rect 5166 6230 5194 6258
rect 5222 6286 5250 6314
rect 5166 6118 5194 6146
rect 5334 6033 5362 6034
rect 5334 6007 5335 6033
rect 5335 6007 5361 6033
rect 5361 6007 5362 6033
rect 5334 6006 5362 6007
rect 5670 6593 5698 6594
rect 5670 6567 5671 6593
rect 5671 6567 5697 6593
rect 5697 6567 5698 6593
rect 5670 6566 5698 6567
rect 5614 6174 5642 6202
rect 5502 6118 5530 6146
rect 5502 5950 5530 5978
rect 5838 6790 5866 6818
rect 5334 5446 5362 5474
rect 5222 5278 5250 5306
rect 5166 5222 5194 5250
rect 4774 4606 4802 4634
rect 4662 4438 4690 4466
rect 4438 4185 4466 4186
rect 4438 4159 4439 4185
rect 4439 4159 4465 4185
rect 4465 4159 4466 4185
rect 4438 4158 4466 4159
rect 4718 4129 4746 4130
rect 4718 4103 4719 4129
rect 4719 4103 4745 4129
rect 4745 4103 4746 4129
rect 4718 4102 4746 4103
rect 4326 3625 4354 3626
rect 4326 3599 4327 3625
rect 4327 3599 4353 3625
rect 4353 3599 4354 3625
rect 4326 3598 4354 3599
rect 5054 4073 5082 4074
rect 5054 4047 5055 4073
rect 5055 4047 5081 4073
rect 5081 4047 5082 4073
rect 5054 4046 5082 4047
rect 5334 4998 5362 5026
rect 5278 4185 5306 4186
rect 5278 4159 5279 4185
rect 5279 4159 5305 4185
rect 5305 4159 5306 4185
rect 5278 4158 5306 4159
rect 5558 4942 5586 4970
rect 5670 5614 5698 5642
rect 5502 4214 5530 4242
rect 5950 6481 5978 6482
rect 5950 6455 5951 6481
rect 5951 6455 5977 6481
rect 5977 6455 5978 6481
rect 5950 6454 5978 6455
rect 6006 6201 6034 6202
rect 6006 6175 6007 6201
rect 6007 6175 6033 6201
rect 6033 6175 6034 6201
rect 6006 6174 6034 6175
rect 5894 5390 5922 5418
rect 6006 5950 6034 5978
rect 5726 4550 5754 4578
rect 5782 5110 5810 5138
rect 5838 5054 5866 5082
rect 5838 4494 5866 4522
rect 6286 6566 6314 6594
rect 6174 6174 6202 6202
rect 6286 5670 6314 5698
rect 6566 6790 6594 6818
rect 6734 6846 6762 6874
rect 6622 6566 6650 6594
rect 6510 6174 6538 6202
rect 6734 6201 6762 6202
rect 6734 6175 6735 6201
rect 6735 6175 6761 6201
rect 6761 6175 6762 6201
rect 6734 6174 6762 6175
rect 6118 5249 6146 5250
rect 6118 5223 6119 5249
rect 6119 5223 6145 5249
rect 6145 5223 6146 5249
rect 6118 5222 6146 5223
rect 6118 4913 6146 4914
rect 6118 4887 6119 4913
rect 6119 4887 6145 4913
rect 6145 4887 6146 4913
rect 6118 4886 6146 4887
rect 6566 5390 6594 5418
rect 6678 4830 6706 4858
rect 6230 4494 6258 4522
rect 5782 4326 5810 4354
rect 5726 4270 5754 4298
rect 5950 3990 5978 4018
rect 7014 6593 7042 6594
rect 7014 6567 7015 6593
rect 7015 6567 7041 6593
rect 7041 6567 7042 6593
rect 7014 6566 7042 6567
rect 6902 4662 6930 4690
rect 6846 3934 6874 3962
rect 7014 5502 7042 5530
rect 7126 6398 7154 6426
rect 7294 6286 7322 6314
rect 7238 6089 7266 6090
rect 7238 6063 7239 6089
rect 7239 6063 7265 6089
rect 7265 6063 7266 6089
rect 7238 6062 7266 6063
rect 7182 5614 7210 5642
rect 7182 5361 7210 5362
rect 7182 5335 7183 5361
rect 7183 5335 7209 5361
rect 7209 5335 7210 5361
rect 7182 5334 7210 5335
rect 7182 5166 7210 5194
rect 7574 6537 7602 6538
rect 7574 6511 7575 6537
rect 7575 6511 7601 6537
rect 7601 6511 7602 6537
rect 7574 6510 7602 6511
rect 7518 5950 7546 5978
rect 7406 5894 7434 5922
rect 7742 6342 7770 6370
rect 7686 6118 7714 6146
rect 7854 6593 7882 6594
rect 7854 6567 7855 6593
rect 7855 6567 7881 6593
rect 7881 6567 7882 6593
rect 7854 6566 7882 6567
rect 7462 5334 7490 5362
rect 7574 4494 7602 4522
rect 7574 4409 7602 4410
rect 7574 4383 7575 4409
rect 7575 4383 7601 4409
rect 7601 4383 7602 4409
rect 7574 4382 7602 4383
rect 7742 5166 7770 5194
rect 7686 5054 7714 5082
rect 7910 5641 7938 5642
rect 7910 5615 7911 5641
rect 7911 5615 7937 5641
rect 7937 5615 7938 5641
rect 7910 5614 7938 5615
rect 8134 6622 8162 6650
rect 8190 6174 8218 6202
rect 8414 6790 8442 6818
rect 8638 6622 8666 6650
rect 8526 6566 8554 6594
rect 8302 6118 8330 6146
rect 8806 6230 8834 6258
rect 8078 5726 8106 5754
rect 7966 5334 7994 5362
rect 8134 5110 8162 5138
rect 7966 4830 7994 4858
rect 7798 4606 7826 4634
rect 7854 4662 7882 4690
rect 8694 5670 8722 5698
rect 8750 5558 8778 5586
rect 8862 6062 8890 6090
rect 8974 5614 9002 5642
rect 8694 4998 8722 5026
rect 8358 4606 8386 4634
rect 8302 4550 8330 4578
rect 7350 4158 7378 4186
rect 7910 4494 7938 4522
rect 7070 4102 7098 4130
rect 6958 3654 6986 3682
rect 7518 3766 7546 3794
rect 4942 3486 4970 3514
rect 6734 3486 6762 3514
rect 4270 3038 4298 3066
rect 2232 1973 2260 1974
rect 2232 1947 2233 1973
rect 2233 1947 2259 1973
rect 2259 1947 2260 1973
rect 2232 1946 2260 1947
rect 2284 1973 2312 1974
rect 2284 1947 2285 1973
rect 2285 1947 2311 1973
rect 2311 1947 2312 1973
rect 2284 1946 2312 1947
rect 2336 1973 2364 1974
rect 2336 1947 2337 1973
rect 2337 1947 2363 1973
rect 2363 1947 2364 1973
rect 3374 1974 3402 2002
rect 2336 1946 2364 1947
rect 1902 1581 1930 1582
rect 1902 1555 1903 1581
rect 1903 1555 1929 1581
rect 1929 1555 1930 1581
rect 1902 1554 1930 1555
rect 1954 1581 1982 1582
rect 1954 1555 1955 1581
rect 1955 1555 1981 1581
rect 1981 1555 1982 1581
rect 1954 1554 1982 1555
rect 2006 1581 2034 1582
rect 2006 1555 2007 1581
rect 2007 1555 2033 1581
rect 2033 1555 2034 1581
rect 2006 1554 2034 1555
rect 1750 630 1778 658
rect 1918 1470 1946 1498
rect 1134 70 1162 98
rect 2232 1189 2260 1190
rect 2232 1163 2233 1189
rect 2233 1163 2259 1189
rect 2259 1163 2260 1189
rect 2232 1162 2260 1163
rect 2284 1189 2312 1190
rect 2284 1163 2285 1189
rect 2285 1163 2311 1189
rect 2311 1163 2312 1189
rect 2284 1162 2312 1163
rect 2336 1189 2364 1190
rect 2336 1163 2337 1189
rect 2337 1163 2363 1189
rect 2363 1163 2364 1189
rect 2336 1162 2364 1163
rect 2478 966 2506 994
rect 1902 797 1930 798
rect 1902 771 1903 797
rect 1903 771 1929 797
rect 1929 771 1930 797
rect 1902 770 1930 771
rect 1954 797 1982 798
rect 1954 771 1955 797
rect 1955 771 1981 797
rect 1981 771 1982 797
rect 1954 770 1982 771
rect 2006 797 2034 798
rect 2006 771 2007 797
rect 2007 771 2033 797
rect 2033 771 2034 797
rect 2006 770 2034 771
rect 2232 405 2260 406
rect 2232 379 2233 405
rect 2233 379 2259 405
rect 2259 379 2260 405
rect 2232 378 2260 379
rect 2284 405 2312 406
rect 2284 379 2285 405
rect 2285 379 2311 405
rect 2311 379 2312 405
rect 2284 378 2312 379
rect 2336 405 2364 406
rect 2336 379 2337 405
rect 2337 379 2363 405
rect 2363 379 2364 405
rect 2336 378 2364 379
rect 7350 3374 7378 3402
rect 7182 3262 7210 3290
rect 7462 3289 7490 3290
rect 7462 3263 7463 3289
rect 7463 3263 7489 3289
rect 7489 3263 7490 3289
rect 7462 3262 7490 3263
rect 7238 3038 7266 3066
rect 7182 2926 7210 2954
rect 7742 3990 7770 4018
rect 7574 3094 7602 3122
rect 7630 2870 7658 2898
rect 7518 2617 7546 2618
rect 7518 2591 7519 2617
rect 7519 2591 7545 2617
rect 7545 2591 7546 2617
rect 7518 2590 7546 2591
rect 6790 2030 6818 2058
rect 7518 2086 7546 2114
rect 7070 1862 7098 1890
rect 7294 1806 7322 1834
rect 7238 1721 7266 1722
rect 7238 1695 7239 1721
rect 7239 1695 7265 1721
rect 7265 1695 7266 1721
rect 7238 1694 7266 1695
rect 7014 1414 7042 1442
rect 7406 1414 7434 1442
rect 7294 1190 7322 1218
rect 6958 1078 6986 1106
rect 3822 854 3850 882
rect 3150 70 3178 98
rect 5558 742 5586 770
rect 5166 630 5194 658
rect 4494 406 4522 434
rect 6566 657 6594 658
rect 6566 631 6567 657
rect 6567 631 6593 657
rect 6593 631 6594 657
rect 6566 630 6594 631
rect 7126 182 7154 210
rect 7686 1385 7714 1386
rect 7686 1359 7687 1385
rect 7687 1359 7713 1385
rect 7713 1359 7714 1385
rect 7686 1358 7714 1359
rect 7798 3737 7826 3738
rect 7798 3711 7799 3737
rect 7799 3711 7825 3737
rect 7825 3711 7826 3737
rect 7798 3710 7826 3711
rect 7854 3430 7882 3458
rect 7910 3318 7938 3346
rect 8078 3878 8106 3906
rect 8470 4102 8498 4130
rect 8190 3822 8218 3850
rect 9198 6566 9226 6594
rect 9422 6902 9450 6930
rect 9310 6062 9338 6090
rect 9254 5502 9282 5530
rect 9086 5305 9114 5306
rect 9086 5279 9087 5305
rect 9087 5279 9113 5305
rect 9113 5279 9114 5305
rect 9086 5278 9114 5279
rect 9254 5249 9282 5250
rect 9254 5223 9255 5249
rect 9255 5223 9281 5249
rect 9281 5223 9282 5249
rect 9254 5222 9282 5223
rect 9030 4718 9058 4746
rect 9086 5166 9114 5194
rect 8974 3710 9002 3738
rect 8918 3374 8946 3402
rect 8022 3318 8050 3346
rect 8302 3038 8330 3066
rect 8078 2561 8106 2562
rect 8078 2535 8079 2561
rect 8079 2535 8105 2561
rect 8105 2535 8106 2561
rect 8078 2534 8106 2535
rect 7798 2254 7826 2282
rect 8134 2225 8162 2226
rect 8134 2199 8135 2225
rect 8135 2199 8161 2225
rect 8161 2199 8162 2225
rect 8134 2198 8162 2199
rect 7854 1974 7882 2002
rect 8134 1273 8162 1274
rect 8134 1247 8135 1273
rect 8135 1247 8161 1273
rect 8161 1247 8162 1273
rect 8134 1246 8162 1247
rect 7966 1078 7994 1106
rect 8078 1049 8106 1050
rect 8078 1023 8079 1049
rect 8079 1023 8105 1049
rect 8105 1023 8106 1049
rect 8078 1022 8106 1023
rect 7798 910 7826 938
rect 7742 742 7770 770
rect 8414 2646 8442 2674
rect 8414 2478 8442 2506
rect 8862 2982 8890 3010
rect 8694 2646 8722 2674
rect 8638 2142 8666 2170
rect 8638 1918 8666 1946
rect 8358 1302 8386 1330
rect 8526 910 8554 938
rect 8302 630 8330 658
rect 7854 601 7882 602
rect 7854 575 7855 601
rect 7855 575 7881 601
rect 7881 575 7882 601
rect 7854 574 7882 575
rect 8358 518 8386 546
rect 8134 489 8162 490
rect 8134 463 8135 489
rect 8135 463 8161 489
rect 8161 463 8162 489
rect 8134 462 8162 463
rect 7574 238 7602 266
rect 7854 182 7882 210
rect 9198 4382 9226 4410
rect 9142 4046 9170 4074
rect 9198 3206 9226 3234
rect 9366 4270 9394 4298
rect 9310 1470 9338 1498
rect 9478 6593 9506 6594
rect 9478 6567 9479 6593
rect 9479 6567 9505 6593
rect 9505 6567 9506 6593
rect 9478 6566 9506 6567
rect 9702 6425 9730 6426
rect 9702 6399 9703 6425
rect 9703 6399 9729 6425
rect 9729 6399 9730 6425
rect 9702 6398 9730 6399
rect 9590 5894 9618 5922
rect 9534 5614 9562 5642
rect 9422 3598 9450 3626
rect 9758 6089 9786 6090
rect 9758 6063 9759 6089
rect 9759 6063 9785 6089
rect 9785 6063 9786 6089
rect 9758 6062 9786 6063
rect 9814 6006 9842 6034
rect 9702 5278 9730 5306
rect 9870 5614 9898 5642
rect 9926 6006 9954 6034
rect 9870 5390 9898 5418
rect 9870 3486 9898 3514
rect 9758 1750 9786 1778
rect 10038 6454 10066 6482
rect 10150 5222 10178 5250
rect 10206 5502 10234 5530
rect 10094 4998 10122 5026
rect 10038 4214 10066 4242
rect 10206 2422 10234 2450
rect 9814 993 9842 994
rect 9814 967 9815 993
rect 9815 967 9841 993
rect 9841 967 9842 993
rect 9814 966 9842 967
rect 10318 5334 10346 5362
rect 10262 1638 10290 1666
rect 10486 6062 10514 6090
rect 10654 6958 10682 6986
rect 10598 6902 10626 6930
rect 10990 6622 11018 6650
rect 10878 6566 10906 6594
rect 11102 6510 11130 6538
rect 10542 5950 10570 5978
rect 10710 5502 10738 5530
rect 10766 5558 10794 5586
rect 10654 5249 10682 5250
rect 10654 5223 10655 5249
rect 10655 5223 10681 5249
rect 10681 5223 10682 5249
rect 10654 5222 10682 5223
rect 10374 5110 10402 5138
rect 10542 5025 10570 5026
rect 10542 4999 10543 5025
rect 10543 4999 10569 5025
rect 10569 4999 10570 5025
rect 10542 4998 10570 4999
rect 10710 4326 10738 4354
rect 10822 4969 10850 4970
rect 10822 4943 10823 4969
rect 10823 4943 10849 4969
rect 10849 4943 10850 4969
rect 10822 4942 10850 4943
rect 11102 6033 11130 6034
rect 11102 6007 11103 6033
rect 11103 6007 11129 6033
rect 11129 6007 11130 6033
rect 11102 6006 11130 6007
rect 10990 5894 11018 5922
rect 11270 6593 11298 6594
rect 11270 6567 11271 6593
rect 11271 6567 11297 6593
rect 11297 6567 11298 6593
rect 11270 6566 11298 6567
rect 11326 6174 11354 6202
rect 11382 6622 11410 6650
rect 11214 5782 11242 5810
rect 11102 5334 11130 5362
rect 11158 5278 11186 5306
rect 10934 4886 10962 4914
rect 10878 4550 10906 4578
rect 10766 3878 10794 3906
rect 10766 2030 10794 2058
rect 10654 1638 10682 1666
rect 9366 406 9394 434
rect 9870 462 9898 490
rect 8918 182 8946 210
rect 9198 238 9226 266
rect 11382 5446 11410 5474
rect 11550 6790 11578 6818
rect 11774 7014 11802 7042
rect 11886 6566 11914 6594
rect 11662 6454 11690 6482
rect 11998 6398 12026 6426
rect 11942 6342 11970 6370
rect 11902 6285 11930 6286
rect 11902 6259 11903 6285
rect 11903 6259 11929 6285
rect 11929 6259 11930 6285
rect 11902 6258 11930 6259
rect 11954 6285 11982 6286
rect 11954 6259 11955 6285
rect 11955 6259 11981 6285
rect 11981 6259 11982 6285
rect 11954 6258 11982 6259
rect 12006 6285 12034 6286
rect 12006 6259 12007 6285
rect 12007 6259 12033 6285
rect 12033 6259 12034 6285
rect 12006 6258 12034 6259
rect 11998 6201 12026 6202
rect 11998 6175 11999 6201
rect 11999 6175 12025 6201
rect 12025 6175 12026 6201
rect 11998 6174 12026 6175
rect 11606 5809 11634 5810
rect 11606 5783 11607 5809
rect 11607 5783 11633 5809
rect 11633 5783 11634 5809
rect 11606 5782 11634 5783
rect 11438 5390 11466 5418
rect 11550 5726 11578 5754
rect 11902 5501 11930 5502
rect 11902 5475 11903 5501
rect 11903 5475 11929 5501
rect 11929 5475 11930 5501
rect 11902 5474 11930 5475
rect 11954 5501 11982 5502
rect 11954 5475 11955 5501
rect 11955 5475 11981 5501
rect 11981 5475 11982 5501
rect 11954 5474 11982 5475
rect 12006 5501 12034 5502
rect 12006 5475 12007 5501
rect 12007 5475 12033 5501
rect 12033 5475 12034 5501
rect 12006 5474 12034 5475
rect 12334 6846 12362 6874
rect 12222 6734 12250 6762
rect 12232 6677 12260 6678
rect 12232 6651 12233 6677
rect 12233 6651 12259 6677
rect 12259 6651 12260 6677
rect 12232 6650 12260 6651
rect 12284 6677 12312 6678
rect 12284 6651 12285 6677
rect 12285 6651 12311 6677
rect 12311 6651 12312 6677
rect 12284 6650 12312 6651
rect 12336 6677 12364 6678
rect 12336 6651 12337 6677
rect 12337 6651 12363 6677
rect 12363 6651 12364 6677
rect 12336 6650 12364 6651
rect 12110 5446 12138 5474
rect 12166 6566 12194 6594
rect 11830 5417 11858 5418
rect 11830 5391 11831 5417
rect 11831 5391 11857 5417
rect 11857 5391 11858 5417
rect 11830 5390 11858 5391
rect 12222 6510 12250 6538
rect 12232 5893 12260 5894
rect 12232 5867 12233 5893
rect 12233 5867 12259 5893
rect 12259 5867 12260 5893
rect 12232 5866 12260 5867
rect 12284 5893 12312 5894
rect 12284 5867 12285 5893
rect 12285 5867 12311 5893
rect 12311 5867 12312 5893
rect 12284 5866 12312 5867
rect 12336 5893 12364 5894
rect 12336 5867 12337 5893
rect 12337 5867 12363 5893
rect 12363 5867 12364 5893
rect 12336 5866 12364 5867
rect 12166 5390 12194 5418
rect 12222 5782 12250 5810
rect 12558 6342 12586 6370
rect 12670 6174 12698 6202
rect 12726 6286 12754 6314
rect 12502 6033 12530 6034
rect 12502 6007 12503 6033
rect 12503 6007 12529 6033
rect 12529 6007 12530 6033
rect 12502 6006 12530 6007
rect 12670 5838 12698 5866
rect 12558 5641 12586 5642
rect 12558 5615 12559 5641
rect 12559 5615 12585 5641
rect 12585 5615 12586 5641
rect 12558 5614 12586 5615
rect 12278 5334 12306 5362
rect 12558 5446 12586 5474
rect 12334 5166 12362 5194
rect 11550 5110 11578 5138
rect 11774 4942 11802 4970
rect 11662 4886 11690 4914
rect 11494 4409 11522 4410
rect 11494 4383 11495 4409
rect 11495 4383 11521 4409
rect 11521 4383 11522 4409
rect 11494 4382 11522 4383
rect 11382 1470 11410 1498
rect 11606 3654 11634 3682
rect 11326 993 11354 994
rect 11326 967 11327 993
rect 11327 967 11353 993
rect 11353 967 11354 993
rect 11326 966 11354 967
rect 10822 854 10850 882
rect 11214 686 11242 714
rect 10542 489 10570 490
rect 10542 463 10543 489
rect 10543 463 10569 489
rect 10569 463 10570 489
rect 10542 462 10570 463
rect 10374 70 10402 98
rect 10542 294 10570 322
rect 11718 4577 11746 4578
rect 11718 4551 11719 4577
rect 11719 4551 11745 4577
rect 11745 4551 11746 4577
rect 11718 4550 11746 4551
rect 11902 4717 11930 4718
rect 11902 4691 11903 4717
rect 11903 4691 11929 4717
rect 11929 4691 11930 4717
rect 11902 4690 11930 4691
rect 11954 4717 11982 4718
rect 11954 4691 11955 4717
rect 11955 4691 11981 4717
rect 11981 4691 11982 4717
rect 11954 4690 11982 4691
rect 12006 4717 12034 4718
rect 12006 4691 12007 4717
rect 12007 4691 12033 4717
rect 12033 4691 12034 4717
rect 12006 4690 12034 4691
rect 12446 5222 12474 5250
rect 12232 5109 12260 5110
rect 12232 5083 12233 5109
rect 12233 5083 12259 5109
rect 12259 5083 12260 5109
rect 12232 5082 12260 5083
rect 12284 5109 12312 5110
rect 12284 5083 12285 5109
rect 12285 5083 12311 5109
rect 12311 5083 12312 5109
rect 12284 5082 12312 5083
rect 12336 5109 12364 5110
rect 12336 5083 12337 5109
rect 12337 5083 12363 5109
rect 12363 5083 12364 5109
rect 12336 5082 12364 5083
rect 12278 4913 12306 4914
rect 12278 4887 12279 4913
rect 12279 4887 12305 4913
rect 12305 4887 12306 4913
rect 12278 4886 12306 4887
rect 11886 4438 11914 4466
rect 11942 4606 11970 4634
rect 12334 4830 12362 4858
rect 12222 4521 12250 4522
rect 12222 4495 12223 4521
rect 12223 4495 12249 4521
rect 12249 4495 12250 4521
rect 12222 4494 12250 4495
rect 12334 4494 12362 4522
rect 11942 4270 11970 4298
rect 12232 4325 12260 4326
rect 12232 4299 12233 4325
rect 12233 4299 12259 4325
rect 12259 4299 12260 4325
rect 12232 4298 12260 4299
rect 12284 4325 12312 4326
rect 12284 4299 12285 4325
rect 12285 4299 12311 4325
rect 12311 4299 12312 4325
rect 12284 4298 12312 4299
rect 12336 4325 12364 4326
rect 12336 4299 12337 4325
rect 12337 4299 12363 4325
rect 12363 4299 12364 4325
rect 12336 4298 12364 4299
rect 12334 4214 12362 4242
rect 11902 3933 11930 3934
rect 11902 3907 11903 3933
rect 11903 3907 11929 3933
rect 11929 3907 11930 3933
rect 11902 3906 11930 3907
rect 11954 3933 11982 3934
rect 11954 3907 11955 3933
rect 11955 3907 11981 3933
rect 11981 3907 11982 3933
rect 11954 3906 11982 3907
rect 12006 3933 12034 3934
rect 12006 3907 12007 3933
rect 12007 3907 12033 3933
rect 12033 3907 12034 3933
rect 12006 3906 12034 3907
rect 12232 3541 12260 3542
rect 12232 3515 12233 3541
rect 12233 3515 12259 3541
rect 12259 3515 12260 3541
rect 12232 3514 12260 3515
rect 12284 3541 12312 3542
rect 12284 3515 12285 3541
rect 12285 3515 12311 3541
rect 12311 3515 12312 3541
rect 12284 3514 12312 3515
rect 12336 3541 12364 3542
rect 12336 3515 12337 3541
rect 12337 3515 12363 3541
rect 12363 3515 12364 3541
rect 12336 3514 12364 3515
rect 11902 3149 11930 3150
rect 11902 3123 11903 3149
rect 11903 3123 11929 3149
rect 11929 3123 11930 3149
rect 11902 3122 11930 3123
rect 11954 3149 11982 3150
rect 11954 3123 11955 3149
rect 11955 3123 11981 3149
rect 11981 3123 11982 3149
rect 11954 3122 11982 3123
rect 12006 3149 12034 3150
rect 12006 3123 12007 3149
rect 12007 3123 12033 3149
rect 12033 3123 12034 3149
rect 12006 3122 12034 3123
rect 12232 2757 12260 2758
rect 12232 2731 12233 2757
rect 12233 2731 12259 2757
rect 12259 2731 12260 2757
rect 12232 2730 12260 2731
rect 12284 2757 12312 2758
rect 12284 2731 12285 2757
rect 12285 2731 12311 2757
rect 12311 2731 12312 2757
rect 12284 2730 12312 2731
rect 12336 2757 12364 2758
rect 12336 2731 12337 2757
rect 12337 2731 12363 2757
rect 12363 2731 12364 2757
rect 12336 2730 12364 2731
rect 11902 2365 11930 2366
rect 11902 2339 11903 2365
rect 11903 2339 11929 2365
rect 11929 2339 11930 2365
rect 11902 2338 11930 2339
rect 11954 2365 11982 2366
rect 11954 2339 11955 2365
rect 11955 2339 11981 2365
rect 11981 2339 11982 2365
rect 11954 2338 11982 2339
rect 12006 2365 12034 2366
rect 12006 2339 12007 2365
rect 12007 2339 12033 2365
rect 12033 2339 12034 2365
rect 12006 2338 12034 2339
rect 12232 1973 12260 1974
rect 12232 1947 12233 1973
rect 12233 1947 12259 1973
rect 12259 1947 12260 1973
rect 12232 1946 12260 1947
rect 12284 1973 12312 1974
rect 12284 1947 12285 1973
rect 12285 1947 12311 1973
rect 12311 1947 12312 1973
rect 12284 1946 12312 1947
rect 12336 1973 12364 1974
rect 12336 1947 12337 1973
rect 12337 1947 12363 1973
rect 12363 1947 12364 1973
rect 12336 1946 12364 1947
rect 12614 5417 12642 5418
rect 12614 5391 12615 5417
rect 12615 5391 12641 5417
rect 12641 5391 12642 5417
rect 12614 5390 12642 5391
rect 12614 4886 12642 4914
rect 12894 6566 12922 6594
rect 12950 6790 12978 6818
rect 13454 7014 13482 7042
rect 12950 6454 12978 6482
rect 13006 6118 13034 6146
rect 12782 4830 12810 4858
rect 12838 5838 12866 5866
rect 12614 3990 12642 4018
rect 12894 4886 12922 4914
rect 14350 6958 14378 6986
rect 13398 6118 13426 6146
rect 13510 6846 13538 6874
rect 13062 5782 13090 5810
rect 13230 5950 13258 5978
rect 13118 5249 13146 5250
rect 13118 5223 13119 5249
rect 13119 5223 13145 5249
rect 13145 5223 13146 5249
rect 13118 5222 13146 5223
rect 13174 4857 13202 4858
rect 13174 4831 13175 4857
rect 13175 4831 13201 4857
rect 13201 4831 13202 4857
rect 13174 4830 13202 4831
rect 13286 5894 13314 5922
rect 12838 3038 12866 3066
rect 11830 1638 11858 1666
rect 11902 1581 11930 1582
rect 11902 1555 11903 1581
rect 11903 1555 11929 1581
rect 11929 1555 11930 1581
rect 11902 1554 11930 1555
rect 11954 1581 11982 1582
rect 11954 1555 11955 1581
rect 11955 1555 11981 1581
rect 11981 1555 11982 1581
rect 11954 1554 11982 1555
rect 12006 1581 12034 1582
rect 12006 1555 12007 1581
rect 12007 1555 12033 1581
rect 12033 1555 12034 1581
rect 12006 1554 12034 1555
rect 11830 1470 11858 1498
rect 12232 1189 12260 1190
rect 12232 1163 12233 1189
rect 12233 1163 12259 1189
rect 12259 1163 12260 1189
rect 12232 1162 12260 1163
rect 12284 1189 12312 1190
rect 12284 1163 12285 1189
rect 12285 1163 12311 1189
rect 12311 1163 12312 1189
rect 12284 1162 12312 1163
rect 12336 1189 12364 1190
rect 12336 1163 12337 1189
rect 12337 1163 12363 1189
rect 12363 1163 12364 1189
rect 12336 1162 12364 1163
rect 11902 797 11930 798
rect 11902 771 11903 797
rect 11903 771 11929 797
rect 11929 771 11930 797
rect 11902 770 11930 771
rect 11954 797 11982 798
rect 11954 771 11955 797
rect 11955 771 11981 797
rect 11981 771 11982 797
rect 11954 770 11982 771
rect 12006 797 12034 798
rect 12006 771 12007 797
rect 12007 771 12033 797
rect 12033 771 12034 797
rect 12006 770 12034 771
rect 13062 4382 13090 4410
rect 13118 3654 13146 3682
rect 13230 2198 13258 2226
rect 13454 5838 13482 5866
rect 13398 5782 13426 5810
rect 14126 6734 14154 6762
rect 13790 6510 13818 6538
rect 13566 6398 13594 6426
rect 13734 6033 13762 6034
rect 13734 6007 13735 6033
rect 13735 6007 13761 6033
rect 13761 6007 13762 6033
rect 13734 6006 13762 6007
rect 13678 5838 13706 5866
rect 13622 5614 13650 5642
rect 13342 3374 13370 3402
rect 13454 1862 13482 1890
rect 13118 910 13146 938
rect 11774 294 11802 322
rect 11382 238 11410 266
rect 12502 686 12530 714
rect 12166 601 12194 602
rect 12166 575 12167 601
rect 12167 575 12193 601
rect 12193 575 12194 601
rect 12166 574 12194 575
rect 12232 405 12260 406
rect 12232 379 12233 405
rect 12233 379 12259 405
rect 12259 379 12260 405
rect 12232 378 12260 379
rect 12284 405 12312 406
rect 12284 379 12285 405
rect 12285 379 12311 405
rect 12311 379 12312 405
rect 12284 378 12312 379
rect 12336 405 12364 406
rect 12336 379 12337 405
rect 12337 379 12363 405
rect 12363 379 12364 405
rect 12336 378 12364 379
rect 12446 238 12474 266
rect 12950 545 12978 546
rect 12950 519 12951 545
rect 12951 519 12977 545
rect 12977 519 12978 545
rect 12950 518 12978 519
rect 13342 1414 13370 1442
rect 13678 4606 13706 4634
rect 13902 5838 13930 5866
rect 13846 5278 13874 5306
rect 13902 4046 13930 4074
rect 13902 3262 13930 3290
rect 13902 2646 13930 2674
rect 13902 2086 13930 2114
rect 13454 1358 13482 1386
rect 13846 1694 13874 1722
rect 13622 686 13650 714
rect 13342 462 13370 490
rect 14126 6342 14154 6370
rect 14294 5894 14322 5922
rect 14910 6593 14938 6594
rect 14910 6567 14911 6593
rect 14911 6567 14937 6593
rect 14937 6567 14938 6593
rect 14910 6566 14938 6567
rect 14518 6201 14546 6202
rect 14518 6175 14519 6201
rect 14519 6175 14545 6201
rect 14545 6175 14546 6201
rect 14518 6174 14546 6175
rect 14462 5670 14490 5698
rect 14406 5390 14434 5418
rect 14294 5166 14322 5194
rect 14014 3766 14042 3794
rect 14126 2030 14154 2058
rect 13958 1694 13986 1722
rect 13902 1302 13930 1330
rect 13734 70 13762 98
rect 13902 70 13930 98
rect 14070 70 14098 98
rect 10094 14 10122 42
rect 14686 5558 14714 5586
rect 14686 4774 14714 4802
rect 14686 4550 14714 4578
rect 14742 4494 14770 4522
rect 14686 4129 14714 4130
rect 14686 4103 14687 4129
rect 14687 4103 14713 4129
rect 14713 4103 14714 4129
rect 14686 4102 14714 4103
rect 14686 3681 14714 3682
rect 14686 3655 14687 3681
rect 14687 3655 14713 3681
rect 14713 3655 14714 3681
rect 14686 3654 14714 3655
rect 14686 3345 14714 3346
rect 14686 3319 14687 3345
rect 14687 3319 14713 3345
rect 14713 3319 14714 3345
rect 14686 3318 14714 3319
rect 14406 3150 14434 3178
rect 14686 2897 14714 2898
rect 14686 2871 14687 2897
rect 14687 2871 14713 2897
rect 14713 2871 14714 2897
rect 14686 2870 14714 2871
rect 14686 2617 14714 2618
rect 14686 2591 14687 2617
rect 14687 2591 14713 2617
rect 14713 2591 14714 2617
rect 14686 2590 14714 2591
rect 14742 2534 14770 2562
rect 14406 2505 14434 2506
rect 14406 2479 14407 2505
rect 14407 2479 14433 2505
rect 14433 2479 14434 2505
rect 14406 2478 14434 2479
rect 14686 2169 14714 2170
rect 14686 2143 14687 2169
rect 14687 2143 14713 2169
rect 14713 2143 14714 2169
rect 14686 2142 14714 2143
rect 14294 1833 14322 1834
rect 14294 1807 14295 1833
rect 14295 1807 14321 1833
rect 14321 1807 14322 1833
rect 14294 1806 14322 1807
rect 14294 1694 14322 1722
rect 14686 1385 14714 1386
rect 14686 1359 14687 1385
rect 14687 1359 14713 1385
rect 14713 1359 14714 1385
rect 14686 1358 14714 1359
rect 14406 1134 14434 1162
rect 14350 910 14378 938
rect 14686 1078 14714 1106
rect 14742 966 14770 994
rect 15302 5950 15330 5978
rect 15190 4942 15218 4970
rect 15078 4718 15106 4746
rect 15190 4494 15218 4522
rect 15078 4270 15106 4298
rect 15134 4046 15162 4074
rect 15190 3822 15218 3850
rect 15190 3598 15218 3626
rect 15134 3374 15162 3402
rect 15078 2926 15106 2954
rect 15134 2702 15162 2730
rect 15190 2254 15218 2282
rect 15134 2030 15162 2058
rect 15078 1582 15106 1610
rect 15190 1358 15218 1386
rect 15022 630 15050 658
<< metal3 >>
rect 11769 7014 11774 7042
rect 11802 7014 12558 7042
rect 12586 7014 12591 7042
rect 13449 7014 13454 7042
rect 13482 7014 14490 7042
rect 0 6986 56 7000
rect 14462 6986 14490 7014
rect 15792 6986 15848 7000
rect 0 6958 70 6986
rect 98 6958 103 6986
rect 10649 6958 10654 6986
rect 10682 6958 14350 6986
rect 14378 6958 14383 6986
rect 14462 6958 15848 6986
rect 0 6944 56 6958
rect 15792 6944 15848 6958
rect 3313 6902 3318 6930
rect 3346 6902 9422 6930
rect 9450 6902 9455 6930
rect 10593 6902 10598 6930
rect 10626 6902 14322 6930
rect 2417 6846 2422 6874
rect 2450 6846 6734 6874
rect 6762 6846 6767 6874
rect 12329 6846 12334 6874
rect 12362 6846 13510 6874
rect 13538 6846 13543 6874
rect 1857 6790 1862 6818
rect 1890 6790 3822 6818
rect 3850 6790 3855 6818
rect 4881 6790 4886 6818
rect 4914 6790 5838 6818
rect 5866 6790 5871 6818
rect 6561 6790 6566 6818
rect 6594 6790 8414 6818
rect 8442 6790 8447 6818
rect 11545 6790 11550 6818
rect 11578 6790 12950 6818
rect 12978 6790 12983 6818
rect 0 6762 56 6776
rect 14294 6762 14322 6902
rect 15792 6762 15848 6776
rect 0 6734 294 6762
rect 322 6734 327 6762
rect 3761 6734 3766 6762
rect 3794 6734 5054 6762
rect 5082 6734 5087 6762
rect 12217 6734 12222 6762
rect 12250 6734 14126 6762
rect 14154 6734 14159 6762
rect 14294 6734 15848 6762
rect 0 6720 56 6734
rect 15792 6720 15848 6734
rect 4153 6678 4158 6706
rect 4186 6678 5166 6706
rect 5194 6678 5199 6706
rect 2227 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2369 6678
rect 12227 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12369 6678
rect 2977 6622 2982 6650
rect 3010 6622 4382 6650
rect 4410 6622 4415 6650
rect 8129 6622 8134 6650
rect 8162 6622 8638 6650
rect 8666 6622 8671 6650
rect 10985 6622 10990 6650
rect 11018 6622 11382 6650
rect 11410 6622 11415 6650
rect 1073 6566 1078 6594
rect 1106 6566 3150 6594
rect 3178 6566 3183 6594
rect 3257 6566 3262 6594
rect 3290 6566 4214 6594
rect 5665 6566 5670 6594
rect 5698 6566 6286 6594
rect 6314 6566 6319 6594
rect 6617 6566 6622 6594
rect 6650 6566 7014 6594
rect 7042 6566 7047 6594
rect 7849 6566 7854 6594
rect 7882 6566 8526 6594
rect 8554 6566 8559 6594
rect 9193 6566 9198 6594
rect 9226 6566 9478 6594
rect 9506 6566 9511 6594
rect 10873 6566 10878 6594
rect 10906 6566 11270 6594
rect 11298 6566 11303 6594
rect 11881 6566 11886 6594
rect 11914 6566 12166 6594
rect 12194 6566 12199 6594
rect 12889 6566 12894 6594
rect 12922 6566 14910 6594
rect 14938 6566 14943 6594
rect 0 6538 56 6552
rect 4186 6538 4214 6566
rect 15792 6538 15848 6552
rect 0 6510 126 6538
rect 154 6510 159 6538
rect 4186 6510 7574 6538
rect 7602 6510 7607 6538
rect 11097 6510 11102 6538
rect 11130 6510 12222 6538
rect 12250 6510 12255 6538
rect 13785 6510 13790 6538
rect 13818 6510 15848 6538
rect 0 6496 56 6510
rect 15792 6496 15848 6510
rect 5945 6454 5950 6482
rect 5978 6454 10038 6482
rect 10066 6454 10071 6482
rect 11657 6454 11662 6482
rect 11690 6454 12950 6482
rect 12978 6454 12983 6482
rect 7121 6398 7126 6426
rect 7154 6398 9702 6426
rect 9730 6398 9735 6426
rect 11993 6398 11998 6426
rect 12026 6398 13566 6426
rect 13594 6398 13599 6426
rect 4769 6342 4774 6370
rect 4802 6342 7742 6370
rect 7770 6342 7775 6370
rect 11769 6342 11774 6370
rect 11802 6342 11942 6370
rect 11970 6342 11975 6370
rect 12553 6342 12558 6370
rect 12586 6342 14126 6370
rect 14154 6342 14159 6370
rect 0 6314 56 6328
rect 15792 6314 15848 6328
rect 0 6286 1246 6314
rect 1274 6286 1279 6314
rect 5217 6286 5222 6314
rect 5250 6286 7294 6314
rect 7322 6286 7327 6314
rect 12721 6286 12726 6314
rect 12754 6286 15848 6314
rect 0 6272 56 6286
rect 1897 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2039 6286
rect 11897 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12039 6286
rect 15792 6272 15848 6286
rect 2753 6230 2758 6258
rect 2786 6230 3150 6258
rect 3178 6230 3183 6258
rect 5161 6230 5166 6258
rect 5194 6230 8806 6258
rect 8834 6230 8839 6258
rect 2529 6174 2534 6202
rect 2562 6174 2926 6202
rect 2954 6174 2959 6202
rect 3649 6174 3654 6202
rect 3682 6174 4718 6202
rect 4746 6174 4751 6202
rect 5049 6174 5054 6202
rect 5082 6174 5614 6202
rect 5642 6174 5647 6202
rect 6001 6174 6006 6202
rect 6034 6174 6174 6202
rect 6202 6174 6207 6202
rect 6505 6174 6510 6202
rect 6538 6174 6734 6202
rect 6762 6174 6767 6202
rect 7126 6174 8190 6202
rect 8218 6174 8223 6202
rect 11321 6174 11326 6202
rect 11354 6174 11998 6202
rect 12026 6174 12031 6202
rect 12665 6174 12670 6202
rect 12698 6174 14518 6202
rect 14546 6174 14551 6202
rect 1913 6118 1918 6146
rect 1946 6118 3374 6146
rect 3402 6118 3407 6146
rect 5161 6118 5166 6146
rect 5194 6118 5502 6146
rect 5530 6118 5535 6146
rect 0 6090 56 6104
rect 7126 6090 7154 6174
rect 7681 6118 7686 6146
rect 7714 6118 8302 6146
rect 8330 6118 8335 6146
rect 13001 6118 13006 6146
rect 13034 6118 13398 6146
rect 13426 6118 13431 6146
rect 15792 6090 15848 6104
rect 0 6062 182 6090
rect 210 6062 215 6090
rect 2641 6062 2646 6090
rect 2674 6062 3598 6090
rect 3626 6062 3631 6090
rect 4433 6062 4438 6090
rect 4466 6062 7154 6090
rect 7233 6062 7238 6090
rect 7266 6062 8862 6090
rect 8890 6062 8895 6090
rect 9305 6062 9310 6090
rect 9338 6062 9758 6090
rect 9786 6062 9791 6090
rect 10481 6062 10486 6090
rect 10514 6062 15848 6090
rect 0 6048 56 6062
rect 15792 6048 15848 6062
rect 2193 6006 2198 6034
rect 2226 6006 4494 6034
rect 4522 6006 4527 6034
rect 5329 6006 5334 6034
rect 5362 6006 9814 6034
rect 9842 6006 9847 6034
rect 9921 6006 9926 6034
rect 9954 6006 11102 6034
rect 11130 6006 11135 6034
rect 12497 6006 12502 6034
rect 12530 6006 13734 6034
rect 13762 6006 13767 6034
rect 3089 5950 3094 5978
rect 3122 5950 3486 5978
rect 3514 5950 3519 5978
rect 3593 5950 3598 5978
rect 3626 5950 5502 5978
rect 5530 5950 5535 5978
rect 6001 5950 6006 5978
rect 6034 5950 7518 5978
rect 7546 5950 7551 5978
rect 10537 5950 10542 5978
rect 10570 5950 12194 5978
rect 13225 5950 13230 5978
rect 13258 5950 15302 5978
rect 15330 5950 15335 5978
rect 2977 5894 2982 5922
rect 3010 5894 4438 5922
rect 4466 5894 4471 5922
rect 4545 5894 4550 5922
rect 4578 5894 7406 5922
rect 7434 5894 7439 5922
rect 9585 5894 9590 5922
rect 9618 5894 10990 5922
rect 11018 5894 11023 5922
rect 0 5866 56 5880
rect 2227 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2369 5894
rect 0 5838 910 5866
rect 938 5838 943 5866
rect 3873 5838 3878 5866
rect 3906 5838 4438 5866
rect 4466 5838 4471 5866
rect 0 5824 56 5838
rect 12166 5810 12194 5950
rect 13281 5894 13286 5922
rect 13314 5894 14294 5922
rect 14322 5894 14327 5922
rect 12227 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12369 5894
rect 15792 5866 15848 5880
rect 12665 5838 12670 5866
rect 12698 5838 12838 5866
rect 12866 5838 12871 5866
rect 13449 5838 13454 5866
rect 13482 5838 13678 5866
rect 13706 5838 13711 5866
rect 13897 5838 13902 5866
rect 13930 5838 15848 5866
rect 15792 5824 15848 5838
rect 1521 5782 1526 5810
rect 1554 5782 9562 5810
rect 11209 5782 11214 5810
rect 11242 5782 11606 5810
rect 11634 5782 11639 5810
rect 12166 5782 12222 5810
rect 12250 5782 12255 5810
rect 13057 5782 13062 5810
rect 13090 5782 13398 5810
rect 13426 5782 13431 5810
rect 9534 5754 9562 5782
rect 2305 5726 2310 5754
rect 2338 5726 3206 5754
rect 3234 5726 3239 5754
rect 5217 5726 5222 5754
rect 5250 5726 8078 5754
rect 8106 5726 8111 5754
rect 9534 5726 11550 5754
rect 11578 5726 11583 5754
rect 2977 5670 2982 5698
rect 3010 5670 3822 5698
rect 3850 5670 3855 5698
rect 4153 5670 4158 5698
rect 4186 5670 6286 5698
rect 6314 5670 6319 5698
rect 8689 5670 8694 5698
rect 8722 5670 14462 5698
rect 14490 5670 14495 5698
rect 0 5642 56 5656
rect 15792 5642 15848 5656
rect 0 5614 406 5642
rect 434 5614 439 5642
rect 5665 5614 5670 5642
rect 5698 5614 7182 5642
rect 7210 5614 7215 5642
rect 7905 5614 7910 5642
rect 7938 5614 8974 5642
rect 9002 5614 9007 5642
rect 9529 5614 9534 5642
rect 9562 5614 9870 5642
rect 9898 5614 9903 5642
rect 12539 5614 12558 5642
rect 12586 5614 12591 5642
rect 13617 5614 13622 5642
rect 13650 5614 15848 5642
rect 0 5600 56 5614
rect 15792 5600 15848 5614
rect 4713 5558 4718 5586
rect 4746 5558 8750 5586
rect 8778 5558 8783 5586
rect 10761 5558 10766 5586
rect 10794 5558 14686 5586
rect 14714 5558 14719 5586
rect 7009 5502 7014 5530
rect 7042 5502 9254 5530
rect 9282 5502 9287 5530
rect 10201 5502 10206 5530
rect 10234 5502 10710 5530
rect 10738 5502 10743 5530
rect 1897 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2039 5502
rect 11897 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12039 5502
rect 4153 5446 4158 5474
rect 4186 5446 5222 5474
rect 5250 5446 5255 5474
rect 5329 5446 5334 5474
rect 5362 5446 11382 5474
rect 11410 5446 11415 5474
rect 12105 5446 12110 5474
rect 12138 5446 12558 5474
rect 12586 5446 12591 5474
rect 0 5418 56 5432
rect 15792 5418 15848 5432
rect 0 5390 1078 5418
rect 1106 5390 1111 5418
rect 1913 5390 1918 5418
rect 1946 5390 2702 5418
rect 2730 5390 2735 5418
rect 3481 5390 3486 5418
rect 3514 5390 4046 5418
rect 4074 5390 4079 5418
rect 4265 5390 4270 5418
rect 4298 5390 4718 5418
rect 4746 5390 4751 5418
rect 5889 5390 5894 5418
rect 5922 5390 6566 5418
rect 6594 5390 6599 5418
rect 9865 5390 9870 5418
rect 9898 5390 11242 5418
rect 11433 5390 11438 5418
rect 11466 5390 11830 5418
rect 11858 5390 11863 5418
rect 12161 5390 12166 5418
rect 12194 5390 12614 5418
rect 12642 5390 12647 5418
rect 14401 5390 14406 5418
rect 14434 5390 15848 5418
rect 0 5376 56 5390
rect 11214 5362 11242 5390
rect 15792 5376 15848 5390
rect 1353 5334 1358 5362
rect 1386 5334 7182 5362
rect 7210 5334 7215 5362
rect 7457 5334 7462 5362
rect 7490 5334 7966 5362
rect 7994 5334 7999 5362
rect 10313 5334 10318 5362
rect 10346 5334 11102 5362
rect 11130 5334 11135 5362
rect 11214 5334 12278 5362
rect 12306 5334 12311 5362
rect 2977 5278 2982 5306
rect 3010 5278 3318 5306
rect 3346 5278 3351 5306
rect 3761 5278 3766 5306
rect 3794 5278 4718 5306
rect 4746 5278 4751 5306
rect 4825 5278 4830 5306
rect 4858 5278 5222 5306
rect 5250 5278 5255 5306
rect 9081 5278 9086 5306
rect 9114 5278 9702 5306
rect 9730 5278 9735 5306
rect 11153 5278 11158 5306
rect 11186 5278 13846 5306
rect 13874 5278 13879 5306
rect 2137 5222 2142 5250
rect 2170 5222 5166 5250
rect 5194 5222 5199 5250
rect 6113 5222 6118 5250
rect 6146 5222 9254 5250
rect 9282 5222 9287 5250
rect 10145 5222 10150 5250
rect 10178 5222 10654 5250
rect 10682 5222 10687 5250
rect 12441 5222 12446 5250
rect 12474 5222 13118 5250
rect 13146 5222 13151 5250
rect 0 5194 56 5208
rect 15792 5194 15848 5208
rect 0 5166 826 5194
rect 7177 5166 7182 5194
rect 7210 5166 7742 5194
rect 7770 5166 7775 5194
rect 9081 5166 9086 5194
rect 9114 5166 12334 5194
rect 12362 5166 12367 5194
rect 14289 5166 14294 5194
rect 14322 5166 15848 5194
rect 0 5152 56 5166
rect 798 5026 826 5166
rect 15792 5152 15848 5166
rect 5777 5110 5782 5138
rect 5810 5110 8134 5138
rect 8162 5110 8167 5138
rect 10369 5110 10374 5138
rect 10402 5110 11550 5138
rect 11578 5110 11583 5138
rect 2227 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2369 5110
rect 12227 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12369 5110
rect 5833 5054 5838 5082
rect 5866 5054 7686 5082
rect 7714 5054 7719 5082
rect 798 4998 4270 5026
rect 4298 4998 4303 5026
rect 5329 4998 5334 5026
rect 5362 4998 8694 5026
rect 8722 4998 8727 5026
rect 10089 4998 10094 5026
rect 10122 4998 10542 5026
rect 10570 4998 10575 5026
rect 0 4970 56 4984
rect 15792 4970 15848 4984
rect 0 4942 4214 4970
rect 4242 4942 4247 4970
rect 5553 4942 5558 4970
rect 5586 4942 10822 4970
rect 10850 4942 10855 4970
rect 11755 4942 11774 4970
rect 11802 4942 11807 4970
rect 15185 4942 15190 4970
rect 15218 4942 15848 4970
rect 0 4928 56 4942
rect 15792 4928 15848 4942
rect 2025 4886 2030 4914
rect 2058 4886 2422 4914
rect 2450 4886 2455 4914
rect 4153 4886 4158 4914
rect 0 4746 56 4760
rect 4186 4746 4214 4914
rect 6113 4886 6118 4914
rect 6146 4886 10934 4914
rect 10962 4886 10967 4914
rect 11657 4886 11662 4914
rect 11690 4886 12278 4914
rect 12306 4886 12311 4914
rect 12609 4886 12614 4914
rect 12642 4886 12894 4914
rect 12922 4886 12927 4914
rect 6673 4830 6678 4858
rect 6706 4830 7882 4858
rect 7961 4830 7966 4858
rect 7994 4830 12334 4858
rect 12362 4830 12367 4858
rect 12777 4830 12782 4858
rect 12810 4830 13174 4858
rect 13202 4830 13207 4858
rect 7854 4746 7882 4830
rect 9142 4774 14686 4802
rect 14714 4774 14719 4802
rect 0 4718 1834 4746
rect 4186 4718 7574 4746
rect 7602 4718 7607 4746
rect 7854 4718 9030 4746
rect 9058 4718 9063 4746
rect 0 4704 56 4718
rect 1806 4634 1834 4718
rect 1897 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2039 4718
rect 9142 4690 9170 4774
rect 15792 4746 15848 4760
rect 15073 4718 15078 4746
rect 15106 4718 15848 4746
rect 11897 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12039 4718
rect 15792 4704 15848 4718
rect 2585 4662 2590 4690
rect 2618 4662 6902 4690
rect 6930 4662 6935 4690
rect 7849 4662 7854 4690
rect 7882 4662 9170 4690
rect 1806 4606 2534 4634
rect 2562 4606 2567 4634
rect 4769 4606 4774 4634
rect 4802 4606 7798 4634
rect 7826 4606 7831 4634
rect 8353 4606 8358 4634
rect 8386 4606 11858 4634
rect 11937 4606 11942 4634
rect 11970 4606 13678 4634
rect 13706 4606 13711 4634
rect 11830 4578 11858 4606
rect 4097 4550 4102 4578
rect 4130 4550 5726 4578
rect 5754 4550 5759 4578
rect 7569 4550 7574 4578
rect 7602 4550 8302 4578
rect 8330 4550 8335 4578
rect 10873 4550 10878 4578
rect 10906 4550 11718 4578
rect 11746 4550 11751 4578
rect 11830 4550 14686 4578
rect 14714 4550 14719 4578
rect 0 4522 56 4536
rect 15792 4522 15848 4536
rect 0 4494 5838 4522
rect 5866 4494 5871 4522
rect 6225 4494 6230 4522
rect 6258 4494 7574 4522
rect 7602 4494 7607 4522
rect 7905 4494 7910 4522
rect 7938 4494 12222 4522
rect 12250 4494 12255 4522
rect 12329 4494 12334 4522
rect 12362 4494 14742 4522
rect 14770 4494 14775 4522
rect 15185 4494 15190 4522
rect 15218 4494 15848 4522
rect 0 4480 56 4494
rect 15792 4480 15848 4494
rect 1857 4438 1862 4466
rect 1890 4438 2590 4466
rect 2618 4438 2623 4466
rect 4657 4438 4662 4466
rect 4690 4438 11886 4466
rect 11914 4438 11919 4466
rect 2086 4382 2450 4410
rect 2529 4382 2534 4410
rect 2562 4382 7574 4410
rect 7602 4382 7607 4410
rect 9193 4382 9198 4410
rect 9226 4382 11494 4410
rect 11522 4382 11527 4410
rect 11718 4382 13062 4410
rect 13090 4382 13095 4410
rect 0 4298 56 4312
rect 2086 4298 2114 4382
rect 2422 4354 2450 4382
rect 11718 4354 11746 4382
rect 2422 4326 5782 4354
rect 5810 4326 5815 4354
rect 10705 4326 10710 4354
rect 10738 4326 11746 4354
rect 2227 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2369 4326
rect 12227 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12369 4326
rect 15792 4298 15848 4312
rect 0 4270 2114 4298
rect 4153 4270 4158 4298
rect 4186 4270 5726 4298
rect 5754 4270 5759 4298
rect 9361 4270 9366 4298
rect 9394 4270 11942 4298
rect 11970 4270 11975 4298
rect 15073 4270 15078 4298
rect 15106 4270 15848 4298
rect 0 4256 56 4270
rect 15792 4256 15848 4270
rect 3257 4214 3262 4242
rect 3290 4214 5502 4242
rect 5530 4214 5535 4242
rect 10033 4214 10038 4242
rect 10066 4214 12334 4242
rect 12362 4214 12367 4242
rect 2025 4158 2030 4186
rect 2058 4158 4438 4186
rect 4466 4158 4471 4186
rect 5273 4158 5278 4186
rect 5306 4158 7350 4186
rect 7378 4158 7383 4186
rect 4713 4102 4718 4130
rect 4746 4102 7070 4130
rect 7098 4102 7103 4130
rect 8465 4102 8470 4130
rect 8498 4102 14686 4130
rect 14714 4102 14719 4130
rect 0 4074 56 4088
rect 15792 4074 15848 4088
rect 0 4046 686 4074
rect 714 4046 719 4074
rect 3985 4046 3990 4074
rect 4018 4046 5054 4074
rect 5082 4046 5087 4074
rect 9137 4046 9142 4074
rect 9170 4046 13902 4074
rect 13930 4046 13935 4074
rect 15129 4046 15134 4074
rect 15162 4046 15848 4074
rect 0 4032 56 4046
rect 15792 4032 15848 4046
rect 3313 3990 3318 4018
rect 3346 3990 5950 4018
rect 5978 3990 5983 4018
rect 7737 3990 7742 4018
rect 7770 3990 12614 4018
rect 12642 3990 12647 4018
rect 2585 3934 2590 3962
rect 2618 3934 6846 3962
rect 6874 3934 6879 3962
rect 1897 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2039 3934
rect 11897 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12039 3934
rect 8073 3878 8078 3906
rect 8106 3878 10766 3906
rect 10794 3878 10799 3906
rect 0 3850 56 3864
rect 15792 3850 15848 3864
rect 0 3822 8190 3850
rect 8218 3822 8223 3850
rect 15185 3822 15190 3850
rect 15218 3822 15848 3850
rect 0 3808 56 3822
rect 15792 3808 15848 3822
rect 7513 3766 7518 3794
rect 7546 3766 14014 3794
rect 14042 3766 14047 3794
rect 4209 3710 4214 3738
rect 4242 3710 7798 3738
rect 7826 3710 7831 3738
rect 8969 3710 8974 3738
rect 9002 3710 13454 3738
rect 13426 3682 13454 3710
rect 401 3654 406 3682
rect 434 3654 3374 3682
rect 3402 3654 3407 3682
rect 3705 3654 3710 3682
rect 3738 3654 6958 3682
rect 6986 3654 6991 3682
rect 11601 3654 11606 3682
rect 11634 3654 13118 3682
rect 13146 3654 13151 3682
rect 13426 3654 14686 3682
rect 14714 3654 14719 3682
rect 0 3626 56 3640
rect 15792 3626 15848 3640
rect 0 3598 2170 3626
rect 4321 3598 4326 3626
rect 4354 3598 9422 3626
rect 9450 3598 9455 3626
rect 15185 3598 15190 3626
rect 15218 3598 15848 3626
rect 0 3584 56 3598
rect 2142 3458 2170 3598
rect 15792 3584 15848 3598
rect 2227 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2369 3542
rect 12227 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12369 3542
rect 3873 3486 3878 3514
rect 3906 3486 4942 3514
rect 4970 3486 4975 3514
rect 6729 3486 6734 3514
rect 6762 3486 9870 3514
rect 9898 3486 9903 3514
rect 2142 3430 7854 3458
rect 7882 3430 7887 3458
rect 0 3402 56 3416
rect 15792 3402 15848 3416
rect 0 3374 7350 3402
rect 7378 3374 7383 3402
rect 8913 3374 8918 3402
rect 8946 3374 13342 3402
rect 13370 3374 13375 3402
rect 15129 3374 15134 3402
rect 15162 3374 15848 3402
rect 0 3360 56 3374
rect 15792 3360 15848 3374
rect 3817 3318 3822 3346
rect 3850 3318 7910 3346
rect 7938 3318 7943 3346
rect 8017 3318 8022 3346
rect 8050 3318 14686 3346
rect 14714 3318 14719 3346
rect 126 3262 7182 3290
rect 7210 3262 7215 3290
rect 7457 3262 7462 3290
rect 7490 3262 13902 3290
rect 13930 3262 13935 3290
rect 0 3178 56 3192
rect 126 3178 154 3262
rect 233 3206 238 3234
rect 266 3206 9198 3234
rect 9226 3206 9231 3234
rect 15792 3178 15848 3192
rect 0 3150 154 3178
rect 14401 3150 14406 3178
rect 14434 3150 15848 3178
rect 0 3136 56 3150
rect 1897 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2039 3150
rect 11897 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12039 3150
rect 15792 3136 15848 3150
rect 4186 3094 7574 3122
rect 7602 3094 7607 3122
rect 4186 3066 4214 3094
rect 681 3038 686 3066
rect 714 3038 4214 3066
rect 4265 3038 4270 3066
rect 4298 3038 7238 3066
rect 7266 3038 7271 3066
rect 8297 3038 8302 3066
rect 8330 3038 12838 3066
rect 12866 3038 12871 3066
rect 1073 2982 1078 3010
rect 1106 2982 8862 3010
rect 8890 2982 8895 3010
rect 0 2954 56 2968
rect 15792 2954 15848 2968
rect 0 2926 7182 2954
rect 7210 2926 7215 2954
rect 15073 2926 15078 2954
rect 15106 2926 15848 2954
rect 0 2912 56 2926
rect 15792 2912 15848 2926
rect 7625 2870 7630 2898
rect 7658 2870 14686 2898
rect 14714 2870 14719 2898
rect 0 2730 56 2744
rect 2227 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2369 2758
rect 12227 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12369 2758
rect 15792 2730 15848 2744
rect 0 2702 2114 2730
rect 15129 2702 15134 2730
rect 15162 2702 15848 2730
rect 0 2688 56 2702
rect 2086 2674 2114 2702
rect 15792 2688 15848 2702
rect 2086 2646 8414 2674
rect 8442 2646 8447 2674
rect 8689 2646 8694 2674
rect 8722 2646 13902 2674
rect 13930 2646 13935 2674
rect 7513 2590 7518 2618
rect 7546 2590 14686 2618
rect 14714 2590 14719 2618
rect 8073 2534 8078 2562
rect 8106 2534 14742 2562
rect 14770 2534 14775 2562
rect 0 2506 56 2520
rect 15792 2506 15848 2520
rect 0 2478 8414 2506
rect 8442 2478 8447 2506
rect 14401 2478 14406 2506
rect 14434 2478 15848 2506
rect 0 2464 56 2478
rect 15792 2464 15848 2478
rect 289 2422 294 2450
rect 322 2422 10206 2450
rect 10234 2422 10239 2450
rect 1897 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2039 2366
rect 11897 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12039 2366
rect 0 2282 56 2296
rect 15792 2282 15848 2296
rect 0 2254 7798 2282
rect 7826 2254 7831 2282
rect 15185 2254 15190 2282
rect 15218 2254 15848 2282
rect 0 2240 56 2254
rect 15792 2240 15848 2254
rect 8129 2198 8134 2226
rect 8162 2198 13230 2226
rect 13258 2198 13263 2226
rect 8633 2142 8638 2170
rect 8666 2142 14686 2170
rect 14714 2142 14719 2170
rect 7513 2086 7518 2114
rect 7546 2086 13902 2114
rect 13930 2086 13935 2114
rect 0 2058 56 2072
rect 15792 2058 15848 2072
rect 0 2030 6790 2058
rect 6818 2030 6823 2058
rect 10761 2030 10766 2058
rect 10794 2030 14126 2058
rect 14154 2030 14159 2058
rect 15129 2030 15134 2058
rect 15162 2030 15848 2058
rect 0 2016 56 2030
rect 15792 2016 15848 2030
rect 3369 1974 3374 2002
rect 3402 1974 7854 2002
rect 7882 1974 7887 2002
rect 2227 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2369 1974
rect 12227 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12369 1974
rect 4186 1918 8638 1946
rect 8666 1918 8671 1946
rect 4186 1890 4214 1918
rect 905 1862 910 1890
rect 938 1862 4214 1890
rect 7065 1862 7070 1890
rect 7098 1862 13454 1890
rect 13482 1862 13487 1890
rect 0 1834 56 1848
rect 15792 1834 15848 1848
rect 0 1806 7294 1834
rect 7322 1806 7327 1834
rect 14289 1806 14294 1834
rect 14322 1806 15848 1834
rect 0 1792 56 1806
rect 15792 1792 15848 1806
rect 1241 1750 1246 1778
rect 1274 1750 9758 1778
rect 9786 1750 9791 1778
rect 7233 1694 7238 1722
rect 7266 1694 13846 1722
rect 13874 1694 13879 1722
rect 13953 1694 13958 1722
rect 13986 1694 14294 1722
rect 14322 1694 14327 1722
rect 121 1638 126 1666
rect 154 1638 10262 1666
rect 10290 1638 10295 1666
rect 10649 1638 10654 1666
rect 10682 1638 11830 1666
rect 11858 1638 11863 1666
rect 0 1610 56 1624
rect 15792 1610 15848 1624
rect 0 1582 1834 1610
rect 15073 1582 15078 1610
rect 15106 1582 15848 1610
rect 0 1568 56 1582
rect 1806 1442 1834 1582
rect 1897 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2039 1582
rect 11897 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12039 1582
rect 15792 1568 15848 1582
rect 1913 1470 1918 1498
rect 1946 1470 9310 1498
rect 9338 1470 9343 1498
rect 11377 1470 11382 1498
rect 11410 1470 11830 1498
rect 11858 1470 11863 1498
rect 1806 1414 7014 1442
rect 7042 1414 7047 1442
rect 7401 1414 7406 1442
rect 7434 1414 13342 1442
rect 13370 1414 13375 1442
rect 0 1386 56 1400
rect 15792 1386 15848 1400
rect 0 1358 7686 1386
rect 7714 1358 7719 1386
rect 13449 1358 13454 1386
rect 13482 1358 14686 1386
rect 14714 1358 14719 1386
rect 15185 1358 15190 1386
rect 15218 1358 15848 1386
rect 0 1344 56 1358
rect 15792 1344 15848 1358
rect 8353 1302 8358 1330
rect 8386 1302 13902 1330
rect 13930 1302 13935 1330
rect 2086 1246 8134 1274
rect 8162 1246 8167 1274
rect 0 1162 56 1176
rect 2086 1162 2114 1246
rect 7289 1190 7294 1218
rect 7322 1190 11970 1218
rect 2227 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2369 1190
rect 0 1134 2114 1162
rect 0 1120 56 1134
rect 11942 1106 11970 1190
rect 12227 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12369 1190
rect 15792 1162 15848 1176
rect 14401 1134 14406 1162
rect 14434 1134 15848 1162
rect 15792 1120 15848 1134
rect 4186 1078 6958 1106
rect 6986 1078 6991 1106
rect 7961 1078 7966 1106
rect 7994 1078 11914 1106
rect 11942 1078 14686 1106
rect 14714 1078 14719 1106
rect 4186 1050 4214 1078
rect 2086 1022 4214 1050
rect 8073 1022 8078 1050
rect 8106 1022 11634 1050
rect 0 938 56 952
rect 2086 938 2114 1022
rect 2473 966 2478 994
rect 2506 966 9814 994
rect 9842 966 9847 994
rect 10066 966 11326 994
rect 11354 966 11359 994
rect 10066 938 10094 966
rect 0 910 2114 938
rect 6001 910 6006 938
rect 6034 910 7798 938
rect 7826 910 7831 938
rect 8521 910 8526 938
rect 8554 910 10094 938
rect 11606 938 11634 1022
rect 11886 994 11914 1078
rect 11886 966 14742 994
rect 14770 966 14775 994
rect 15792 938 15848 952
rect 11606 910 13118 938
rect 13146 910 13151 938
rect 14345 910 14350 938
rect 14378 910 15848 938
rect 0 896 56 910
rect 15792 896 15848 910
rect 1806 854 2114 882
rect 3817 854 3822 882
rect 3850 854 10822 882
rect 10850 854 10855 882
rect 1806 826 1834 854
rect 65 798 70 826
rect 98 798 1834 826
rect 2086 826 2114 854
rect 2086 798 10094 826
rect 1897 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2039 798
rect 5553 742 5558 770
rect 5586 742 7742 770
rect 7770 742 7775 770
rect 0 714 56 728
rect 0 686 6006 714
rect 6034 686 6039 714
rect 0 672 56 686
rect 10066 658 10094 798
rect 11897 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12039 798
rect 15792 714 15848 728
rect 11209 686 11214 714
rect 11242 686 12502 714
rect 12530 686 12535 714
rect 13617 686 13622 714
rect 13650 686 15848 714
rect 15792 672 15848 686
rect 1745 630 1750 658
rect 1778 630 5166 658
rect 5194 630 5199 658
rect 6561 630 6566 658
rect 6594 630 8302 658
rect 8330 630 8335 658
rect 10066 630 15022 658
rect 15050 630 15055 658
rect 7849 574 7854 602
rect 7882 574 12166 602
rect 12194 574 12199 602
rect 8353 518 8358 546
rect 8386 518 12950 546
rect 12978 518 12983 546
rect 0 490 56 504
rect 15792 490 15848 504
rect 0 462 8134 490
rect 8162 462 8167 490
rect 9865 462 9870 490
rect 9898 462 10542 490
rect 10570 462 10575 490
rect 13337 462 13342 490
rect 13370 462 15848 490
rect 0 448 56 462
rect 15792 448 15848 462
rect 4489 406 4494 434
rect 4522 406 9366 434
rect 9394 406 9399 434
rect 2227 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2369 406
rect 12227 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12369 406
rect 10537 294 10542 322
rect 10570 294 11774 322
rect 11802 294 11807 322
rect 0 266 56 280
rect 15792 266 15848 280
rect 0 238 7574 266
rect 7602 238 7607 266
rect 9193 238 9198 266
rect 9226 238 11382 266
rect 11410 238 11415 266
rect 12441 238 12446 266
rect 12474 238 15848 266
rect 0 224 56 238
rect 15792 224 15848 238
rect 4186 182 7126 210
rect 7154 182 7159 210
rect 7849 182 7854 210
rect 7882 182 8918 210
rect 8946 182 8951 210
rect 4186 154 4214 182
rect 1022 126 4214 154
rect 0 42 56 56
rect 1022 42 1050 126
rect 1129 70 1134 98
rect 1162 70 1167 98
rect 3145 70 3150 98
rect 3178 70 10374 98
rect 10402 70 10407 98
rect 13729 70 13734 98
rect 13762 70 13767 98
rect 13897 70 13902 98
rect 13930 70 14070 98
rect 14098 70 14103 98
rect 0 14 1050 42
rect 1134 42 1162 70
rect 13734 42 13762 70
rect 15792 42 15848 56
rect 1134 14 10094 42
rect 10122 14 10127 42
rect 13734 14 15848 42
rect 0 0 56 14
rect 15792 0 15848 14
<< via3 >>
rect 12558 7014 12586 7042
rect 2232 6650 2260 6678
rect 2284 6650 2312 6678
rect 2336 6650 2364 6678
rect 12232 6650 12260 6678
rect 12284 6650 12312 6678
rect 12336 6650 12364 6678
rect 11774 6342 11802 6370
rect 1902 6258 1930 6286
rect 1954 6258 1982 6286
rect 2006 6258 2034 6286
rect 11902 6258 11930 6286
rect 11954 6258 11982 6286
rect 12006 6258 12034 6286
rect 3598 6062 3626 6090
rect 4438 6062 4466 6090
rect 3598 5950 3626 5978
rect 4438 5894 4466 5922
rect 2232 5866 2260 5894
rect 2284 5866 2312 5894
rect 2336 5866 2364 5894
rect 12232 5866 12260 5894
rect 12284 5866 12312 5894
rect 12336 5866 12364 5894
rect 5222 5726 5250 5754
rect 12558 5614 12586 5642
rect 4718 5558 4746 5586
rect 1902 5474 1930 5502
rect 1954 5474 1982 5502
rect 2006 5474 2034 5502
rect 11902 5474 11930 5502
rect 11954 5474 11982 5502
rect 12006 5474 12034 5502
rect 5222 5446 5250 5474
rect 4718 5278 4746 5306
rect 2232 5082 2260 5110
rect 2284 5082 2312 5110
rect 2336 5082 2364 5110
rect 12232 5082 12260 5110
rect 12284 5082 12312 5110
rect 12336 5082 12364 5110
rect 11774 4942 11802 4970
rect 7574 4718 7602 4746
rect 1902 4690 1930 4718
rect 1954 4690 1982 4718
rect 2006 4690 2034 4718
rect 11902 4690 11930 4718
rect 11954 4690 11982 4718
rect 12006 4690 12034 4718
rect 2534 4606 2562 4634
rect 7574 4550 7602 4578
rect 2534 4382 2562 4410
rect 2232 4298 2260 4326
rect 2284 4298 2312 4326
rect 2336 4298 2364 4326
rect 12232 4298 12260 4326
rect 12284 4298 12312 4326
rect 12336 4298 12364 4326
rect 1902 3906 1930 3934
rect 1954 3906 1982 3934
rect 2006 3906 2034 3934
rect 11902 3906 11930 3934
rect 11954 3906 11982 3934
rect 12006 3906 12034 3934
rect 2232 3514 2260 3542
rect 2284 3514 2312 3542
rect 2336 3514 2364 3542
rect 12232 3514 12260 3542
rect 12284 3514 12312 3542
rect 12336 3514 12364 3542
rect 1902 3122 1930 3150
rect 1954 3122 1982 3150
rect 2006 3122 2034 3150
rect 11902 3122 11930 3150
rect 11954 3122 11982 3150
rect 12006 3122 12034 3150
rect 2232 2730 2260 2758
rect 2284 2730 2312 2758
rect 2336 2730 2364 2758
rect 12232 2730 12260 2758
rect 12284 2730 12312 2758
rect 12336 2730 12364 2758
rect 1902 2338 1930 2366
rect 1954 2338 1982 2366
rect 2006 2338 2034 2366
rect 11902 2338 11930 2366
rect 11954 2338 11982 2366
rect 12006 2338 12034 2366
rect 2232 1946 2260 1974
rect 2284 1946 2312 1974
rect 2336 1946 2364 1974
rect 12232 1946 12260 1974
rect 12284 1946 12312 1974
rect 12336 1946 12364 1974
rect 1902 1554 1930 1582
rect 1954 1554 1982 1582
rect 2006 1554 2034 1582
rect 11902 1554 11930 1582
rect 11954 1554 11982 1582
rect 12006 1554 12034 1582
rect 2232 1162 2260 1190
rect 2284 1162 2312 1190
rect 2336 1162 2364 1190
rect 12232 1162 12260 1190
rect 12284 1162 12312 1190
rect 12336 1162 12364 1190
rect 6006 910 6034 938
rect 1902 770 1930 798
rect 1954 770 1982 798
rect 2006 770 2034 798
rect 6006 686 6034 714
rect 11902 770 11930 798
rect 11954 770 11982 798
rect 12006 770 12034 798
rect 2232 378 2260 406
rect 2284 378 2312 406
rect 2336 378 2364 406
rect 12232 378 12260 406
rect 12284 378 12312 406
rect 12336 378 12364 406
<< metal4 >>
rect 1888 6286 2048 7112
rect 1888 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2048 6286
rect 1888 5502 2048 6258
rect 1888 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2048 5502
rect 1888 4718 2048 5474
rect 1888 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2048 4718
rect 1888 3934 2048 4690
rect 1888 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2048 3934
rect 1888 3150 2048 3906
rect 1888 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2048 3150
rect 1888 2366 2048 3122
rect 1888 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2048 2366
rect 1888 1582 2048 2338
rect 1888 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2048 1582
rect 1888 798 2048 1554
rect 1888 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2048 798
rect 1888 0 2048 770
rect 2218 6678 2378 7112
rect 2218 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2378 6678
rect 2218 5894 2378 6650
rect 11774 6370 11802 6375
rect 3598 6090 3626 6095
rect 3598 5978 3626 6062
rect 3598 5945 3626 5950
rect 4438 6090 4466 6095
rect 2218 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2378 5894
rect 4438 5922 4466 6062
rect 4438 5889 4466 5894
rect 2218 5110 2378 5866
rect 5222 5754 5250 5759
rect 4718 5586 4746 5591
rect 4718 5306 4746 5558
rect 5222 5474 5250 5726
rect 5222 5441 5250 5446
rect 4718 5273 4746 5278
rect 2218 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2378 5110
rect 2218 4326 2378 5082
rect 11774 4970 11802 6342
rect 11774 4937 11802 4942
rect 11888 6286 12048 7112
rect 11888 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12048 6286
rect 11888 5502 12048 6258
rect 11888 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12048 5502
rect 7574 4746 7602 4751
rect 2534 4634 2562 4639
rect 2534 4410 2562 4606
rect 7574 4578 7602 4718
rect 7574 4545 7602 4550
rect 11888 4718 12048 5474
rect 11888 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12048 4718
rect 2534 4377 2562 4382
rect 2218 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2378 4326
rect 2218 3542 2378 4298
rect 2218 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2378 3542
rect 2218 2758 2378 3514
rect 2218 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2378 2758
rect 2218 1974 2378 2730
rect 2218 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2378 1974
rect 2218 1190 2378 1946
rect 2218 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2378 1190
rect 2218 406 2378 1162
rect 11888 3934 12048 4690
rect 11888 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12048 3934
rect 11888 3150 12048 3906
rect 11888 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12048 3150
rect 11888 2366 12048 3122
rect 11888 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12048 2366
rect 11888 1582 12048 2338
rect 11888 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12048 1582
rect 6006 938 6034 943
rect 6006 714 6034 910
rect 6006 681 6034 686
rect 11888 798 12048 1554
rect 11888 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12048 798
rect 2218 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2378 406
rect 2218 0 2378 378
rect 11888 0 12048 770
rect 12218 6678 12378 7112
rect 12218 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12378 6678
rect 12218 5894 12378 6650
rect 12218 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12378 5894
rect 12218 5110 12378 5866
rect 12558 7042 12586 7047
rect 12558 5642 12586 7014
rect 12558 5609 12586 5614
rect 12218 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12378 5110
rect 12218 4326 12378 5082
rect 12218 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12378 4326
rect 12218 3542 12378 4298
rect 12218 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12378 3542
rect 12218 2758 12378 3514
rect 12218 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12378 2758
rect 12218 1974 12378 2730
rect 12218 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12378 1974
rect 12218 1190 12378 1946
rect 12218 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12378 1190
rect 12218 406 12378 1162
rect 12218 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12378 406
rect 12218 0 12378 378
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _00_
timestamp 1486834041
transform 1 0 7056 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _01_
timestamp 1486834041
transform 1 0 7504 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _02_
timestamp 1486834041
transform 1 0 8064 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _03_
timestamp 1486834041
transform 1 0 7728 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _04_
timestamp 1486834041
transform 1 0 6888 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _05_
timestamp 1486834041
transform 1 0 8064 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _06_
timestamp 1486834041
transform 1 0 7616 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _07_
timestamp 1486834041
transform 1 0 6944 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _08_
timestamp 1486834041
transform 1 0 7224 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _09_
timestamp 1486834041
transform 1 0 6720 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _10_
timestamp 1486834041
transform 1 0 7728 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _11_
timestamp 1486834041
transform 1 0 8344 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _12_
timestamp 1486834041
transform 1 0 8288 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _13_
timestamp 1486834041
transform 1 0 7168 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _14_
timestamp 1486834041
transform 1 0 7112 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _15_
timestamp 1486834041
transform 1 0 7280 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _16_
timestamp 1486834041
transform 1 0 7728 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _17_
timestamp 1486834041
transform 1 0 8120 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _18_
timestamp 1486834041
transform 1 0 7560 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _19_
timestamp 1486834041
transform 1 0 8064 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _20_
timestamp 1486834041
transform 1 0 7616 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _21_
timestamp 1486834041
transform 1 0 7504 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _22_
timestamp 1486834041
transform 1 0 7728 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _23_
timestamp 1486834041
transform 1 0 7168 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _24_
timestamp 1486834041
transform 1 0 8792 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _25_
timestamp 1486834041
transform 1 0 7784 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _26_
timestamp 1486834041
transform 1 0 8568 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _27_
timestamp 1486834041
transform 1 0 11424 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _28_
timestamp 1486834041
transform 1 0 9688 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _29_
timestamp 1486834041
transform 1 0 10136 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _30_
timestamp 1486834041
transform 1 0 10640 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _31_
timestamp 1486834041
transform 1 0 14952 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _32_
timestamp 1486834041
transform 1 0 9240 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _33_
timestamp 1486834041
transform 1 0 9744 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _34_
timestamp 1486834041
transform 1 0 10304 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _35_
timestamp 1486834041
transform 1 0 10752 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _36_
timestamp 1486834041
transform 1 0 13384 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _37_
timestamp 1486834041
transform -1 0 1904 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _38_
timestamp 1486834041
transform -1 0 5880 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _39_
timestamp 1486834041
transform 1 0 6216 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _40_
timestamp 1486834041
transform -1 0 7056 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _41_
timestamp 1486834041
transform 1 0 8848 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _42_
timestamp 1486834041
transform 1 0 11256 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _43_
timestamp 1486834041
transform 1 0 11312 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _44_
timestamp 1486834041
transform 1 0 10472 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _45_
timestamp 1486834041
transform 1 0 11704 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _46_
timestamp 1486834041
transform 1 0 12488 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _47_
timestamp 1486834041
transform -1 0 11480 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _48_
timestamp 1486834041
transform 1 0 12656 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _49_
timestamp 1486834041
transform 1 0 13216 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _50_
timestamp 1486834041
transform 1 0 14168 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _51_
timestamp 1486834041
transform -1 0 14616 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _52_
timestamp 1486834041
transform -1 0 4816 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _53_
timestamp 1486834041
transform -1 0 3808 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _54_
timestamp 1486834041
transform -1 0 2688 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _55_
timestamp 1486834041
transform -1 0 2240 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _56_
timestamp 1486834041
transform -1 0 7560 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _57_
timestamp 1486834041
transform -1 0 7280 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _58_
timestamp 1486834041
transform -1 0 4872 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _59_
timestamp 1486834041
transform -1 0 6328 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _60_
timestamp 1486834041
transform -1 0 6104 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _61_
timestamp 1486834041
transform -1 0 5376 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _62_
timestamp 1486834041
transform -1 0 5544 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _63_
timestamp 1486834041
transform -1 0 5880 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _64_
timestamp 1486834041
transform -1 0 9128 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _65_
timestamp 1486834041
transform -1 0 8680 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _66_
timestamp 1486834041
transform -1 0 8232 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _67_
timestamp 1486834041
transform -1 0 7952 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _68_
timestamp 1486834041
transform -1 0 6664 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _69_
timestamp 1486834041
transform -1 0 7784 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _70_
timestamp 1486834041
transform -1 0 3080 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _71_
timestamp 1486834041
transform -1 0 4256 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _72_
timestamp 1486834041
transform 1 0 14168 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _73_
timestamp 1486834041
transform 1 0 11872 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _74_
timestamp 1486834041
transform 1 0 11480 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _75_
timestamp 1486834041
transform 1 0 11032 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _76_
timestamp 1486834041
transform 1 0 10584 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _77_
timestamp 1486834041
transform 1 0 10472 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _78_
timestamp 1486834041
transform -1 0 10136 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _79_
timestamp 1486834041
transform -1 0 9632 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _80_
timestamp 1486834041
transform -1 0 9184 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _81_
timestamp 1486834041
transform -1 0 9576 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _82_
timestamp 1486834041
transform -1 0 4424 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _83_
timestamp 1486834041
transform -1 0 3080 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _84_
timestamp 1486834041
transform 1 0 9688 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _85_
timestamp 1486834041
transform 1 0 9408 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _86_
timestamp 1486834041
transform -1 0 9240 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _87_
timestamp 1486834041
transform -1 0 6832 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _88_
timestamp 1486834041
transform 1 0 9968 0 1 392
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2
timestamp 1486834041
transform 1 0 448 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36
timestamp 1486834041
transform 1 0 2352 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70
timestamp 1486834041
transform 1 0 4256 0 1 392
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86
timestamp 1486834041
transform 1 0 5152 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90
timestamp 1486834041
transform 1 0 5376 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99
timestamp 1486834041
transform 1 0 5880 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101
timestamp 1486834041
transform 1 0 5992 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1486834041
transform 1 0 6160 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_113
timestamp 1486834041
transform 1 0 6664 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_121
timestamp 1486834041
transform 1 0 7112 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_125
timestamp 1486834041
transform 1 0 7336 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_127
timestamp 1486834041
transform 1 0 7448 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_146
timestamp 1486834041
transform 1 0 8512 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_150
timestamp 1486834041
transform 1 0 8736 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_160
timestamp 1486834041
transform 1 0 9296 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_168
timestamp 1486834041
transform 1 0 9744 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_178
timestamp 1486834041
transform 1 0 10304 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_180
timestamp 1486834041
transform 1 0 10416 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189
timestamp 1486834041
transform 1 0 10920 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_193
timestamp 1486834041
transform 1 0 11144 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195
timestamp 1486834041
transform 1 0 11256 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_206
timestamp 1486834041
transform 1 0 11872 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_240
timestamp 1486834041
transform 1 0 13776 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2
timestamp 1486834041
transform 1 0 448 0 -1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1486834041
transform 1 0 4032 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_72
timestamp 1486834041
transform 1 0 4368 0 -1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_104
timestamp 1486834041
transform 1 0 6160 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_128
timestamp 1486834041
transform 1 0 7504 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_142
timestamp 1486834041
transform 1 0 8288 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_158
timestamp 1486834041
transform 1 0 9184 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_167
timestamp 1486834041
transform 1 0 9688 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_176
timestamp 1486834041
transform 1 0 10192 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_194
timestamp 1486834041
transform 1 0 11200 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_203
timestamp 1486834041
transform 1 0 11704 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_207
timestamp 1486834041
transform 1 0 11928 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_209
timestamp 1486834041
transform 1 0 12040 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_212
timestamp 1486834041
transform 1 0 12208 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_216
timestamp 1486834041
transform 1 0 12432 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_225
timestamp 1486834041
transform 1 0 12936 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1486834041
transform 1 0 448 0 1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1486834041
transform 1 0 2240 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1486834041
transform 1 0 2408 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1486834041
transform 1 0 5992 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_107
timestamp 1486834041
transform 1 0 6328 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_115
timestamp 1486834041
transform 1 0 6776 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_117
timestamp 1486834041
transform 1 0 6888 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_126
timestamp 1486834041
transform 1 0 7392 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_146
timestamp 1486834041
transform 1 0 8512 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_155
timestamp 1486834041
transform 1 0 9016 0 1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 9912 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_177
timestamp 1486834041
transform 1 0 10248 0 1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_193
timestamp 1486834041
transform 1 0 11144 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_201
timestamp 1486834041
transform 1 0 11592 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_211
timestamp 1486834041
transform 1 0 12152 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_219
timestamp 1486834041
transform 1 0 12600 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_228
timestamp 1486834041
transform 1 0 13104 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_230
timestamp 1486834041
transform 1 0 13216 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1486834041
transform 1 0 448 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1486834041
transform 1 0 4032 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_72
timestamp 1486834041
transform 1 0 4368 0 -1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_104
timestamp 1486834041
transform 1 0 6160 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_112
timestamp 1486834041
transform 1 0 6608 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_116
timestamp 1486834041
transform 1 0 6832 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_125
timestamp 1486834041
transform 1 0 7336 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_133
timestamp 1486834041
transform 1 0 7784 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_137
timestamp 1486834041
transform 1 0 8008 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_139
timestamp 1486834041
transform 1 0 8120 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_142
timestamp 1486834041
transform 1 0 8288 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_206
timestamp 1486834041
transform 1 0 11872 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_212
timestamp 1486834041
transform 1 0 12208 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_228
timestamp 1486834041
transform 1 0 13104 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_238
timestamp 1486834041
transform 1 0 13664 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_240
timestamp 1486834041
transform 1 0 13776 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1486834041
transform 1 0 448 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 2240 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1486834041
transform 1 0 2408 0 1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1486834041
transform 1 0 5992 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_107
timestamp 1486834041
transform 1 0 6328 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_131
timestamp 1486834041
transform 1 0 7672 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_141
timestamp 1486834041
transform 1 0 8232 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_173
timestamp 1486834041
transform 1 0 10024 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_177
timestamp 1486834041
transform 1 0 10248 0 1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_241
timestamp 1486834041
transform 1 0 13832 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_247
timestamp 1486834041
transform 1 0 14168 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1486834041
transform 1 0 448 0 -1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1486834041
transform 1 0 4032 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_72
timestamp 1486834041
transform 1 0 4368 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_104
timestamp 1486834041
transform 1 0 6160 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_112
timestamp 1486834041
transform 1 0 6608 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_130
timestamp 1486834041
transform 1 0 7616 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_142
timestamp 1486834041
transform 1 0 8288 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_159
timestamp 1486834041
transform 1 0 9240 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_191
timestamp 1486834041
transform 1 0 11032 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_207
timestamp 1486834041
transform 1 0 11928 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_209
timestamp 1486834041
transform 1 0 12040 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_212
timestamp 1486834041
transform 1 0 12208 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_228
timestamp 1486834041
transform 1 0 13104 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_236
timestamp 1486834041
transform 1 0 13552 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_240
timestamp 1486834041
transform 1 0 13776 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1486834041
transform 1 0 448 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 2240 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1486834041
transform 1 0 2408 0 1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1486834041
transform 1 0 5992 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_107
timestamp 1486834041
transform 1 0 6328 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_115
timestamp 1486834041
transform 1 0 6776 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_119
timestamp 1486834041
transform 1 0 7000 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_121
timestamp 1486834041
transform 1 0 7112 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_130
timestamp 1486834041
transform 1 0 7616 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_162
timestamp 1486834041
transform 1 0 9408 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_170
timestamp 1486834041
transform 1 0 9856 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_174
timestamp 1486834041
transform 1 0 10080 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_177
timestamp 1486834041
transform 1 0 10248 0 1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_241
timestamp 1486834041
transform 1 0 13832 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_247
timestamp 1486834041
transform 1 0 14168 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_2
timestamp 1486834041
transform 1 0 448 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_34
timestamp 1486834041
transform 1 0 2240 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_50
timestamp 1486834041
transform 1 0 3136 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_58
timestamp 1486834041
transform 1 0 3584 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_72
timestamp 1486834041
transform 1 0 4368 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_104
timestamp 1486834041
transform 1 0 6160 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_120
timestamp 1486834041
transform 1 0 7056 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_129
timestamp 1486834041
transform 1 0 7560 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_137
timestamp 1486834041
transform 1 0 8008 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_139
timestamp 1486834041
transform 1 0 8120 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_150
timestamp 1486834041
transform 1 0 8736 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_182
timestamp 1486834041
transform 1 0 10528 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_198
timestamp 1486834041
transform 1 0 11424 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_206
timestamp 1486834041
transform 1 0 11872 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_212
timestamp 1486834041
transform 1 0 12208 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_220
timestamp 1486834041
transform 1 0 12656 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_224
timestamp 1486834041
transform 1 0 12880 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_226
timestamp 1486834041
transform 1 0 12992 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1486834041
transform 1 0 448 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 2240 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_37
timestamp 1486834041
transform 1 0 2408 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_53
timestamp 1486834041
transform 1 0 3304 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_62
timestamp 1486834041
transform 1 0 3808 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_64
timestamp 1486834041
transform 1 0 3920 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_73
timestamp 1486834041
transform 1 0 4424 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_81
timestamp 1486834041
transform 1 0 4872 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_93
timestamp 1486834041
transform 1 0 5544 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1486834041
transform 1 0 5992 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_107
timestamp 1486834041
transform 1 0 6328 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_123
timestamp 1486834041
transform 1 0 7224 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_140
timestamp 1486834041
transform 1 0 8176 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_172
timestamp 1486834041
transform 1 0 9968 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_174
timestamp 1486834041
transform 1 0 10080 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_177
timestamp 1486834041
transform 1 0 10248 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_209
timestamp 1486834041
transform 1 0 12040 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_247
timestamp 1486834041
transform 1 0 14168 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_2
timestamp 1486834041
transform 1 0 448 0 -1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_80
timestamp 1486834041
transform 1 0 4816 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_90
timestamp 1486834041
transform 1 0 5376 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_107
timestamp 1486834041
transform 1 0 6328 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_123
timestamp 1486834041
transform 1 0 7224 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_131
timestamp 1486834041
transform 1 0 7672 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_142
timestamp 1486834041
transform 1 0 8288 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_206
timestamp 1486834041
transform 1 0 11872 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1486834041
transform 1 0 12208 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_2
timestamp 1486834041
transform 1 0 448 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_18
timestamp 1486834041
transform 1 0 1344 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1486834041
transform 1 0 2240 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_37
timestamp 1486834041
transform 1 0 2408 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_103
timestamp 1486834041
transform 1 0 6104 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_107
timestamp 1486834041
transform 1 0 6328 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_123
timestamp 1486834041
transform 1 0 7224 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_127
timestamp 1486834041
transform 1 0 7448 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_136
timestamp 1486834041
transform 1 0 7952 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_138
timestamp 1486834041
transform 1 0 8064 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_147
timestamp 1486834041
transform 1 0 8568 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_163
timestamp 1486834041
transform 1 0 9464 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_171
timestamp 1486834041
transform 1 0 9912 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_177
timestamp 1486834041
transform 1 0 10248 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_193
timestamp 1486834041
transform 1 0 11144 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_197
timestamp 1486834041
transform 1 0 11368 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_214
timestamp 1486834041
transform 1 0 12320 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_216
timestamp 1486834041
transform 1 0 12432 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_2
timestamp 1486834041
transform 1 0 448 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_18
timestamp 1486834041
transform 1 0 1344 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_26
timestamp 1486834041
transform 1 0 1792 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_72
timestamp 1486834041
transform 1 0 4368 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_76
timestamp 1486834041
transform 1 0 4592 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_105
timestamp 1486834041
transform 1 0 6216 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_107
timestamp 1486834041
transform 1 0 6328 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_124
timestamp 1486834041
transform 1 0 7280 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_142
timestamp 1486834041
transform 1 0 8288 0 -1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_174
timestamp 1486834041
transform 1 0 10080 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_178
timestamp 1486834041
transform 1 0 10304 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_180
timestamp 1486834041
transform 1 0 10416 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_189
timestamp 1486834041
transform 1 0 10920 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_207
timestamp 1486834041
transform 1 0 11928 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_209
timestamp 1486834041
transform 1 0 12040 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_240
timestamp 1486834041
transform 1 0 13776 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_2
timestamp 1486834041
transform 1 0 448 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_18
timestamp 1486834041
transform 1 0 1344 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_20
timestamp 1486834041
transform 1 0 1456 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_37
timestamp 1486834041
transform 1 0 2408 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_129
timestamp 1486834041
transform 1 0 7560 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_146
timestamp 1486834041
transform 1 0 8512 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_166
timestamp 1486834041
transform 1 0 9632 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_241
timestamp 1486834041
transform 1 0 13832 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_2
timestamp 1486834041
transform 1 0 448 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_18
timestamp 1486834041
transform 1 0 1344 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_72
timestamp 1486834041
transform 1 0 4368 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_123
timestamp 1486834041
transform 1 0 7224 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_127
timestamp 1486834041
transform 1 0 7448 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_137
timestamp 1486834041
transform 1 0 8008 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_139
timestamp 1486834041
transform 1 0 8120 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_142
timestamp 1486834041
transform 1 0 8288 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_158
timestamp 1486834041
transform 1 0 9184 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_166
timestamp 1486834041
transform 1 0 9632 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_183
timestamp 1486834041
transform 1 0 10584 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_192
timestamp 1486834041
transform 1 0 11088 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_194
timestamp 1486834041
transform 1 0 11200 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_209
timestamp 1486834041
transform 1 0 12040 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_254
timestamp 1486834041
transform 1 0 14560 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_2
timestamp 1486834041
transform 1 0 448 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_18
timestamp 1486834041
transform 1 0 1344 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_20
timestamp 1486834041
transform 1 0 1456 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_37
timestamp 1486834041
transform 1 0 2408 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_107
timestamp 1486834041
transform 1 0 6328 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_165
timestamp 1486834041
transform 1 0 9576 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_241
timestamp 1486834041
transform 1 0 13832 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_2
timestamp 1486834041
transform 1 0 448 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_36
timestamp 1486834041
transform 1 0 2352 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_70
timestamp 1486834041
transform 1 0 4256 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_104
timestamp 1486834041
transform 1 0 6160 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_127
timestamp 1486834041
transform 1 0 7448 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_138
timestamp 1486834041
transform 1 0 8064 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_146
timestamp 1486834041
transform 1 0 8512 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_150
timestamp 1486834041
transform 1 0 8736 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_159
timestamp 1486834041
transform 1 0 9240 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_161
timestamp 1486834041
transform 1 0 9352 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_172
timestamp 1486834041
transform 1 0 9968 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_174
timestamp 1486834041
transform 1 0 10080 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_203
timestamp 1486834041
transform 1 0 11704 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_234
timestamp 1486834041
transform 1 0 13440 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_268
timestamp 1486834041
transform 1 0 15344 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform 1 0 13272 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform 1 0 14616 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform 1 0 13832 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform 1 0 14616 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform 1 0 14616 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform 1 0 13832 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform 1 0 14616 0 1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform 1 0 14616 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform 1 0 14616 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform 1 0 14616 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform 1 0 14616 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform 1 0 12096 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform 1 0 14616 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform 1 0 14616 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 14616 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 13832 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform 1 0 13832 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 13048 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform 1 0 13272 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform -1 0 10920 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform 1 0 12264 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform 1 0 13048 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 12880 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform -1 0 11032 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform -1 0 13272 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 13048 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 13832 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 13832 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 14616 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 14616 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform 1 0 13832 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 14616 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform 1 0 10920 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform 1 0 12992 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform 1 0 12208 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform 1 0 13776 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform 1 0 13048 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform -1 0 13272 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform 1 0 13776 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform 1 0 14168 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform -1 0 13776 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform 1 0 14560 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform -1 0 14056 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform 1 0 11032 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform 1 0 11872 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform 1 0 11256 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform -1 0 12600 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform 1 0 11480 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform 1 0 12656 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform 1 0 12600 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform 1 0 12208 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform 1 0 12264 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform -1 0 2296 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform -1 0 3472 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform 1 0 1904 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform 1 0 2520 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform -1 0 1456 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform -1 0 2688 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform -1 0 2296 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform -1 0 3472 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform -1 0 4256 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform -1 0 4088 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform -1 0 2240 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform -1 0 3472 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform -1 0 3864 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform -1 0 4256 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform -1 0 4872 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform -1 0 3360 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform -1 0 4256 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform -1 0 4648 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform 1 0 3080 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform 1 0 4872 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform -1 0 5432 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform 1 0 5656 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform 1 0 5432 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform -1 0 6048 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform -1 0 7224 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform -1 0 7336 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform 1 0 6664 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform -1 0 4144 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform -1 0 4648 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform -1 0 5432 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform -1 0 6216 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform -1 0 5656 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform -1 0 5432 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform -1 0 6216 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform -1 0 5264 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform -1 0 7112 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output89
timestamp 1486834041
transform 1 0 10248 0 1 5096
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_16
timestamp 1486834041
transform 1 0 336 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 15512 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_17
timestamp 1486834041
transform 1 0 336 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 15512 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_18
timestamp 1486834041
transform 1 0 336 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 15512 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_19
timestamp 1486834041
transform 1 0 336 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 15512 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_20
timestamp 1486834041
transform 1 0 336 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 15512 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_21
timestamp 1486834041
transform 1 0 336 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 15512 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_22
timestamp 1486834041
transform 1 0 336 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 15512 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_23
timestamp 1486834041
transform 1 0 336 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 15512 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_24
timestamp 1486834041
transform 1 0 336 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 15512 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_25
timestamp 1486834041
transform 1 0 336 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 15512 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_26
timestamp 1486834041
transform 1 0 336 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 15512 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_27
timestamp 1486834041
transform 1 0 336 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 15512 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_28
timestamp 1486834041
transform 1 0 336 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 15512 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_29
timestamp 1486834041
transform 1 0 336 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 15512 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_30
timestamp 1486834041
transform 1 0 336 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 15512 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_31
timestamp 1486834041
transform 1 0 336 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 15512 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_32
timestamp 1486834041
transform 1 0 2240 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_33
timestamp 1486834041
transform 1 0 4144 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34
timestamp 1486834041
transform 1 0 6048 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1486834041
transform 1 0 7952 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1486834041
transform 1 0 9856 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1486834041
transform 1 0 11760 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1486834041
transform 1 0 13664 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_39
timestamp 1486834041
transform 1 0 4256 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_40
timestamp 1486834041
transform 1 0 8176 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_41
timestamp 1486834041
transform 1 0 12096 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_42
timestamp 1486834041
transform 1 0 2296 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_43
timestamp 1486834041
transform 1 0 6216 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_44
timestamp 1486834041
transform 1 0 10136 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_45
timestamp 1486834041
transform 1 0 14056 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_46
timestamp 1486834041
transform 1 0 4256 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_47
timestamp 1486834041
transform 1 0 8176 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_48
timestamp 1486834041
transform 1 0 12096 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_49
timestamp 1486834041
transform 1 0 2296 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_50
timestamp 1486834041
transform 1 0 6216 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_51
timestamp 1486834041
transform 1 0 10136 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_52
timestamp 1486834041
transform 1 0 14056 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_53
timestamp 1486834041
transform 1 0 4256 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_54
timestamp 1486834041
transform 1 0 8176 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_55
timestamp 1486834041
transform 1 0 12096 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_56
timestamp 1486834041
transform 1 0 2296 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_57
timestamp 1486834041
transform 1 0 6216 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_58
timestamp 1486834041
transform 1 0 10136 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_59
timestamp 1486834041
transform 1 0 14056 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_60
timestamp 1486834041
transform 1 0 4256 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_61
timestamp 1486834041
transform 1 0 8176 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_62
timestamp 1486834041
transform 1 0 12096 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_63
timestamp 1486834041
transform 1 0 2296 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_64
timestamp 1486834041
transform 1 0 6216 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_65
timestamp 1486834041
transform 1 0 10136 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_66
timestamp 1486834041
transform 1 0 14056 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_67
timestamp 1486834041
transform 1 0 4256 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_68
timestamp 1486834041
transform 1 0 8176 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_69
timestamp 1486834041
transform 1 0 12096 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_70
timestamp 1486834041
transform 1 0 2296 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_71
timestamp 1486834041
transform 1 0 6216 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_72
timestamp 1486834041
transform 1 0 10136 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_73
timestamp 1486834041
transform 1 0 14056 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_74
timestamp 1486834041
transform 1 0 4256 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_75
timestamp 1486834041
transform 1 0 8176 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_76
timestamp 1486834041
transform 1 0 12096 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_77
timestamp 1486834041
transform 1 0 2296 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_78
timestamp 1486834041
transform 1 0 6216 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_79
timestamp 1486834041
transform 1 0 10136 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_80
timestamp 1486834041
transform 1 0 14056 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_81
timestamp 1486834041
transform 1 0 4256 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_82
timestamp 1486834041
transform 1 0 8176 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_83
timestamp 1486834041
transform 1 0 12096 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_84
timestamp 1486834041
transform 1 0 2296 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_85
timestamp 1486834041
transform 1 0 6216 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_86
timestamp 1486834041
transform 1 0 10136 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_87
timestamp 1486834041
transform 1 0 14056 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_88
timestamp 1486834041
transform 1 0 2240 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_89
timestamp 1486834041
transform 1 0 4144 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_90
timestamp 1486834041
transform 1 0 6048 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_91
timestamp 1486834041
transform 1 0 7952 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_92
timestamp 1486834041
transform 1 0 9856 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_93
timestamp 1486834041
transform 1 0 11760 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_94
timestamp 1486834041
transform 1 0 13664 0 -1 6664
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 0 56 56 0 FreeSans 224 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 2240 56 2296 0 FreeSans 224 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 2464 56 2520 0 FreeSans 224 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 2688 56 2744 0 FreeSans 224 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 2912 56 2968 0 FreeSans 224 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 3136 56 3192 0 FreeSans 224 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 3360 56 3416 0 FreeSans 224 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 3584 56 3640 0 FreeSans 224 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 3808 56 3864 0 FreeSans 224 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 4032 56 4088 0 FreeSans 224 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 4256 56 4312 0 FreeSans 224 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 224 56 280 0 FreeSans 224 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 4480 56 4536 0 FreeSans 224 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 4704 56 4760 0 FreeSans 224 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 4928 56 4984 0 FreeSans 224 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 5152 56 5208 0 FreeSans 224 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 5376 56 5432 0 FreeSans 224 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 5600 56 5656 0 FreeSans 224 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 5824 56 5880 0 FreeSans 224 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 6048 56 6104 0 FreeSans 224 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 6272 56 6328 0 FreeSans 224 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 6496 56 6552 0 FreeSans 224 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 448 56 504 0 FreeSans 224 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 6720 56 6776 0 FreeSans 224 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 6944 56 7000 0 FreeSans 224 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 672 56 728 0 FreeSans 224 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 896 56 952 0 FreeSans 224 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 1120 56 1176 0 FreeSans 224 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 1344 56 1400 0 FreeSans 224 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 1568 56 1624 0 FreeSans 224 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 1792 56 1848 0 FreeSans 224 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 2016 56 2072 0 FreeSans 224 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 15792 0 15848 56 0 FreeSans 224 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 15792 2240 15848 2296 0 FreeSans 224 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 15792 2464 15848 2520 0 FreeSans 224 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 15792 2688 15848 2744 0 FreeSans 224 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 15792 2912 15848 2968 0 FreeSans 224 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 15792 3136 15848 3192 0 FreeSans 224 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 15792 3360 15848 3416 0 FreeSans 224 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 15792 3584 15848 3640 0 FreeSans 224 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 15792 3808 15848 3864 0 FreeSans 224 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 15792 4032 15848 4088 0 FreeSans 224 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 15792 4256 15848 4312 0 FreeSans 224 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 15792 224 15848 280 0 FreeSans 224 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 15792 4480 15848 4536 0 FreeSans 224 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 15792 4704 15848 4760 0 FreeSans 224 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 15792 4928 15848 4984 0 FreeSans 224 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 15792 5152 15848 5208 0 FreeSans 224 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 15792 5376 15848 5432 0 FreeSans 224 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 15792 5600 15848 5656 0 FreeSans 224 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 15792 5824 15848 5880 0 FreeSans 224 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 15792 6048 15848 6104 0 FreeSans 224 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 15792 6272 15848 6328 0 FreeSans 224 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 15792 6496 15848 6552 0 FreeSans 224 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 15792 448 15848 504 0 FreeSans 224 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 15792 6720 15848 6776 0 FreeSans 224 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 15792 6944 15848 7000 0 FreeSans 224 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 15792 672 15848 728 0 FreeSans 224 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 15792 896 15848 952 0 FreeSans 224 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 15792 1120 15848 1176 0 FreeSans 224 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 15792 1344 15848 1400 0 FreeSans 224 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 15792 1568 15848 1624 0 FreeSans 224 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 15792 1792 15848 1848 0 FreeSans 224 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 15792 2016 15848 2072 0 FreeSans 224 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 1792 0 1848 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 8512 0 8568 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 9184 0 9240 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 9856 0 9912 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 10528 0 10584 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 11200 0 11256 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 11872 0 11928 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 12544 0 12600 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 13216 0 13272 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 13888 0 13944 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 14560 0 14616 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 2464 0 2520 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 3136 0 3192 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 3808 0 3864 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 4480 0 4536 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 5152 0 5208 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 5824 0 5880 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 6496 0 6552 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 7168 0 7224 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 7840 0 7896 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 10864 7056 10920 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 11984 7056 12040 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 12096 7056 12152 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 12208 7056 12264 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 12320 7056 12376 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 12432 7056 12488 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 12544 7056 12600 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 12656 7056 12712 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 12768 7056 12824 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 12880 7056 12936 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 12992 7056 13048 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 10976 7056 11032 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 11088 7056 11144 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 11200 7056 11256 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 11312 7056 11368 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 11424 7056 11480 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 11536 7056 11592 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 11648 7056 11704 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 11760 7056 11816 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 11872 7056 11928 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 2688 7056 2744 7112 0 FreeSans 224 0 0 0 N1BEG[0]
port 104 nsew signal output
flabel metal2 s 2800 7056 2856 7112 0 FreeSans 224 0 0 0 N1BEG[1]
port 105 nsew signal output
flabel metal2 s 2912 7056 2968 7112 0 FreeSans 224 0 0 0 N1BEG[2]
port 106 nsew signal output
flabel metal2 s 3024 7056 3080 7112 0 FreeSans 224 0 0 0 N1BEG[3]
port 107 nsew signal output
flabel metal2 s 3136 7056 3192 7112 0 FreeSans 224 0 0 0 N2BEG[0]
port 108 nsew signal output
flabel metal2 s 3248 7056 3304 7112 0 FreeSans 224 0 0 0 N2BEG[1]
port 109 nsew signal output
flabel metal2 s 3360 7056 3416 7112 0 FreeSans 224 0 0 0 N2BEG[2]
port 110 nsew signal output
flabel metal2 s 3472 7056 3528 7112 0 FreeSans 224 0 0 0 N2BEG[3]
port 111 nsew signal output
flabel metal2 s 3584 7056 3640 7112 0 FreeSans 224 0 0 0 N2BEG[4]
port 112 nsew signal output
flabel metal2 s 3696 7056 3752 7112 0 FreeSans 224 0 0 0 N2BEG[5]
port 113 nsew signal output
flabel metal2 s 3808 7056 3864 7112 0 FreeSans 224 0 0 0 N2BEG[6]
port 114 nsew signal output
flabel metal2 s 3920 7056 3976 7112 0 FreeSans 224 0 0 0 N2BEG[7]
port 115 nsew signal output
flabel metal2 s 4032 7056 4088 7112 0 FreeSans 224 0 0 0 N2BEGb[0]
port 116 nsew signal output
flabel metal2 s 4144 7056 4200 7112 0 FreeSans 224 0 0 0 N2BEGb[1]
port 117 nsew signal output
flabel metal2 s 4256 7056 4312 7112 0 FreeSans 224 0 0 0 N2BEGb[2]
port 118 nsew signal output
flabel metal2 s 4368 7056 4424 7112 0 FreeSans 224 0 0 0 N2BEGb[3]
port 119 nsew signal output
flabel metal2 s 4480 7056 4536 7112 0 FreeSans 224 0 0 0 N2BEGb[4]
port 120 nsew signal output
flabel metal2 s 4592 7056 4648 7112 0 FreeSans 224 0 0 0 N2BEGb[5]
port 121 nsew signal output
flabel metal2 s 4704 7056 4760 7112 0 FreeSans 224 0 0 0 N2BEGb[6]
port 122 nsew signal output
flabel metal2 s 4816 7056 4872 7112 0 FreeSans 224 0 0 0 N2BEGb[7]
port 123 nsew signal output
flabel metal2 s 4928 7056 4984 7112 0 FreeSans 224 0 0 0 N4BEG[0]
port 124 nsew signal output
flabel metal2 s 6048 7056 6104 7112 0 FreeSans 224 0 0 0 N4BEG[10]
port 125 nsew signal output
flabel metal2 s 6160 7056 6216 7112 0 FreeSans 224 0 0 0 N4BEG[11]
port 126 nsew signal output
flabel metal2 s 6272 7056 6328 7112 0 FreeSans 224 0 0 0 N4BEG[12]
port 127 nsew signal output
flabel metal2 s 6384 7056 6440 7112 0 FreeSans 224 0 0 0 N4BEG[13]
port 128 nsew signal output
flabel metal2 s 6496 7056 6552 7112 0 FreeSans 224 0 0 0 N4BEG[14]
port 129 nsew signal output
flabel metal2 s 6608 7056 6664 7112 0 FreeSans 224 0 0 0 N4BEG[15]
port 130 nsew signal output
flabel metal2 s 5040 7056 5096 7112 0 FreeSans 224 0 0 0 N4BEG[1]
port 131 nsew signal output
flabel metal2 s 5152 7056 5208 7112 0 FreeSans 224 0 0 0 N4BEG[2]
port 132 nsew signal output
flabel metal2 s 5264 7056 5320 7112 0 FreeSans 224 0 0 0 N4BEG[3]
port 133 nsew signal output
flabel metal2 s 5376 7056 5432 7112 0 FreeSans 224 0 0 0 N4BEG[4]
port 134 nsew signal output
flabel metal2 s 5488 7056 5544 7112 0 FreeSans 224 0 0 0 N4BEG[5]
port 135 nsew signal output
flabel metal2 s 5600 7056 5656 7112 0 FreeSans 224 0 0 0 N4BEG[6]
port 136 nsew signal output
flabel metal2 s 5712 7056 5768 7112 0 FreeSans 224 0 0 0 N4BEG[7]
port 137 nsew signal output
flabel metal2 s 5824 7056 5880 7112 0 FreeSans 224 0 0 0 N4BEG[8]
port 138 nsew signal output
flabel metal2 s 5936 7056 5992 7112 0 FreeSans 224 0 0 0 N4BEG[9]
port 139 nsew signal output
flabel metal2 s 6720 7056 6776 7112 0 FreeSans 224 0 0 0 S1END[0]
port 140 nsew signal input
flabel metal2 s 6832 7056 6888 7112 0 FreeSans 224 0 0 0 S1END[1]
port 141 nsew signal input
flabel metal2 s 6944 7056 7000 7112 0 FreeSans 224 0 0 0 S1END[2]
port 142 nsew signal input
flabel metal2 s 7056 7056 7112 7112 0 FreeSans 224 0 0 0 S1END[3]
port 143 nsew signal input
flabel metal2 s 8064 7056 8120 7112 0 FreeSans 224 0 0 0 S2END[0]
port 144 nsew signal input
flabel metal2 s 8176 7056 8232 7112 0 FreeSans 224 0 0 0 S2END[1]
port 145 nsew signal input
flabel metal2 s 8288 7056 8344 7112 0 FreeSans 224 0 0 0 S2END[2]
port 146 nsew signal input
flabel metal2 s 8400 7056 8456 7112 0 FreeSans 224 0 0 0 S2END[3]
port 147 nsew signal input
flabel metal2 s 8512 7056 8568 7112 0 FreeSans 224 0 0 0 S2END[4]
port 148 nsew signal input
flabel metal2 s 8624 7056 8680 7112 0 FreeSans 224 0 0 0 S2END[5]
port 149 nsew signal input
flabel metal2 s 8736 7056 8792 7112 0 FreeSans 224 0 0 0 S2END[6]
port 150 nsew signal input
flabel metal2 s 8848 7056 8904 7112 0 FreeSans 224 0 0 0 S2END[7]
port 151 nsew signal input
flabel metal2 s 7168 7056 7224 7112 0 FreeSans 224 0 0 0 S2MID[0]
port 152 nsew signal input
flabel metal2 s 7280 7056 7336 7112 0 FreeSans 224 0 0 0 S2MID[1]
port 153 nsew signal input
flabel metal2 s 7392 7056 7448 7112 0 FreeSans 224 0 0 0 S2MID[2]
port 154 nsew signal input
flabel metal2 s 7504 7056 7560 7112 0 FreeSans 224 0 0 0 S2MID[3]
port 155 nsew signal input
flabel metal2 s 7616 7056 7672 7112 0 FreeSans 224 0 0 0 S2MID[4]
port 156 nsew signal input
flabel metal2 s 7728 7056 7784 7112 0 FreeSans 224 0 0 0 S2MID[5]
port 157 nsew signal input
flabel metal2 s 7840 7056 7896 7112 0 FreeSans 224 0 0 0 S2MID[6]
port 158 nsew signal input
flabel metal2 s 7952 7056 8008 7112 0 FreeSans 224 0 0 0 S2MID[7]
port 159 nsew signal input
flabel metal2 s 8960 7056 9016 7112 0 FreeSans 224 0 0 0 S4END[0]
port 160 nsew signal input
flabel metal2 s 10080 7056 10136 7112 0 FreeSans 224 0 0 0 S4END[10]
port 161 nsew signal input
flabel metal2 s 10192 7056 10248 7112 0 FreeSans 224 0 0 0 S4END[11]
port 162 nsew signal input
flabel metal2 s 10304 7056 10360 7112 0 FreeSans 224 0 0 0 S4END[12]
port 163 nsew signal input
flabel metal2 s 10416 7056 10472 7112 0 FreeSans 224 0 0 0 S4END[13]
port 164 nsew signal input
flabel metal2 s 10528 7056 10584 7112 0 FreeSans 224 0 0 0 S4END[14]
port 165 nsew signal input
flabel metal2 s 10640 7056 10696 7112 0 FreeSans 224 0 0 0 S4END[15]
port 166 nsew signal input
flabel metal2 s 9072 7056 9128 7112 0 FreeSans 224 0 0 0 S4END[1]
port 167 nsew signal input
flabel metal2 s 9184 7056 9240 7112 0 FreeSans 224 0 0 0 S4END[2]
port 168 nsew signal input
flabel metal2 s 9296 7056 9352 7112 0 FreeSans 224 0 0 0 S4END[3]
port 169 nsew signal input
flabel metal2 s 9408 7056 9464 7112 0 FreeSans 224 0 0 0 S4END[4]
port 170 nsew signal input
flabel metal2 s 9520 7056 9576 7112 0 FreeSans 224 0 0 0 S4END[5]
port 171 nsew signal input
flabel metal2 s 9632 7056 9688 7112 0 FreeSans 224 0 0 0 S4END[6]
port 172 nsew signal input
flabel metal2 s 9744 7056 9800 7112 0 FreeSans 224 0 0 0 S4END[7]
port 173 nsew signal input
flabel metal2 s 9856 7056 9912 7112 0 FreeSans 224 0 0 0 S4END[8]
port 174 nsew signal input
flabel metal2 s 9968 7056 10024 7112 0 FreeSans 224 0 0 0 S4END[9]
port 175 nsew signal input
flabel metal2 s 1120 0 1176 56 0 FreeSans 224 0 0 0 UserCLK
port 176 nsew signal input
flabel metal2 s 10752 7056 10808 7112 0 FreeSans 224 0 0 0 UserCLKo
port 177 nsew signal output
flabel metal4 s 1888 0 2048 7112 0 FreeSans 736 90 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 1888 0 2048 28 0 FreeSans 184 0 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 1888 7084 2048 7112 0 FreeSans 184 0 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 11888 0 12048 7112 0 FreeSans 736 90 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 11888 0 12048 28 0 FreeSans 184 0 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 11888 7084 12048 7112 0 FreeSans 184 0 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 2218 0 2378 7112 0 FreeSans 736 90 0 0 VSS
port 179 nsew ground bidirectional
flabel metal4 s 2218 0 2378 28 0 FreeSans 184 0 0 0 VSS
port 179 nsew ground bidirectional
flabel metal4 s 2218 7084 2378 7112 0 FreeSans 184 0 0 0 VSS
port 179 nsew ground bidirectional
flabel metal4 s 12218 0 12378 7112 0 FreeSans 736 90 0 0 VSS
port 179 nsew ground bidirectional
flabel metal4 s 12218 0 12378 28 0 FreeSans 184 0 0 0 VSS
port 179 nsew ground bidirectional
flabel metal4 s 12218 7084 12378 7112 0 FreeSans 184 0 0 0 VSS
port 179 nsew ground bidirectional
rlabel metal1 7924 6272 7924 6272 0 VDD
rlabel metal1 7924 6664 7924 6664 0 VSS
rlabel metal3 539 28 539 28 0 FrameData[0]
rlabel metal2 7812 2408 7812 2408 0 FrameData[10]
rlabel metal2 8428 2520 8428 2520 0 FrameData[11]
rlabel metal3 1071 2716 1071 2716 0 FrameData[12]
rlabel metal2 7196 2800 7196 2800 0 FrameData[13]
rlabel metal3 91 3164 91 3164 0 FrameData[14]
rlabel metal2 7364 3500 7364 3500 0 FrameData[15]
rlabel metal3 1099 3612 1099 3612 0 FrameData[16]
rlabel metal2 8204 4116 8204 4116 0 FrameData[17]
rlabel metal3 371 4060 371 4060 0 FrameData[18]
rlabel metal3 1071 4284 1071 4284 0 FrameData[19]
rlabel metal2 7588 364 7588 364 0 FrameData[1]
rlabel metal2 5852 4788 5852 4788 0 FrameData[20]
rlabel metal3 931 4732 931 4732 0 FrameData[21]
rlabel metal3 2135 4956 2135 4956 0 FrameData[22]
rlabel metal3 427 5180 427 5180 0 FrameData[23]
rlabel metal3 567 5404 567 5404 0 FrameData[24]
rlabel metal3 1904 3668 1904 3668 0 FrameData[25]
rlabel metal3 483 5852 483 5852 0 FrameData[26]
rlabel metal2 224 4116 224 4116 0 FrameData[27]
rlabel metal3 651 6300 651 6300 0 FrameData[28]
rlabel metal3 91 6524 91 6524 0 FrameData[29]
rlabel metal3 4095 476 4095 476 0 FrameData[2]
rlabel metal3 175 6748 175 6748 0 FrameData[30]
rlabel metal3 952 812 952 812 0 FrameData[31]
rlabel metal4 6020 812 6020 812 0 FrameData[3]
rlabel metal3 1071 924 1071 924 0 FrameData[4]
rlabel metal3 1071 1148 1071 1148 0 FrameData[5]
rlabel metal3 3871 1372 3871 1372 0 FrameData[6]
rlabel metal3 931 1596 931 1596 0 FrameData[7]
rlabel metal2 7308 1932 7308 1932 0 FrameData[8]
rlabel metal2 6804 2296 6804 2296 0 FrameData[9]
rlabel metal3 14777 28 14777 28 0 FrameData_O[0]
rlabel metal2 15204 1988 15204 1988 0 FrameData_O[10]
rlabel metal3 15113 2492 15113 2492 0 FrameData_O[11]
rlabel metal2 15148 2464 15148 2464 0 FrameData_O[12]
rlabel metal2 15092 2772 15092 2772 0 FrameData_O[13]
rlabel metal3 15113 3164 15113 3164 0 FrameData_O[14]
rlabel metal2 15148 3192 15148 3192 0 FrameData_O[15]
rlabel metal2 15204 3444 15204 3444 0 FrameData_O[16]
rlabel metal3 15505 3836 15505 3836 0 FrameData_O[17]
rlabel metal2 15148 3920 15148 3920 0 FrameData_O[18]
rlabel metal3 15449 4284 15449 4284 0 FrameData_O[19]
rlabel metal3 14133 252 14133 252 0 FrameData_O[1]
rlabel metal3 15505 4508 15505 4508 0 FrameData_O[20]
rlabel metal3 15449 4732 15449 4732 0 FrameData_O[21]
rlabel metal3 15505 4956 15505 4956 0 FrameData_O[22]
rlabel metal2 14308 5068 14308 5068 0 FrameData_O[23]
rlabel metal3 15113 5404 15113 5404 0 FrameData_O[24]
rlabel metal3 14721 5628 14721 5628 0 FrameData_O[25]
rlabel metal2 13860 4018 13860 4018 0 FrameData_O[26]
rlabel metal2 10500 6244 10500 6244 0 FrameData_O[27]
rlabel metal2 12740 5236 12740 5236 0 FrameData_O[28]
rlabel metal2 13664 3276 13664 3276 0 FrameData_O[29]
rlabel metal3 14581 476 14581 476 0 FrameData_O[2]
rlabel metal3 15057 6748 15057 6748 0 FrameData_O[30]
rlabel metal3 15141 6972 15141 6972 0 FrameData_O[31]
rlabel metal3 14721 700 14721 700 0 FrameData_O[3]
rlabel metal2 14364 784 14364 784 0 FrameData_O[4]
rlabel metal2 14420 1036 14420 1036 0 FrameData_O[5]
rlabel metal2 15204 1036 15204 1036 0 FrameData_O[6]
rlabel metal2 15092 1316 15092 1316 0 FrameData_O[7]
rlabel metal3 15057 1820 15057 1820 0 FrameData_O[8]
rlabel metal2 15148 1736 15148 1736 0 FrameData_O[9]
rlabel metal2 1820 763 1820 763 0 FrameStrobe[0]
rlabel metal3 10710 980 10710 980 0 FrameStrobe[10]
rlabel metal2 11396 364 11396 364 0 FrameStrobe[11]
rlabel metal2 9884 259 9884 259 0 FrameStrobe[12]
rlabel metal2 10556 175 10556 175 0 FrameStrobe[13]
rlabel metal2 11228 371 11228 371 0 FrameStrobe[14]
rlabel metal2 11900 371 11900 371 0 FrameStrobe[15]
rlabel metal2 12572 455 12572 455 0 FrameStrobe[16]
rlabel metal2 13244 203 13244 203 0 FrameStrobe[17]
rlabel metal2 13916 63 13916 63 0 FrameStrobe[18]
rlabel metal2 14588 651 14588 651 0 FrameStrobe[19]
rlabel metal2 2492 511 2492 511 0 FrameStrobe[1]
rlabel metal2 3164 63 3164 63 0 FrameStrobe[2]
rlabel metal2 3836 455 3836 455 0 FrameStrobe[3]
rlabel metal2 13692 5236 13692 5236 0 FrameStrobe[4]
rlabel metal2 1764 3164 1764 3164 0 FrameStrobe[5]
rlabel metal2 5852 259 5852 259 0 FrameStrobe[6]
rlabel metal2 6524 315 6524 315 0 FrameStrobe[7]
rlabel metal2 7196 567 7196 567 0 FrameStrobe[8]
rlabel metal2 7868 119 7868 119 0 FrameStrobe[9]
rlabel metal2 10892 6825 10892 6825 0 FrameStrobe_O[0]
rlabel metal2 13580 6020 13580 6020 0 FrameStrobe_O[10]
rlabel metal2 12124 6265 12124 6265 0 FrameStrobe_O[11]
rlabel metal2 14140 6664 14140 6664 0 FrameStrobe_O[12]
rlabel metal2 13524 6104 13524 6104 0 FrameStrobe_O[13]
rlabel metal2 12684 5180 12684 5180 0 FrameStrobe_O[14]
rlabel metal2 14140 6076 14140 6076 0 FrameStrobe_O[15]
rlabel metal2 12684 6629 12684 6629 0 FrameStrobe_O[16]
rlabel metal2 12796 5957 12796 5957 0 FrameStrobe_O[17]
rlabel metal2 12908 6825 12908 6825 0 FrameStrobe_O[18]
rlabel metal2 13468 5180 13468 5180 0 FrameStrobe_O[19]
rlabel metal2 11004 6853 11004 6853 0 FrameStrobe_O[1]
rlabel metal2 11116 6797 11116 6797 0 FrameStrobe_O[2]
rlabel metal2 11228 6433 11228 6433 0 FrameStrobe_O[3]
rlabel metal3 11676 6188 11676 6188 0 FrameStrobe_O[4]
rlabel metal2 11452 6237 11452 6237 0 FrameStrobe_O[5]
rlabel metal2 11564 6937 11564 6937 0 FrameStrobe_O[6]
rlabel metal2 11676 6769 11676 6769 0 FrameStrobe_O[7]
rlabel metal4 12572 6328 12572 6328 0 FrameStrobe_O[8]
rlabel metal2 11900 6825 11900 6825 0 FrameStrobe_O[9]
rlabel metal2 2716 6237 2716 6237 0 N1BEG[0]
rlabel metal2 2828 6545 2828 6545 0 N1BEG[1]
rlabel metal2 2492 5348 2492 5348 0 N1BEG[2]
rlabel metal2 3052 5817 3052 5817 0 N1BEG[3]
rlabel metal3 2128 6580 2128 6580 0 N2BEG[0]
rlabel metal2 2324 5768 2324 5768 0 N2BEG[1]
rlabel metal2 3388 6601 3388 6601 0 N2BEG[2]
rlabel metal2 3108 5488 3108 5488 0 N2BEG[3]
rlabel metal2 3668 4130 3668 4130 0 N2BEG[4]
rlabel metal2 3724 5845 3724 5845 0 N2BEG[5]
rlabel metal2 1876 6692 1876 6692 0 N2BEG[6]
rlabel metal3 3416 5684 3416 5684 0 N2BEG[7]
rlabel metal2 4060 6237 4060 6237 0 N2BEGb[0]
rlabel metal2 3892 5152 3892 5152 0 N2BEGb[1]
rlabel metal2 4340 5152 4340 5152 0 N2BEGb[2]
rlabel metal2 2996 6608 2996 6608 0 N2BEGb[3]
rlabel metal2 3892 5824 3892 5824 0 N2BEGb[4]
rlabel metal3 4508 5404 4508 5404 0 N2BEGb[5]
rlabel metal2 4732 6629 4732 6629 0 N2BEGb[6]
rlabel metal2 4844 6181 4844 6181 0 N2BEGb[7]
rlabel metal2 4956 6013 4956 6013 0 N4BEG[0]
rlabel metal2 6076 6349 6076 6349 0 N4BEG[10]
rlabel metal3 6104 6188 6104 6188 0 N4BEG[11]
rlabel metal3 5992 6580 5992 6580 0 N4BEG[12]
rlabel metal2 6412 6349 6412 6349 0 N4BEG[13]
rlabel metal3 6636 6188 6636 6188 0 N4BEG[14]
rlabel metal2 6636 6825 6636 6825 0 N4BEG[15]
rlabel metal2 3780 6664 3780 6664 0 N4BEG[1]
rlabel metal2 4172 6412 4172 6412 0 N4BEG[2]
rlabel metal2 5292 6825 5292 6825 0 N4BEG[3]
rlabel metal2 5404 6489 5404 6489 0 N4BEG[4]
rlabel metal2 5180 5936 5180 5936 0 N4BEG[5]
rlabel metal2 5628 6629 5628 6629 0 N4BEG[6]
rlabel metal2 5796 5600 5796 5600 0 N4BEG[7]
rlabel metal2 4900 6692 4900 6692 0 N4BEG[8]
rlabel metal2 6580 5376 6580 5376 0 N4BEG[9]
rlabel metal2 2156 4760 2156 4760 0 S1END[0]
rlabel metal2 2604 4032 2604 4032 0 S1END[1]
rlabel metal3 5348 3668 5348 3668 0 S1END[2]
rlabel metal3 5908 4116 5908 4116 0 S1END[3]
rlabel metal2 4088 3332 4088 3332 0 S2END[0]
rlabel metal2 2996 5936 2996 5936 0 S2END[1]
rlabel metal2 7700 6104 7700 6104 0 S2END[2]
rlabel metal2 6580 6692 6580 6692 0 S2END[3]
rlabel metal2 8540 6825 8540 6825 0 S2END[4]
rlabel metal2 8148 6356 8148 6356 0 S2END[5]
rlabel metal2 8596 6300 8596 6300 0 S2END[6]
rlabel metal2 8988 6300 8988 6300 0 S2END[7]
rlabel metal2 5796 4214 5796 4214 0 S2MID[0]
rlabel metal2 7308 6685 7308 6685 0 S2MID[1]
rlabel metal3 6328 4172 6328 4172 0 S2MID[2]
rlabel metal2 6020 5236 6020 5236 0 S2MID[3]
rlabel metal2 6244 4368 6244 4368 0 S2MID[4]
rlabel metal2 4788 6076 4788 6076 0 S2MID[5]
rlabel metal2 7196 5096 7196 5096 0 S2MID[6]
rlabel metal2 7476 5320 7476 5320 0 S2MID[7]
rlabel metal2 6692 4872 6692 4872 0 S4END[0]
rlabel metal2 10108 6041 10108 6041 0 S4END[10]
rlabel metal3 10416 5236 10416 5236 0 S4END[11]
rlabel metal2 11116 5320 11116 5320 0 S4END[12]
rlabel metal2 10444 6993 10444 6993 0 S4END[13]
rlabel metal2 12012 4564 12012 4564 0 S4END[14]
rlabel metal2 14336 5292 14336 5292 0 S4END[15]
rlabel metal2 9100 6769 9100 6769 0 S4END[1]
rlabel metal2 9212 6825 9212 6825 0 S4END[2]
rlabel metal3 9548 6076 9548 6076 0 S4END[3]
rlabel metal3 3164 5292 3164 5292 0 S4END[4]
rlabel metal2 9548 6881 9548 6881 0 S4END[5]
rlabel metal2 9492 6272 9492 6272 0 S4END[6]
rlabel metal3 9408 5292 9408 5292 0 S4END[7]
rlabel metal2 9548 5460 9548 5460 0 S4END[8]
rlabel metal2 9996 6181 9996 6181 0 S4END[9]
rlabel metal2 1148 63 1148 63 0 UserCLK
rlabel metal2 10472 5236 10472 5236 0 UserCLKo
rlabel metal2 13356 1400 13356 1400 0 net1
rlabel metal3 14070 3668 14070 3668 0 net10
rlabel metal2 14700 4536 14700 4536 0 net11
rlabel metal3 10024 588 10024 588 0 net12
rlabel metal2 14756 4704 14756 4704 0 net13
rlabel metal2 14700 5012 14700 5012 0 net14
rlabel metal2 14700 5628 14700 5628 0 net15
rlabel metal2 14028 4340 14028 4340 0 net16
rlabel metal2 13916 4088 13916 4088 0 net17
rlabel metal3 10696 2212 10696 2212 0 net18
rlabel metal3 11144 3388 11144 3388 0 net19
rlabel metal2 14756 2156 14756 2156 0 net2
rlabel metal3 11312 4564 11312 4564 0 net20
rlabel metal2 10052 4928 10052 4928 0 net21
rlabel metal2 10500 5488 10500 5488 0 net22
rlabel metal2 8372 588 8372 588 0 net23
rlabel metal2 10948 5824 10948 5824 0 net24
rlabel metal2 15316 5992 15316 5992 0 net25
rlabel metal3 11620 980 11620 980 0 net26
rlabel metal2 13860 1148 13860 1148 0 net27
rlabel metal2 13916 1176 13916 1176 0 net28
rlabel metal3 11900 1036 11900 1036 0 net29
rlabel metal2 13916 2632 13916 2632 0 net3
rlabel metal3 11956 1148 11956 1148 0 net30
rlabel metal2 13916 1960 13916 1960 0 net31
rlabel metal2 13468 1624 13468 1624 0 net32
rlabel metal3 10304 5908 10304 5908 0 net33
rlabel metal3 12376 3668 12376 3668 0 net34
rlabel metal3 11984 4900 11984 4900 0 net35
rlabel metal2 14140 3122 14140 3122 0 net36
rlabel metal2 12096 1428 12096 1428 0 net37
rlabel metal2 12908 1036 12908 1036 0 net38
rlabel metal2 13860 5488 13860 5488 0 net39
rlabel metal2 8652 2716 8652 2716 0 net4
rlabel metal2 14308 5992 14308 5992 0 net40
rlabel metal2 13580 3360 13580 3360 0 net41
rlabel metal2 14560 4564 14560 4564 0 net42
rlabel metal2 14308 1568 14308 1568 0 net43
rlabel metal2 10052 1302 10052 1302 0 net44
rlabel metal3 11256 1652 11256 1652 0 net45
rlabel metal2 11116 1358 11116 1358 0 net46
rlabel metal3 13132 6020 13132 6020 0 net47
rlabel metal2 1540 5768 1540 5768 0 net48
rlabel metal2 5572 700 5572 700 0 net49
rlabel metal3 11116 2604 11116 2604 0 net5
rlabel metal3 7448 644 7448 644 0 net50
rlabel metal2 6748 2212 6748 2212 0 net51
rlabel metal2 9128 644 9128 644 0 net52
rlabel metal2 2044 4186 2044 4186 0 net53
rlabel metal2 3416 3780 3416 3780 0 net54
rlabel metal2 2324 4186 2324 4186 0 net55
rlabel metal3 2240 4452 2240 4452 0 net56
rlabel metal2 1372 5908 1372 5908 0 net57
rlabel metal2 2604 5180 2604 5180 0 net58
rlabel metal2 4508 5880 4508 5880 0 net59
rlabel metal2 13916 3304 13916 3304 0 net6
rlabel metal2 3332 4452 3332 4452 0 net60
rlabel metal2 4172 4228 4172 4228 0 net61
rlabel metal2 4004 4256 4004 4256 0 net62
rlabel metal2 2156 5852 2156 5852 0 net63
rlabel metal2 3276 4956 3276 4956 0 net64
rlabel metal4 4732 5432 4732 5432 0 net65
rlabel metal3 4186 4900 4186 4900 0 net66
rlabel metal2 4788 4564 4788 4564 0 net67
rlabel metal2 3276 6552 3276 6552 0 net68
rlabel metal2 6300 6048 6300 6048 0 net69
rlabel metal2 7644 3276 7644 3276 0 net7
rlabel metal2 4564 5600 4564 5600 0 net70
rlabel metal2 2772 6188 2772 6188 0 net71
rlabel metal2 3892 3416 3892 3416 0 net72
rlabel metal2 14476 5516 14476 5516 0 net73
rlabel metal2 4116 4172 4116 4172 0 net74
rlabel metal2 2688 5292 2688 5292 0 net75
rlabel metal2 10052 6300 10052 6300 0 net76
rlabel metal2 7140 6076 7140 6076 0 net77
rlabel metal2 8876 6244 8876 6244 0 net78
rlabel metal2 6524 5180 6524 5180 0 net79
rlabel metal2 8036 3696 8036 3696 0 net8
rlabel metal2 3892 5348 3892 5348 0 net80
rlabel metal2 4676 5236 4676 5236 0 net81
rlabel metal2 5348 5376 5348 5376 0 net82
rlabel metal2 10948 5068 10948 5068 0 net83
rlabel metal2 5572 5320 5572 5320 0 net84
rlabel metal2 9828 5684 9828 5684 0 net85
rlabel metal3 7700 5236 7700 5236 0 net86
rlabel metal2 5180 6356 5180 6356 0 net87
rlabel metal2 7028 5404 7028 5404 0 net88
rlabel metal2 10220 896 10220 896 0 net89
rlabel metal2 8484 4284 8484 4284 0 net9
<< properties >>
string FIXED_BBOX 0 0 15848 7112
<< end >>
