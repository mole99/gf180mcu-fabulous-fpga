VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO eFPGA
  CLASS BLOCK ;
  FOREIGN eFPGA ;
  ORIGIN 0.000 0.000 ;
  SIZE 2324.560 BY 3595.760 ;
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3524.080 0.560 3524.640 ;
    END
  END FrameData[0]
  PIN FrameData[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2816.800 1.120 2817.360 ;
    END
  END FrameData[100]
  PIN FrameData[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2821.280 1.120 2821.840 ;
    END
  END FrameData[101]
  PIN FrameData[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2825.760 1.120 2826.320 ;
    END
  END FrameData[102]
  PIN FrameData[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2830.240 1.120 2830.800 ;
    END
  END FrameData[103]
  PIN FrameData[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2834.720 1.120 2835.280 ;
    END
  END FrameData[104]
  PIN FrameData[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2839.200 1.120 2839.760 ;
    END
  END FrameData[105]
  PIN FrameData[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2843.680 1.120 2844.240 ;
    END
  END FrameData[106]
  PIN FrameData[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2848.160 1.120 2848.720 ;
    END
  END FrameData[107]
  PIN FrameData[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2852.640 1.120 2853.200 ;
    END
  END FrameData[108]
  PIN FrameData[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2857.120 1.120 2857.680 ;
    END
  END FrameData[109]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3546.480 0.560 3547.040 ;
    END
  END FrameData[10]
  PIN FrameData[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2861.600 1.120 2862.160 ;
    END
  END FrameData[110]
  PIN FrameData[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2866.080 1.120 2866.640 ;
    END
  END FrameData[111]
  PIN FrameData[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2870.560 1.120 2871.120 ;
    END
  END FrameData[112]
  PIN FrameData[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2875.040 1.120 2875.600 ;
    END
  END FrameData[113]
  PIN FrameData[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2879.520 1.120 2880.080 ;
    END
  END FrameData[114]
  PIN FrameData[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2884.000 1.120 2884.560 ;
    END
  END FrameData[115]
  PIN FrameData[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2888.480 1.120 2889.040 ;
    END
  END FrameData[116]
  PIN FrameData[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2892.960 1.120 2893.520 ;
    END
  END FrameData[117]
  PIN FrameData[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2897.440 1.120 2898.000 ;
    END
  END FrameData[118]
  PIN FrameData[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2901.920 1.120 2902.480 ;
    END
  END FrameData[119]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3548.720 0.560 3549.280 ;
    END
  END FrameData[11]
  PIN FrameData[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2906.400 1.120 2906.960 ;
    END
  END FrameData[120]
  PIN FrameData[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2910.880 1.120 2911.440 ;
    END
  END FrameData[121]
  PIN FrameData[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2915.360 1.120 2915.920 ;
    END
  END FrameData[122]
  PIN FrameData[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2919.840 1.120 2920.400 ;
    END
  END FrameData[123]
  PIN FrameData[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2924.320 1.120 2924.880 ;
    END
  END FrameData[124]
  PIN FrameData[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2928.800 1.120 2929.360 ;
    END
  END FrameData[125]
  PIN FrameData[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2933.280 1.120 2933.840 ;
    END
  END FrameData[126]
  PIN FrameData[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2937.760 1.120 2938.320 ;
    END
  END FrameData[127]
  PIN FrameData[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2511.600 1.120 2512.160 ;
    END
  END FrameData[128]
  PIN FrameData[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2516.080 1.120 2516.640 ;
    END
  END FrameData[129]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3550.960 0.560 3551.520 ;
    END
  END FrameData[12]
  PIN FrameData[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2520.560 1.120 2521.120 ;
    END
  END FrameData[130]
  PIN FrameData[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2525.040 1.120 2525.600 ;
    END
  END FrameData[131]
  PIN FrameData[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2529.520 1.120 2530.080 ;
    END
  END FrameData[132]
  PIN FrameData[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2534.000 1.120 2534.560 ;
    END
  END FrameData[133]
  PIN FrameData[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2538.480 1.120 2539.040 ;
    END
  END FrameData[134]
  PIN FrameData[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2542.960 1.120 2543.520 ;
    END
  END FrameData[135]
  PIN FrameData[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2547.440 1.120 2548.000 ;
    END
  END FrameData[136]
  PIN FrameData[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2551.920 1.120 2552.480 ;
    END
  END FrameData[137]
  PIN FrameData[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2556.400 1.120 2556.960 ;
    END
  END FrameData[138]
  PIN FrameData[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2560.880 1.120 2561.440 ;
    END
  END FrameData[139]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3553.200 0.560 3553.760 ;
    END
  END FrameData[13]
  PIN FrameData[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2565.360 1.120 2565.920 ;
    END
  END FrameData[140]
  PIN FrameData[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2569.840 1.120 2570.400 ;
    END
  END FrameData[141]
  PIN FrameData[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2574.320 1.120 2574.880 ;
    END
  END FrameData[142]
  PIN FrameData[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2578.800 1.120 2579.360 ;
    END
  END FrameData[143]
  PIN FrameData[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2583.280 1.120 2583.840 ;
    END
  END FrameData[144]
  PIN FrameData[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2587.760 1.120 2588.320 ;
    END
  END FrameData[145]
  PIN FrameData[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2592.240 1.120 2592.800 ;
    END
  END FrameData[146]
  PIN FrameData[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2596.720 1.120 2597.280 ;
    END
  END FrameData[147]
  PIN FrameData[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2601.200 1.120 2601.760 ;
    END
  END FrameData[148]
  PIN FrameData[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2605.680 1.120 2606.240 ;
    END
  END FrameData[149]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3555.440 0.560 3556.000 ;
    END
  END FrameData[14]
  PIN FrameData[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2610.160 1.120 2610.720 ;
    END
  END FrameData[150]
  PIN FrameData[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2614.640 1.120 2615.200 ;
    END
  END FrameData[151]
  PIN FrameData[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2619.120 1.120 2619.680 ;
    END
  END FrameData[152]
  PIN FrameData[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2623.600 1.120 2624.160 ;
    END
  END FrameData[153]
  PIN FrameData[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2628.080 1.120 2628.640 ;
    END
  END FrameData[154]
  PIN FrameData[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2632.560 1.120 2633.120 ;
    END
  END FrameData[155]
  PIN FrameData[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2637.040 1.120 2637.600 ;
    END
  END FrameData[156]
  PIN FrameData[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2641.520 1.120 2642.080 ;
    END
  END FrameData[157]
  PIN FrameData[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2646.000 1.120 2646.560 ;
    END
  END FrameData[158]
  PIN FrameData[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2650.480 1.120 2651.040 ;
    END
  END FrameData[159]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3557.680 0.560 3558.240 ;
    END
  END FrameData[15]
  PIN FrameData[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2224.320 1.120 2224.880 ;
    END
  END FrameData[160]
  PIN FrameData[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2228.800 1.120 2229.360 ;
    END
  END FrameData[161]
  PIN FrameData[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2233.280 1.120 2233.840 ;
    END
  END FrameData[162]
  PIN FrameData[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2237.760 1.120 2238.320 ;
    END
  END FrameData[163]
  PIN FrameData[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2242.240 1.120 2242.800 ;
    END
  END FrameData[164]
  PIN FrameData[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2246.720 1.120 2247.280 ;
    END
  END FrameData[165]
  PIN FrameData[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2251.200 1.120 2251.760 ;
    END
  END FrameData[166]
  PIN FrameData[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2255.680 1.120 2256.240 ;
    END
  END FrameData[167]
  PIN FrameData[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2260.160 1.120 2260.720 ;
    END
  END FrameData[168]
  PIN FrameData[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2264.640 1.120 2265.200 ;
    END
  END FrameData[169]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3559.920 0.560 3560.480 ;
    END
  END FrameData[16]
  PIN FrameData[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2269.120 1.120 2269.680 ;
    END
  END FrameData[170]
  PIN FrameData[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2273.600 1.120 2274.160 ;
    END
  END FrameData[171]
  PIN FrameData[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2278.080 1.120 2278.640 ;
    END
  END FrameData[172]
  PIN FrameData[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2282.560 1.120 2283.120 ;
    END
  END FrameData[173]
  PIN FrameData[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2287.040 1.120 2287.600 ;
    END
  END FrameData[174]
  PIN FrameData[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2291.520 1.120 2292.080 ;
    END
  END FrameData[175]
  PIN FrameData[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2296.000 1.120 2296.560 ;
    END
  END FrameData[176]
  PIN FrameData[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2300.480 1.120 2301.040 ;
    END
  END FrameData[177]
  PIN FrameData[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2304.960 1.120 2305.520 ;
    END
  END FrameData[178]
  PIN FrameData[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2309.440 1.120 2310.000 ;
    END
  END FrameData[179]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3562.160 0.560 3562.720 ;
    END
  END FrameData[17]
  PIN FrameData[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2313.920 1.120 2314.480 ;
    END
  END FrameData[180]
  PIN FrameData[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2318.400 1.120 2318.960 ;
    END
  END FrameData[181]
  PIN FrameData[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2322.880 1.120 2323.440 ;
    END
  END FrameData[182]
  PIN FrameData[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2327.360 1.120 2327.920 ;
    END
  END FrameData[183]
  PIN FrameData[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2331.840 1.120 2332.400 ;
    END
  END FrameData[184]
  PIN FrameData[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2336.320 1.120 2336.880 ;
    END
  END FrameData[185]
  PIN FrameData[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2340.800 1.120 2341.360 ;
    END
  END FrameData[186]
  PIN FrameData[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2345.280 1.120 2345.840 ;
    END
  END FrameData[187]
  PIN FrameData[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2349.760 1.120 2350.320 ;
    END
  END FrameData[188]
  PIN FrameData[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2354.240 1.120 2354.800 ;
    END
  END FrameData[189]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3564.400 0.560 3564.960 ;
    END
  END FrameData[18]
  PIN FrameData[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2358.720 1.120 2359.280 ;
    END
  END FrameData[190]
  PIN FrameData[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2363.200 1.120 2363.760 ;
    END
  END FrameData[191]
  PIN FrameData[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1937.040 1.120 1937.600 ;
    END
  END FrameData[192]
  PIN FrameData[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1941.520 1.120 1942.080 ;
    END
  END FrameData[193]
  PIN FrameData[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1946.000 1.120 1946.560 ;
    END
  END FrameData[194]
  PIN FrameData[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1950.480 1.120 1951.040 ;
    END
  END FrameData[195]
  PIN FrameData[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1954.960 1.120 1955.520 ;
    END
  END FrameData[196]
  PIN FrameData[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1959.440 1.120 1960.000 ;
    END
  END FrameData[197]
  PIN FrameData[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1963.920 1.120 1964.480 ;
    END
  END FrameData[198]
  PIN FrameData[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1968.400 1.120 1968.960 ;
    END
  END FrameData[199]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3566.640 0.560 3567.200 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3526.320 0.560 3526.880 ;
    END
  END FrameData[1]
  PIN FrameData[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1972.880 1.120 1973.440 ;
    END
  END FrameData[200]
  PIN FrameData[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1977.360 1.120 1977.920 ;
    END
  END FrameData[201]
  PIN FrameData[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1981.840 1.120 1982.400 ;
    END
  END FrameData[202]
  PIN FrameData[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1986.320 1.120 1986.880 ;
    END
  END FrameData[203]
  PIN FrameData[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1990.800 1.120 1991.360 ;
    END
  END FrameData[204]
  PIN FrameData[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1995.280 1.120 1995.840 ;
    END
  END FrameData[205]
  PIN FrameData[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1999.760 1.120 2000.320 ;
    END
  END FrameData[206]
  PIN FrameData[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2004.240 1.120 2004.800 ;
    END
  END FrameData[207]
  PIN FrameData[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2008.720 1.120 2009.280 ;
    END
  END FrameData[208]
  PIN FrameData[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2013.200 1.120 2013.760 ;
    END
  END FrameData[209]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3568.880 0.560 3569.440 ;
    END
  END FrameData[20]
  PIN FrameData[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2017.680 1.120 2018.240 ;
    END
  END FrameData[210]
  PIN FrameData[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2022.160 1.120 2022.720 ;
    END
  END FrameData[211]
  PIN FrameData[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2026.640 1.120 2027.200 ;
    END
  END FrameData[212]
  PIN FrameData[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2031.120 1.120 2031.680 ;
    END
  END FrameData[213]
  PIN FrameData[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2035.600 1.120 2036.160 ;
    END
  END FrameData[214]
  PIN FrameData[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2040.080 1.120 2040.640 ;
    END
  END FrameData[215]
  PIN FrameData[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2044.560 1.120 2045.120 ;
    END
  END FrameData[216]
  PIN FrameData[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2049.040 1.120 2049.600 ;
    END
  END FrameData[217]
  PIN FrameData[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2053.520 1.120 2054.080 ;
    END
  END FrameData[218]
  PIN FrameData[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2058.000 1.120 2058.560 ;
    END
  END FrameData[219]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3571.120 0.560 3571.680 ;
    END
  END FrameData[21]
  PIN FrameData[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2062.480 1.120 2063.040 ;
    END
  END FrameData[220]
  PIN FrameData[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2066.960 1.120 2067.520 ;
    END
  END FrameData[221]
  PIN FrameData[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2071.440 1.120 2072.000 ;
    END
  END FrameData[222]
  PIN FrameData[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2075.920 1.120 2076.480 ;
    END
  END FrameData[223]
  PIN FrameData[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1649.760 1.120 1650.320 ;
    END
  END FrameData[224]
  PIN FrameData[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1654.240 1.120 1654.800 ;
    END
  END FrameData[225]
  PIN FrameData[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1658.720 1.120 1659.280 ;
    END
  END FrameData[226]
  PIN FrameData[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1663.200 1.120 1663.760 ;
    END
  END FrameData[227]
  PIN FrameData[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1667.680 1.120 1668.240 ;
    END
  END FrameData[228]
  PIN FrameData[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1672.160 1.120 1672.720 ;
    END
  END FrameData[229]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3573.360 0.560 3573.920 ;
    END
  END FrameData[22]
  PIN FrameData[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1676.640 1.120 1677.200 ;
    END
  END FrameData[230]
  PIN FrameData[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1681.120 1.120 1681.680 ;
    END
  END FrameData[231]
  PIN FrameData[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1685.600 1.120 1686.160 ;
    END
  END FrameData[232]
  PIN FrameData[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1690.080 1.120 1690.640 ;
    END
  END FrameData[233]
  PIN FrameData[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1694.560 1.120 1695.120 ;
    END
  END FrameData[234]
  PIN FrameData[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1699.040 1.120 1699.600 ;
    END
  END FrameData[235]
  PIN FrameData[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1703.520 1.120 1704.080 ;
    END
  END FrameData[236]
  PIN FrameData[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1708.000 1.120 1708.560 ;
    END
  END FrameData[237]
  PIN FrameData[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1712.480 1.120 1713.040 ;
    END
  END FrameData[238]
  PIN FrameData[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1716.960 1.120 1717.520 ;
    END
  END FrameData[239]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3575.600 0.560 3576.160 ;
    END
  END FrameData[23]
  PIN FrameData[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1721.440 1.120 1722.000 ;
    END
  END FrameData[240]
  PIN FrameData[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1725.920 1.120 1726.480 ;
    END
  END FrameData[241]
  PIN FrameData[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1730.400 1.120 1730.960 ;
    END
  END FrameData[242]
  PIN FrameData[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1734.880 1.120 1735.440 ;
    END
  END FrameData[243]
  PIN FrameData[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1739.360 1.120 1739.920 ;
    END
  END FrameData[244]
  PIN FrameData[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1743.840 1.120 1744.400 ;
    END
  END FrameData[245]
  PIN FrameData[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1748.320 1.120 1748.880 ;
    END
  END FrameData[246]
  PIN FrameData[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1752.800 1.120 1753.360 ;
    END
  END FrameData[247]
  PIN FrameData[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1757.280 1.120 1757.840 ;
    END
  END FrameData[248]
  PIN FrameData[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1761.760 1.120 1762.320 ;
    END
  END FrameData[249]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3577.840 0.560 3578.400 ;
    END
  END FrameData[24]
  PIN FrameData[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1766.240 1.120 1766.800 ;
    END
  END FrameData[250]
  PIN FrameData[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1770.720 1.120 1771.280 ;
    END
  END FrameData[251]
  PIN FrameData[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1775.200 1.120 1775.760 ;
    END
  END FrameData[252]
  PIN FrameData[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1779.680 1.120 1780.240 ;
    END
  END FrameData[253]
  PIN FrameData[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1784.160 1.120 1784.720 ;
    END
  END FrameData[254]
  PIN FrameData[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1788.640 1.120 1789.200 ;
    END
  END FrameData[255]
  PIN FrameData[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1362.480 1.120 1363.040 ;
    END
  END FrameData[256]
  PIN FrameData[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1366.960 1.120 1367.520 ;
    END
  END FrameData[257]
  PIN FrameData[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1371.440 1.120 1372.000 ;
    END
  END FrameData[258]
  PIN FrameData[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1375.920 1.120 1376.480 ;
    END
  END FrameData[259]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3580.080 0.560 3580.640 ;
    END
  END FrameData[25]
  PIN FrameData[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1380.400 1.120 1380.960 ;
    END
  END FrameData[260]
  PIN FrameData[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1384.880 1.120 1385.440 ;
    END
  END FrameData[261]
  PIN FrameData[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1389.360 1.120 1389.920 ;
    END
  END FrameData[262]
  PIN FrameData[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1393.840 1.120 1394.400 ;
    END
  END FrameData[263]
  PIN FrameData[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1398.320 1.120 1398.880 ;
    END
  END FrameData[264]
  PIN FrameData[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1402.800 1.120 1403.360 ;
    END
  END FrameData[265]
  PIN FrameData[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1407.280 1.120 1407.840 ;
    END
  END FrameData[266]
  PIN FrameData[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1411.760 1.120 1412.320 ;
    END
  END FrameData[267]
  PIN FrameData[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1416.240 1.120 1416.800 ;
    END
  END FrameData[268]
  PIN FrameData[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1420.720 1.120 1421.280 ;
    END
  END FrameData[269]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3582.320 0.560 3582.880 ;
    END
  END FrameData[26]
  PIN FrameData[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1425.200 1.120 1425.760 ;
    END
  END FrameData[270]
  PIN FrameData[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1429.680 1.120 1430.240 ;
    END
  END FrameData[271]
  PIN FrameData[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1434.160 1.120 1434.720 ;
    END
  END FrameData[272]
  PIN FrameData[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1438.640 1.120 1439.200 ;
    END
  END FrameData[273]
  PIN FrameData[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1443.120 1.120 1443.680 ;
    END
  END FrameData[274]
  PIN FrameData[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1447.600 1.120 1448.160 ;
    END
  END FrameData[275]
  PIN FrameData[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1452.080 1.120 1452.640 ;
    END
  END FrameData[276]
  PIN FrameData[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1456.560 1.120 1457.120 ;
    END
  END FrameData[277]
  PIN FrameData[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1461.040 1.120 1461.600 ;
    END
  END FrameData[278]
  PIN FrameData[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1465.520 1.120 1466.080 ;
    END
  END FrameData[279]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3584.560 0.560 3585.120 ;
    END
  END FrameData[27]
  PIN FrameData[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1470.000 1.120 1470.560 ;
    END
  END FrameData[280]
  PIN FrameData[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1474.480 1.120 1475.040 ;
    END
  END FrameData[281]
  PIN FrameData[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1478.960 1.120 1479.520 ;
    END
  END FrameData[282]
  PIN FrameData[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1483.440 1.120 1484.000 ;
    END
  END FrameData[283]
  PIN FrameData[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1487.920 1.120 1488.480 ;
    END
  END FrameData[284]
  PIN FrameData[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1492.400 1.120 1492.960 ;
    END
  END FrameData[285]
  PIN FrameData[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1496.880 1.120 1497.440 ;
    END
  END FrameData[286]
  PIN FrameData[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1501.360 1.120 1501.920 ;
    END
  END FrameData[287]
  PIN FrameData[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1075.200 1.120 1075.760 ;
    END
  END FrameData[288]
  PIN FrameData[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1079.680 1.120 1080.240 ;
    END
  END FrameData[289]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3586.800 0.560 3587.360 ;
    END
  END FrameData[28]
  PIN FrameData[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1084.160 1.120 1084.720 ;
    END
  END FrameData[290]
  PIN FrameData[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1088.640 1.120 1089.200 ;
    END
  END FrameData[291]
  PIN FrameData[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1093.120 1.120 1093.680 ;
    END
  END FrameData[292]
  PIN FrameData[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1097.600 1.120 1098.160 ;
    END
  END FrameData[293]
  PIN FrameData[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1102.080 1.120 1102.640 ;
    END
  END FrameData[294]
  PIN FrameData[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1106.560 1.120 1107.120 ;
    END
  END FrameData[295]
  PIN FrameData[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1111.040 1.120 1111.600 ;
    END
  END FrameData[296]
  PIN FrameData[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1115.520 1.120 1116.080 ;
    END
  END FrameData[297]
  PIN FrameData[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1120.000 1.120 1120.560 ;
    END
  END FrameData[298]
  PIN FrameData[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1124.480 1.120 1125.040 ;
    END
  END FrameData[299]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3589.040 0.560 3589.600 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3528.560 0.560 3529.120 ;
    END
  END FrameData[2]
  PIN FrameData[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1128.960 1.120 1129.520 ;
    END
  END FrameData[300]
  PIN FrameData[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1133.440 1.120 1134.000 ;
    END
  END FrameData[301]
  PIN FrameData[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1137.920 1.120 1138.480 ;
    END
  END FrameData[302]
  PIN FrameData[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1142.400 1.120 1142.960 ;
    END
  END FrameData[303]
  PIN FrameData[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1146.880 1.120 1147.440 ;
    END
  END FrameData[304]
  PIN FrameData[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1151.360 1.120 1151.920 ;
    END
  END FrameData[305]
  PIN FrameData[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1155.840 1.120 1156.400 ;
    END
  END FrameData[306]
  PIN FrameData[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1160.320 1.120 1160.880 ;
    END
  END FrameData[307]
  PIN FrameData[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1164.800 1.120 1165.360 ;
    END
  END FrameData[308]
  PIN FrameData[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1169.280 1.120 1169.840 ;
    END
  END FrameData[309]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3591.280 0.560 3591.840 ;
    END
  END FrameData[30]
  PIN FrameData[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1173.760 1.120 1174.320 ;
    END
  END FrameData[310]
  PIN FrameData[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1178.240 1.120 1178.800 ;
    END
  END FrameData[311]
  PIN FrameData[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1182.720 1.120 1183.280 ;
    END
  END FrameData[312]
  PIN FrameData[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1187.200 1.120 1187.760 ;
    END
  END FrameData[313]
  PIN FrameData[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1191.680 1.120 1192.240 ;
    END
  END FrameData[314]
  PIN FrameData[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1196.160 1.120 1196.720 ;
    END
  END FrameData[315]
  PIN FrameData[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1200.640 1.120 1201.200 ;
    END
  END FrameData[316]
  PIN FrameData[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1205.120 1.120 1205.680 ;
    END
  END FrameData[317]
  PIN FrameData[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1209.600 1.120 1210.160 ;
    END
  END FrameData[318]
  PIN FrameData[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1214.080 1.120 1214.640 ;
    END
  END FrameData[319]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3593.520 0.560 3594.080 ;
    END
  END FrameData[31]
  PIN FrameData[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 787.920 1.120 788.480 ;
    END
  END FrameData[320]
  PIN FrameData[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 792.400 1.120 792.960 ;
    END
  END FrameData[321]
  PIN FrameData[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 796.880 1.120 797.440 ;
    END
  END FrameData[322]
  PIN FrameData[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 801.360 1.120 801.920 ;
    END
  END FrameData[323]
  PIN FrameData[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 805.840 1.120 806.400 ;
    END
  END FrameData[324]
  PIN FrameData[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 810.320 1.120 810.880 ;
    END
  END FrameData[325]
  PIN FrameData[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 814.800 1.120 815.360 ;
    END
  END FrameData[326]
  PIN FrameData[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 819.280 1.120 819.840 ;
    END
  END FrameData[327]
  PIN FrameData[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 823.760 1.120 824.320 ;
    END
  END FrameData[328]
  PIN FrameData[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 828.240 1.120 828.800 ;
    END
  END FrameData[329]
  PIN FrameData[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3373.440 1.120 3374.000 ;
    END
  END FrameData[32]
  PIN FrameData[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 832.720 1.120 833.280 ;
    END
  END FrameData[330]
  PIN FrameData[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 837.200 1.120 837.760 ;
    END
  END FrameData[331]
  PIN FrameData[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 841.680 1.120 842.240 ;
    END
  END FrameData[332]
  PIN FrameData[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 846.160 1.120 846.720 ;
    END
  END FrameData[333]
  PIN FrameData[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 850.640 1.120 851.200 ;
    END
  END FrameData[334]
  PIN FrameData[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 855.120 1.120 855.680 ;
    END
  END FrameData[335]
  PIN FrameData[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 859.600 1.120 860.160 ;
    END
  END FrameData[336]
  PIN FrameData[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 864.080 1.120 864.640 ;
    END
  END FrameData[337]
  PIN FrameData[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 868.560 1.120 869.120 ;
    END
  END FrameData[338]
  PIN FrameData[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 873.040 1.120 873.600 ;
    END
  END FrameData[339]
  PIN FrameData[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3377.920 1.120 3378.480 ;
    END
  END FrameData[33]
  PIN FrameData[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 877.520 1.120 878.080 ;
    END
  END FrameData[340]
  PIN FrameData[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 882.000 1.120 882.560 ;
    END
  END FrameData[341]
  PIN FrameData[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 886.480 1.120 887.040 ;
    END
  END FrameData[342]
  PIN FrameData[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 890.960 1.120 891.520 ;
    END
  END FrameData[343]
  PIN FrameData[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 895.440 1.120 896.000 ;
    END
  END FrameData[344]
  PIN FrameData[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 899.920 1.120 900.480 ;
    END
  END FrameData[345]
  PIN FrameData[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 904.400 1.120 904.960 ;
    END
  END FrameData[346]
  PIN FrameData[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 908.880 1.120 909.440 ;
    END
  END FrameData[347]
  PIN FrameData[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 913.360 1.120 913.920 ;
    END
  END FrameData[348]
  PIN FrameData[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 917.840 1.120 918.400 ;
    END
  END FrameData[349]
  PIN FrameData[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3382.400 1.120 3382.960 ;
    END
  END FrameData[34]
  PIN FrameData[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 922.320 1.120 922.880 ;
    END
  END FrameData[350]
  PIN FrameData[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 926.800 1.120 927.360 ;
    END
  END FrameData[351]
  PIN FrameData[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 500.640 1.120 501.200 ;
    END
  END FrameData[352]
  PIN FrameData[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 505.120 1.120 505.680 ;
    END
  END FrameData[353]
  PIN FrameData[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 509.600 1.120 510.160 ;
    END
  END FrameData[354]
  PIN FrameData[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 514.080 1.120 514.640 ;
    END
  END FrameData[355]
  PIN FrameData[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 518.560 1.120 519.120 ;
    END
  END FrameData[356]
  PIN FrameData[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 523.040 1.120 523.600 ;
    END
  END FrameData[357]
  PIN FrameData[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 527.520 1.120 528.080 ;
    END
  END FrameData[358]
  PIN FrameData[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 532.000 1.120 532.560 ;
    END
  END FrameData[359]
  PIN FrameData[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3386.880 1.120 3387.440 ;
    END
  END FrameData[35]
  PIN FrameData[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 536.480 1.120 537.040 ;
    END
  END FrameData[360]
  PIN FrameData[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 540.960 1.120 541.520 ;
    END
  END FrameData[361]
  PIN FrameData[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 545.440 1.120 546.000 ;
    END
  END FrameData[362]
  PIN FrameData[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 549.920 1.120 550.480 ;
    END
  END FrameData[363]
  PIN FrameData[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 554.400 1.120 554.960 ;
    END
  END FrameData[364]
  PIN FrameData[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 558.880 1.120 559.440 ;
    END
  END FrameData[365]
  PIN FrameData[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 563.360 1.120 563.920 ;
    END
  END FrameData[366]
  PIN FrameData[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 567.840 1.120 568.400 ;
    END
  END FrameData[367]
  PIN FrameData[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 572.320 1.120 572.880 ;
    END
  END FrameData[368]
  PIN FrameData[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 576.800 1.120 577.360 ;
    END
  END FrameData[369]
  PIN FrameData[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3391.360 1.120 3391.920 ;
    END
  END FrameData[36]
  PIN FrameData[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 581.280 1.120 581.840 ;
    END
  END FrameData[370]
  PIN FrameData[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 585.760 1.120 586.320 ;
    END
  END FrameData[371]
  PIN FrameData[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 590.240 1.120 590.800 ;
    END
  END FrameData[372]
  PIN FrameData[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 594.720 1.120 595.280 ;
    END
  END FrameData[373]
  PIN FrameData[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 599.200 1.120 599.760 ;
    END
  END FrameData[374]
  PIN FrameData[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 603.680 1.120 604.240 ;
    END
  END FrameData[375]
  PIN FrameData[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 608.160 1.120 608.720 ;
    END
  END FrameData[376]
  PIN FrameData[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 612.640 1.120 613.200 ;
    END
  END FrameData[377]
  PIN FrameData[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 617.120 1.120 617.680 ;
    END
  END FrameData[378]
  PIN FrameData[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 621.600 1.120 622.160 ;
    END
  END FrameData[379]
  PIN FrameData[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3395.840 1.120 3396.400 ;
    END
  END FrameData[37]
  PIN FrameData[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 626.080 1.120 626.640 ;
    END
  END FrameData[380]
  PIN FrameData[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 630.560 1.120 631.120 ;
    END
  END FrameData[381]
  PIN FrameData[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 635.040 1.120 635.600 ;
    END
  END FrameData[382]
  PIN FrameData[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 639.520 1.120 640.080 ;
    END
  END FrameData[383]
  PIN FrameData[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 213.360 1.120 213.920 ;
    END
  END FrameData[384]
  PIN FrameData[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 217.840 1.120 218.400 ;
    END
  END FrameData[385]
  PIN FrameData[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 222.320 1.120 222.880 ;
    END
  END FrameData[386]
  PIN FrameData[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 226.800 1.120 227.360 ;
    END
  END FrameData[387]
  PIN FrameData[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 231.280 1.120 231.840 ;
    END
  END FrameData[388]
  PIN FrameData[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 235.760 1.120 236.320 ;
    END
  END FrameData[389]
  PIN FrameData[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3400.320 1.120 3400.880 ;
    END
  END FrameData[38]
  PIN FrameData[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 240.240 1.120 240.800 ;
    END
  END FrameData[390]
  PIN FrameData[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 244.720 1.120 245.280 ;
    END
  END FrameData[391]
  PIN FrameData[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 249.200 1.120 249.760 ;
    END
  END FrameData[392]
  PIN FrameData[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 253.680 1.120 254.240 ;
    END
  END FrameData[393]
  PIN FrameData[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 258.160 1.120 258.720 ;
    END
  END FrameData[394]
  PIN FrameData[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.640 1.120 263.200 ;
    END
  END FrameData[395]
  PIN FrameData[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 267.120 1.120 267.680 ;
    END
  END FrameData[396]
  PIN FrameData[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 271.600 1.120 272.160 ;
    END
  END FrameData[397]
  PIN FrameData[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 276.080 1.120 276.640 ;
    END
  END FrameData[398]
  PIN FrameData[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 280.560 1.120 281.120 ;
    END
  END FrameData[399]
  PIN FrameData[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3404.800 1.120 3405.360 ;
    END
  END FrameData[39]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3530.800 0.560 3531.360 ;
    END
  END FrameData[3]
  PIN FrameData[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.040 1.120 285.600 ;
    END
  END FrameData[400]
  PIN FrameData[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 289.520 1.120 290.080 ;
    END
  END FrameData[401]
  PIN FrameData[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 1.120 294.560 ;
    END
  END FrameData[402]
  PIN FrameData[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 298.480 1.120 299.040 ;
    END
  END FrameData[403]
  PIN FrameData[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.960 1.120 303.520 ;
    END
  END FrameData[404]
  PIN FrameData[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 307.440 1.120 308.000 ;
    END
  END FrameData[405]
  PIN FrameData[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 311.920 1.120 312.480 ;
    END
  END FrameData[406]
  PIN FrameData[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 316.400 1.120 316.960 ;
    END
  END FrameData[407]
  PIN FrameData[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 320.880 1.120 321.440 ;
    END
  END FrameData[408]
  PIN FrameData[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 325.360 1.120 325.920 ;
    END
  END FrameData[409]
  PIN FrameData[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3409.280 1.120 3409.840 ;
    END
  END FrameData[40]
  PIN FrameData[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 329.840 1.120 330.400 ;
    END
  END FrameData[410]
  PIN FrameData[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.320 1.120 334.880 ;
    END
  END FrameData[411]
  PIN FrameData[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 338.800 1.120 339.360 ;
    END
  END FrameData[412]
  PIN FrameData[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 343.280 1.120 343.840 ;
    END
  END FrameData[413]
  PIN FrameData[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 347.760 1.120 348.320 ;
    END
  END FrameData[414]
  PIN FrameData[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 352.240 1.120 352.800 ;
    END
  END FrameData[415]
  PIN FrameData[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 5.600 0.560 6.160 ;
    END
  END FrameData[416]
  PIN FrameData[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 7.840 0.560 8.400 ;
    END
  END FrameData[417]
  PIN FrameData[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 10.080 0.560 10.640 ;
    END
  END FrameData[418]
  PIN FrameData[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 12.320 0.560 12.880 ;
    END
  END FrameData[419]
  PIN FrameData[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3413.760 1.120 3414.320 ;
    END
  END FrameData[41]
  PIN FrameData[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 14.560 0.560 15.120 ;
    END
  END FrameData[420]
  PIN FrameData[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 16.800 0.560 17.360 ;
    END
  END FrameData[421]
  PIN FrameData[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.040 0.560 19.600 ;
    END
  END FrameData[422]
  PIN FrameData[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 21.280 0.560 21.840 ;
    END
  END FrameData[423]
  PIN FrameData[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.520 0.560 24.080 ;
    END
  END FrameData[424]
  PIN FrameData[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 25.760 0.560 26.320 ;
    END
  END FrameData[425]
  PIN FrameData[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 28.000 0.560 28.560 ;
    END
  END FrameData[426]
  PIN FrameData[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.240 0.560 30.800 ;
    END
  END FrameData[427]
  PIN FrameData[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 32.480 0.560 33.040 ;
    END
  END FrameData[428]
  PIN FrameData[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 34.720 0.560 35.280 ;
    END
  END FrameData[429]
  PIN FrameData[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3418.240 1.120 3418.800 ;
    END
  END FrameData[42]
  PIN FrameData[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 36.960 0.560 37.520 ;
    END
  END FrameData[430]
  PIN FrameData[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.200 0.560 39.760 ;
    END
  END FrameData[431]
  PIN FrameData[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 41.440 0.560 42.000 ;
    END
  END FrameData[432]
  PIN FrameData[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.680 0.560 44.240 ;
    END
  END FrameData[433]
  PIN FrameData[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 45.920 0.560 46.480 ;
    END
  END FrameData[434]
  PIN FrameData[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.160 0.560 48.720 ;
    END
  END FrameData[435]
  PIN FrameData[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.400 0.560 50.960 ;
    END
  END FrameData[436]
  PIN FrameData[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 52.640 0.560 53.200 ;
    END
  END FrameData[437]
  PIN FrameData[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 54.880 0.560 55.440 ;
    END
  END FrameData[438]
  PIN FrameData[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 0.560 57.680 ;
    END
  END FrameData[439]
  PIN FrameData[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3422.720 1.120 3423.280 ;
    END
  END FrameData[43]
  PIN FrameData[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.360 0.560 59.920 ;
    END
  END FrameData[440]
  PIN FrameData[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.600 0.560 62.160 ;
    END
  END FrameData[441]
  PIN FrameData[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 63.840 0.560 64.400 ;
    END
  END FrameData[442]
  PIN FrameData[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.080 0.560 66.640 ;
    END
  END FrameData[443]
  PIN FrameData[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 68.320 0.560 68.880 ;
    END
  END FrameData[444]
  PIN FrameData[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.560 0.560 71.120 ;
    END
  END FrameData[445]
  PIN FrameData[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 72.800 0.560 73.360 ;
    END
  END FrameData[446]
  PIN FrameData[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.654000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 75.040 0.560 75.600 ;
    END
  END FrameData[447]
  PIN FrameData[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3427.200 1.120 3427.760 ;
    END
  END FrameData[44]
  PIN FrameData[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3431.680 1.120 3432.240 ;
    END
  END FrameData[45]
  PIN FrameData[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3436.160 1.120 3436.720 ;
    END
  END FrameData[46]
  PIN FrameData[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3440.640 1.120 3441.200 ;
    END
  END FrameData[47]
  PIN FrameData[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3445.120 1.120 3445.680 ;
    END
  END FrameData[48]
  PIN FrameData[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3449.600 1.120 3450.160 ;
    END
  END FrameData[49]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3533.040 0.560 3533.600 ;
    END
  END FrameData[4]
  PIN FrameData[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3454.080 1.120 3454.640 ;
    END
  END FrameData[50]
  PIN FrameData[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3458.560 1.120 3459.120 ;
    END
  END FrameData[51]
  PIN FrameData[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3463.040 1.120 3463.600 ;
    END
  END FrameData[52]
  PIN FrameData[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3467.520 1.120 3468.080 ;
    END
  END FrameData[53]
  PIN FrameData[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3472.000 1.120 3472.560 ;
    END
  END FrameData[54]
  PIN FrameData[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3476.480 1.120 3477.040 ;
    END
  END FrameData[55]
  PIN FrameData[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3480.960 1.120 3481.520 ;
    END
  END FrameData[56]
  PIN FrameData[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3485.440 1.120 3486.000 ;
    END
  END FrameData[57]
  PIN FrameData[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3489.920 1.120 3490.480 ;
    END
  END FrameData[58]
  PIN FrameData[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3494.400 1.120 3494.960 ;
    END
  END FrameData[59]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3535.280 0.560 3535.840 ;
    END
  END FrameData[5]
  PIN FrameData[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3498.880 1.120 3499.440 ;
    END
  END FrameData[60]
  PIN FrameData[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3503.360 1.120 3503.920 ;
    END
  END FrameData[61]
  PIN FrameData[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3507.840 1.120 3508.400 ;
    END
  END FrameData[62]
  PIN FrameData[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3512.320 1.120 3512.880 ;
    END
  END FrameData[63]
  PIN FrameData[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3086.160 1.120 3086.720 ;
    END
  END FrameData[64]
  PIN FrameData[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3090.640 1.120 3091.200 ;
    END
  END FrameData[65]
  PIN FrameData[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3095.120 1.120 3095.680 ;
    END
  END FrameData[66]
  PIN FrameData[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3099.600 1.120 3100.160 ;
    END
  END FrameData[67]
  PIN FrameData[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3104.080 1.120 3104.640 ;
    END
  END FrameData[68]
  PIN FrameData[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3108.560 1.120 3109.120 ;
    END
  END FrameData[69]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3537.520 0.560 3538.080 ;
    END
  END FrameData[6]
  PIN FrameData[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3113.040 1.120 3113.600 ;
    END
  END FrameData[70]
  PIN FrameData[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3117.520 1.120 3118.080 ;
    END
  END FrameData[71]
  PIN FrameData[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3122.000 1.120 3122.560 ;
    END
  END FrameData[72]
  PIN FrameData[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3126.480 1.120 3127.040 ;
    END
  END FrameData[73]
  PIN FrameData[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3130.960 1.120 3131.520 ;
    END
  END FrameData[74]
  PIN FrameData[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3135.440 1.120 3136.000 ;
    END
  END FrameData[75]
  PIN FrameData[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3139.920 1.120 3140.480 ;
    END
  END FrameData[76]
  PIN FrameData[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3144.400 1.120 3144.960 ;
    END
  END FrameData[77]
  PIN FrameData[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3148.880 1.120 3149.440 ;
    END
  END FrameData[78]
  PIN FrameData[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3153.360 1.120 3153.920 ;
    END
  END FrameData[79]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3539.760 0.560 3540.320 ;
    END
  END FrameData[7]
  PIN FrameData[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3157.840 1.120 3158.400 ;
    END
  END FrameData[80]
  PIN FrameData[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3162.320 1.120 3162.880 ;
    END
  END FrameData[81]
  PIN FrameData[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3166.800 1.120 3167.360 ;
    END
  END FrameData[82]
  PIN FrameData[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3171.280 1.120 3171.840 ;
    END
  END FrameData[83]
  PIN FrameData[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3175.760 1.120 3176.320 ;
    END
  END FrameData[84]
  PIN FrameData[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3180.240 1.120 3180.800 ;
    END
  END FrameData[85]
  PIN FrameData[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3184.720 1.120 3185.280 ;
    END
  END FrameData[86]
  PIN FrameData[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3189.200 1.120 3189.760 ;
    END
  END FrameData[87]
  PIN FrameData[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3193.680 1.120 3194.240 ;
    END
  END FrameData[88]
  PIN FrameData[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3198.160 1.120 3198.720 ;
    END
  END FrameData[89]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3542.000 0.560 3542.560 ;
    END
  END FrameData[8]
  PIN FrameData[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3202.640 1.120 3203.200 ;
    END
  END FrameData[90]
  PIN FrameData[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3207.120 1.120 3207.680 ;
    END
  END FrameData[91]
  PIN FrameData[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3211.600 1.120 3212.160 ;
    END
  END FrameData[92]
  PIN FrameData[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3216.080 1.120 3216.640 ;
    END
  END FrameData[93]
  PIN FrameData[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3220.560 1.120 3221.120 ;
    END
  END FrameData[94]
  PIN FrameData[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.862000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3225.040 1.120 3225.600 ;
    END
  END FrameData[95]
  PIN FrameData[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2798.880 1.120 2799.440 ;
    END
  END FrameData[96]
  PIN FrameData[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2803.360 1.120 2803.920 ;
    END
  END FrameData[97]
  PIN FrameData[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2807.840 1.120 2808.400 ;
    END
  END FrameData[98]
  PIN FrameData[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.310000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2812.320 1.120 2812.880 ;
    END
  END FrameData[99]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3544.240 0.560 3544.800 ;
    END
  END FrameData[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.640 0.000 11.200 0.560 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1349.600 0.000 1350.160 0.560 ;
    END
  END FrameStrobe[100]
  PIN FrameStrobe[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1363.040 0.000 1363.600 0.560 ;
    END
  END FrameStrobe[101]
  PIN FrameStrobe[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1376.480 0.000 1377.040 0.560 ;
    END
  END FrameStrobe[102]
  PIN FrameStrobe[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1389.920 0.000 1390.480 0.560 ;
    END
  END FrameStrobe[103]
  PIN FrameStrobe[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1403.360 0.000 1403.920 0.560 ;
    END
  END FrameStrobe[104]
  PIN FrameStrobe[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1416.800 0.000 1417.360 0.560 ;
    END
  END FrameStrobe[105]
  PIN FrameStrobe[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1430.240 0.000 1430.800 0.560 ;
    END
  END FrameStrobe[106]
  PIN FrameStrobe[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1443.680 0.000 1444.240 0.560 ;
    END
  END FrameStrobe[107]
  PIN FrameStrobe[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1457.120 0.000 1457.680 0.560 ;
    END
  END FrameStrobe[108]
  PIN FrameStrobe[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1470.560 0.000 1471.120 0.560 ;
    END
  END FrameStrobe[109]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 77.840 0.000 78.400 0.560 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1484.000 0.000 1484.560 0.560 ;
    END
  END FrameStrobe[110]
  PIN FrameStrobe[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1497.440 0.000 1498.000 0.560 ;
    END
  END FrameStrobe[111]
  PIN FrameStrobe[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1510.880 0.000 1511.440 0.560 ;
    END
  END FrameStrobe[112]
  PIN FrameStrobe[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1524.320 0.000 1524.880 0.560 ;
    END
  END FrameStrobe[113]
  PIN FrameStrobe[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1537.760 0.000 1538.320 0.560 ;
    END
  END FrameStrobe[114]
  PIN FrameStrobe[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1551.200 0.000 1551.760 0.560 ;
    END
  END FrameStrobe[115]
  PIN FrameStrobe[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1564.640 0.000 1565.200 0.560 ;
    END
  END FrameStrobe[116]
  PIN FrameStrobe[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1578.080 0.000 1578.640 0.560 ;
    END
  END FrameStrobe[117]
  PIN FrameStrobe[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1591.520 0.000 1592.080 0.560 ;
    END
  END FrameStrobe[118]
  PIN FrameStrobe[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1604.960 0.000 1605.520 0.560 ;
    END
  END FrameStrobe[119]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 84.560 0.000 85.120 0.560 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1634.640 0.000 1635.200 0.560 ;
    END
  END FrameStrobe[120]
  PIN FrameStrobe[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1646.960 0.000 1647.520 0.560 ;
    END
  END FrameStrobe[121]
  PIN FrameStrobe[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1659.280 0.000 1659.840 0.560 ;
    END
  END FrameStrobe[122]
  PIN FrameStrobe[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1671.600 0.000 1672.160 0.560 ;
    END
  END FrameStrobe[123]
  PIN FrameStrobe[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1683.920 0.000 1684.480 0.560 ;
    END
  END FrameStrobe[124]
  PIN FrameStrobe[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1696.240 0.000 1696.800 0.560 ;
    END
  END FrameStrobe[125]
  PIN FrameStrobe[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1708.560 0.000 1709.120 0.560 ;
    END
  END FrameStrobe[126]
  PIN FrameStrobe[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1720.880 0.000 1721.440 0.560 ;
    END
  END FrameStrobe[127]
  PIN FrameStrobe[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1733.200 0.000 1733.760 0.560 ;
    END
  END FrameStrobe[128]
  PIN FrameStrobe[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1745.520 0.000 1746.080 0.560 ;
    END
  END FrameStrobe[129]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 91.280 0.000 91.840 0.560 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1757.840 0.000 1758.400 0.560 ;
    END
  END FrameStrobe[130]
  PIN FrameStrobe[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1770.160 0.000 1770.720 0.560 ;
    END
  END FrameStrobe[131]
  PIN FrameStrobe[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1782.480 0.000 1783.040 0.560 ;
    END
  END FrameStrobe[132]
  PIN FrameStrobe[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1794.800 0.000 1795.360 0.560 ;
    END
  END FrameStrobe[133]
  PIN FrameStrobe[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1807.120 0.000 1807.680 0.560 ;
    END
  END FrameStrobe[134]
  PIN FrameStrobe[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1819.440 0.000 1820.000 0.560 ;
    END
  END FrameStrobe[135]
  PIN FrameStrobe[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1831.760 0.000 1832.320 0.560 ;
    END
  END FrameStrobe[136]
  PIN FrameStrobe[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1844.080 0.000 1844.640 0.560 ;
    END
  END FrameStrobe[137]
  PIN FrameStrobe[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1856.400 0.000 1856.960 0.560 ;
    END
  END FrameStrobe[138]
  PIN FrameStrobe[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1868.720 0.000 1869.280 0.560 ;
    END
  END FrameStrobe[139]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 98.000 0.000 98.560 0.560 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1900.640 0.000 1901.200 0.560 ;
    END
  END FrameStrobe[140]
  PIN FrameStrobe[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1914.080 0.000 1914.640 0.560 ;
    END
  END FrameStrobe[141]
  PIN FrameStrobe[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1927.520 0.000 1928.080 0.560 ;
    END
  END FrameStrobe[142]
  PIN FrameStrobe[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1940.960 0.000 1941.520 0.560 ;
    END
  END FrameStrobe[143]
  PIN FrameStrobe[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1954.400 0.000 1954.960 0.560 ;
    END
  END FrameStrobe[144]
  PIN FrameStrobe[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1967.840 0.000 1968.400 0.560 ;
    END
  END FrameStrobe[145]
  PIN FrameStrobe[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1981.280 0.000 1981.840 0.560 ;
    END
  END FrameStrobe[146]
  PIN FrameStrobe[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1994.720 0.000 1995.280 0.560 ;
    END
  END FrameStrobe[147]
  PIN FrameStrobe[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2008.160 0.000 2008.720 0.560 ;
    END
  END FrameStrobe[148]
  PIN FrameStrobe[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2021.600 0.000 2022.160 0.560 ;
    END
  END FrameStrobe[149]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 104.720 0.000 105.280 0.560 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2035.040 0.000 2035.600 0.560 ;
    END
  END FrameStrobe[150]
  PIN FrameStrobe[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2048.480 0.000 2049.040 0.560 ;
    END
  END FrameStrobe[151]
  PIN FrameStrobe[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2061.920 0.000 2062.480 0.560 ;
    END
  END FrameStrobe[152]
  PIN FrameStrobe[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2075.360 0.000 2075.920 0.560 ;
    END
  END FrameStrobe[153]
  PIN FrameStrobe[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2088.800 0.000 2089.360 0.560 ;
    END
  END FrameStrobe[154]
  PIN FrameStrobe[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2102.240 0.000 2102.800 0.560 ;
    END
  END FrameStrobe[155]
  PIN FrameStrobe[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2115.680 0.000 2116.240 0.560 ;
    END
  END FrameStrobe[156]
  PIN FrameStrobe[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2129.120 0.000 2129.680 0.560 ;
    END
  END FrameStrobe[157]
  PIN FrameStrobe[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2142.560 0.000 2143.120 0.560 ;
    END
  END FrameStrobe[158]
  PIN FrameStrobe[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2156.000 0.000 2156.560 0.560 ;
    END
  END FrameStrobe[159]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 111.440 0.000 112.000 0.560 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2183.440 0.000 2184.000 0.560 ;
    END
  END FrameStrobe[160]
  PIN FrameStrobe[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2190.160 0.000 2190.720 0.560 ;
    END
  END FrameStrobe[161]
  PIN FrameStrobe[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2196.880 0.000 2197.440 0.560 ;
    END
  END FrameStrobe[162]
  PIN FrameStrobe[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2203.600 0.000 2204.160 0.560 ;
    END
  END FrameStrobe[163]
  PIN FrameStrobe[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2210.320 0.000 2210.880 0.560 ;
    END
  END FrameStrobe[164]
  PIN FrameStrobe[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2217.040 0.000 2217.600 0.560 ;
    END
  END FrameStrobe[165]
  PIN FrameStrobe[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2223.760 0.000 2224.320 0.560 ;
    END
  END FrameStrobe[166]
  PIN FrameStrobe[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2230.480 0.000 2231.040 0.560 ;
    END
  END FrameStrobe[167]
  PIN FrameStrobe[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2241.120 0.000 2241.680 0.560 ;
    END
  END FrameStrobe[168]
  PIN FrameStrobe[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2243.920 0.000 2244.480 0.560 ;
    END
  END FrameStrobe[169]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 118.160 0.000 118.720 0.560 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2250.640 0.000 2251.200 0.560 ;
    END
  END FrameStrobe[170]
  PIN FrameStrobe[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2257.360 0.000 2257.920 0.560 ;
    END
  END FrameStrobe[171]
  PIN FrameStrobe[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2264.080 0.000 2264.640 0.560 ;
    END
  END FrameStrobe[172]
  PIN FrameStrobe[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2270.800 0.000 2271.360 0.560 ;
    END
  END FrameStrobe[173]
  PIN FrameStrobe[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2277.520 0.000 2278.080 0.560 ;
    END
  END FrameStrobe[174]
  PIN FrameStrobe[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2284.240 0.000 2284.800 0.560 ;
    END
  END FrameStrobe[175]
  PIN FrameStrobe[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2290.960 0.000 2291.520 0.560 ;
    END
  END FrameStrobe[176]
  PIN FrameStrobe[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2297.680 0.000 2298.240 0.560 ;
    END
  END FrameStrobe[177]
  PIN FrameStrobe[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2304.400 0.000 2304.960 0.560 ;
    END
  END FrameStrobe[178]
  PIN FrameStrobe[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2311.120 0.000 2311.680 0.560 ;
    END
  END FrameStrobe[179]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 124.880 0.000 125.440 0.560 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 131.600 0.000 132.160 0.560 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 138.320 0.000 138.880 0.560 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 17.360 0.000 17.920 0.560 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 230.720 0.000 231.280 0.560 ;
    END
  END FrameStrobe[20]
  PIN FrameStrobe[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 240.800 0.000 241.360 0.560 ;
    END
  END FrameStrobe[21]
  PIN FrameStrobe[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 250.880 0.000 251.440 0.560 ;
    END
  END FrameStrobe[22]
  PIN FrameStrobe[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 0.000 261.520 0.560 ;
    END
  END FrameStrobe[23]
  PIN FrameStrobe[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 271.040 0.000 271.600 0.560 ;
    END
  END FrameStrobe[24]
  PIN FrameStrobe[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 0.000 281.680 0.560 ;
    END
  END FrameStrobe[25]
  PIN FrameStrobe[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 291.200 0.000 291.760 0.560 ;
    END
  END FrameStrobe[26]
  PIN FrameStrobe[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 301.280 0.000 301.840 0.560 ;
    END
  END FrameStrobe[27]
  PIN FrameStrobe[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 311.360 0.000 311.920 0.560 ;
    END
  END FrameStrobe[28]
  PIN FrameStrobe[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 321.440 0.000 322.000 0.560 ;
    END
  END FrameStrobe[29]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 24.080 0.000 24.640 0.560 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 331.520 0.000 332.080 0.560 ;
    END
  END FrameStrobe[30]
  PIN FrameStrobe[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 341.600 0.000 342.160 0.560 ;
    END
  END FrameStrobe[31]
  PIN FrameStrobe[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 351.680 0.000 352.240 0.560 ;
    END
  END FrameStrobe[32]
  PIN FrameStrobe[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 361.760 0.000 362.320 0.560 ;
    END
  END FrameStrobe[33]
  PIN FrameStrobe[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 371.840 0.000 372.400 0.560 ;
    END
  END FrameStrobe[34]
  PIN FrameStrobe[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 381.920 0.000 382.480 0.560 ;
    END
  END FrameStrobe[35]
  PIN FrameStrobe[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 392.000 0.000 392.560 0.560 ;
    END
  END FrameStrobe[36]
  PIN FrameStrobe[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 402.080 0.000 402.640 0.560 ;
    END
  END FrameStrobe[37]
  PIN FrameStrobe[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 412.160 0.000 412.720 0.560 ;
    END
  END FrameStrobe[38]
  PIN FrameStrobe[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 422.240 0.000 422.800 0.560 ;
    END
  END FrameStrobe[39]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.510000 ;
    PORT
      LAYER Metal2 ;
        RECT 30.800 0.000 31.360 0.560 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 453.040 0.000 453.600 0.560 ;
    END
  END FrameStrobe[40]
  PIN FrameStrobe[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 466.480 0.000 467.040 0.560 ;
    END
  END FrameStrobe[41]
  PIN FrameStrobe[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 479.920 0.000 480.480 0.560 ;
    END
  END FrameStrobe[42]
  PIN FrameStrobe[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 493.360 0.000 493.920 0.560 ;
    END
  END FrameStrobe[43]
  PIN FrameStrobe[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 506.800 0.000 507.360 0.560 ;
    END
  END FrameStrobe[44]
  PIN FrameStrobe[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 520.240 0.000 520.800 0.560 ;
    END
  END FrameStrobe[45]
  PIN FrameStrobe[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 533.680 0.000 534.240 0.560 ;
    END
  END FrameStrobe[46]
  PIN FrameStrobe[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 547.120 0.000 547.680 0.560 ;
    END
  END FrameStrobe[47]
  PIN FrameStrobe[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 560.560 0.000 561.120 0.560 ;
    END
  END FrameStrobe[48]
  PIN FrameStrobe[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 574.000 0.000 574.560 0.560 ;
    END
  END FrameStrobe[49]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.412000 ;
    PORT
      LAYER Metal2 ;
        RECT 37.520 0.000 38.080 0.560 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 587.440 0.000 588.000 0.560 ;
    END
  END FrameStrobe[50]
  PIN FrameStrobe[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 600.880 0.000 601.440 0.560 ;
    END
  END FrameStrobe[51]
  PIN FrameStrobe[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 614.320 0.000 614.880 0.560 ;
    END
  END FrameStrobe[52]
  PIN FrameStrobe[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 627.760 0.000 628.320 0.560 ;
    END
  END FrameStrobe[53]
  PIN FrameStrobe[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 641.200 0.000 641.760 0.560 ;
    END
  END FrameStrobe[54]
  PIN FrameStrobe[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 654.640 0.000 655.200 0.560 ;
    END
  END FrameStrobe[55]
  PIN FrameStrobe[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 668.080 0.000 668.640 0.560 ;
    END
  END FrameStrobe[56]
  PIN FrameStrobe[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 681.520 0.000 682.080 0.560 ;
    END
  END FrameStrobe[57]
  PIN FrameStrobe[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 694.960 0.000 695.520 0.560 ;
    END
  END FrameStrobe[58]
  PIN FrameStrobe[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 708.400 0.000 708.960 0.560 ;
    END
  END FrameStrobe[59]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 44.240 0.000 44.800 0.560 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 740.320 0.000 740.880 0.560 ;
    END
  END FrameStrobe[60]
  PIN FrameStrobe[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 753.760 0.000 754.320 0.560 ;
    END
  END FrameStrobe[61]
  PIN FrameStrobe[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 767.200 0.000 767.760 0.560 ;
    END
  END FrameStrobe[62]
  PIN FrameStrobe[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 780.640 0.000 781.200 0.560 ;
    END
  END FrameStrobe[63]
  PIN FrameStrobe[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 794.080 0.000 794.640 0.560 ;
    END
  END FrameStrobe[64]
  PIN FrameStrobe[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 807.520 0.000 808.080 0.560 ;
    END
  END FrameStrobe[65]
  PIN FrameStrobe[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 820.960 0.000 821.520 0.560 ;
    END
  END FrameStrobe[66]
  PIN FrameStrobe[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 834.400 0.000 834.960 0.560 ;
    END
  END FrameStrobe[67]
  PIN FrameStrobe[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 847.840 0.000 848.400 0.560 ;
    END
  END FrameStrobe[68]
  PIN FrameStrobe[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 861.280 0.000 861.840 0.560 ;
    END
  END FrameStrobe[69]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 50.960 0.000 51.520 0.560 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 874.720 0.000 875.280 0.560 ;
    END
  END FrameStrobe[70]
  PIN FrameStrobe[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 888.160 0.000 888.720 0.560 ;
    END
  END FrameStrobe[71]
  PIN FrameStrobe[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 901.600 0.000 902.160 0.560 ;
    END
  END FrameStrobe[72]
  PIN FrameStrobe[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 915.040 0.000 915.600 0.560 ;
    END
  END FrameStrobe[73]
  PIN FrameStrobe[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 928.480 0.000 929.040 0.560 ;
    END
  END FrameStrobe[74]
  PIN FrameStrobe[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 941.920 0.000 942.480 0.560 ;
    END
  END FrameStrobe[75]
  PIN FrameStrobe[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 955.360 0.000 955.920 0.560 ;
    END
  END FrameStrobe[76]
  PIN FrameStrobe[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 968.800 0.000 969.360 0.560 ;
    END
  END FrameStrobe[77]
  PIN FrameStrobe[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 982.240 0.000 982.800 0.560 ;
    END
  END FrameStrobe[78]
  PIN FrameStrobe[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 995.680 0.000 996.240 0.560 ;
    END
  END FrameStrobe[79]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 57.680 0.000 58.240 0.560 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1034.320 0.000 1034.880 0.560 ;
    END
  END FrameStrobe[80]
  PIN FrameStrobe[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1048.880 0.000 1049.440 0.560 ;
    END
  END FrameStrobe[81]
  PIN FrameStrobe[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1063.440 0.000 1064.000 0.560 ;
    END
  END FrameStrobe[82]
  PIN FrameStrobe[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1078.000 0.000 1078.560 0.560 ;
    END
  END FrameStrobe[83]
  PIN FrameStrobe[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1092.560 0.000 1093.120 0.560 ;
    END
  END FrameStrobe[84]
  PIN FrameStrobe[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1107.120 0.000 1107.680 0.560 ;
    END
  END FrameStrobe[85]
  PIN FrameStrobe[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1121.680 0.000 1122.240 0.560 ;
    END
  END FrameStrobe[86]
  PIN FrameStrobe[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1136.240 0.000 1136.800 0.560 ;
    END
  END FrameStrobe[87]
  PIN FrameStrobe[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1150.800 0.000 1151.360 0.560 ;
    END
  END FrameStrobe[88]
  PIN FrameStrobe[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1165.360 0.000 1165.920 0.560 ;
    END
  END FrameStrobe[89]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 64.400 0.000 64.960 0.560 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1179.920 0.000 1180.480 0.560 ;
    END
  END FrameStrobe[90]
  PIN FrameStrobe[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1194.480 0.000 1195.040 0.560 ;
    END
  END FrameStrobe[91]
  PIN FrameStrobe[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1209.040 0.000 1209.600 0.560 ;
    END
  END FrameStrobe[92]
  PIN FrameStrobe[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1223.600 0.000 1224.160 0.560 ;
    END
  END FrameStrobe[93]
  PIN FrameStrobe[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1238.160 0.000 1238.720 0.560 ;
    END
  END FrameStrobe[94]
  PIN FrameStrobe[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1252.720 0.000 1253.280 0.560 ;
    END
  END FrameStrobe[95]
  PIN FrameStrobe[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1267.280 0.000 1267.840 0.560 ;
    END
  END FrameStrobe[96]
  PIN FrameStrobe[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1281.840 0.000 1282.400 0.560 ;
    END
  END FrameStrobe[97]
  PIN FrameStrobe[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1296.400 0.000 1296.960 0.560 ;
    END
  END FrameStrobe[98]
  PIN FrameStrobe[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1310.960 0.000 1311.520 0.560 ;
    END
  END FrameStrobe[99]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 71.120 0.000 71.680 0.560 ;
    END
  END FrameStrobe[9]
  PIN Tile_X0Y10_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 666.960 1.120 667.520 ;
    END
  END Tile_X0Y10_A_I_top
  PIN Tile_X0Y10_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 662.480 1.120 663.040 ;
    END
  END Tile_X0Y10_A_O_top
  PIN Tile_X0Y10_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 671.440 1.120 672.000 ;
    END
  END Tile_X0Y10_A_T_top
  PIN Tile_X0Y10_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 716.240 1.120 716.800 ;
    END
  END Tile_X0Y10_A_config_C_bit0
  PIN Tile_X0Y10_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 720.720 1.120 721.280 ;
    END
  END Tile_X0Y10_A_config_C_bit1
  PIN Tile_X0Y10_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 725.200 1.120 725.760 ;
    END
  END Tile_X0Y10_A_config_C_bit2
  PIN Tile_X0Y10_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 729.680 1.120 730.240 ;
    END
  END Tile_X0Y10_A_config_C_bit3
  PIN Tile_X0Y10_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 680.400 1.120 680.960 ;
    END
  END Tile_X0Y10_B_I_top
  PIN Tile_X0Y10_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 675.920 1.120 676.480 ;
    END
  END Tile_X0Y10_B_O_top
  PIN Tile_X0Y10_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 684.880 1.120 685.440 ;
    END
  END Tile_X0Y10_B_T_top
  PIN Tile_X0Y10_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 734.160 1.120 734.720 ;
    END
  END Tile_X0Y10_B_config_C_bit0
  PIN Tile_X0Y10_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 738.640 1.120 739.200 ;
    END
  END Tile_X0Y10_B_config_C_bit1
  PIN Tile_X0Y10_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 743.120 1.120 743.680 ;
    END
  END Tile_X0Y10_B_config_C_bit2
  PIN Tile_X0Y10_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 747.600 1.120 748.160 ;
    END
  END Tile_X0Y10_B_config_C_bit3
  PIN Tile_X0Y10_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 693.840 1.120 694.400 ;
    END
  END Tile_X0Y10_C_I_top
  PIN Tile_X0Y10_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 689.360 1.120 689.920 ;
    END
  END Tile_X0Y10_C_O_top
  PIN Tile_X0Y10_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 698.320 1.120 698.880 ;
    END
  END Tile_X0Y10_C_T_top
  PIN Tile_X0Y10_C_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 752.080 1.120 752.640 ;
    END
  END Tile_X0Y10_C_config_C_bit0
  PIN Tile_X0Y10_C_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 756.560 1.120 757.120 ;
    END
  END Tile_X0Y10_C_config_C_bit1
  PIN Tile_X0Y10_C_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 761.040 1.120 761.600 ;
    END
  END Tile_X0Y10_C_config_C_bit2
  PIN Tile_X0Y10_C_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 765.520 1.120 766.080 ;
    END
  END Tile_X0Y10_C_config_C_bit3
  PIN Tile_X0Y10_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 707.280 1.120 707.840 ;
    END
  END Tile_X0Y10_D_I_top
  PIN Tile_X0Y10_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 702.800 1.120 703.360 ;
    END
  END Tile_X0Y10_D_O_top
  PIN Tile_X0Y10_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 711.760 1.120 712.320 ;
    END
  END Tile_X0Y10_D_T_top
  PIN Tile_X0Y10_D_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 770.000 1.120 770.560 ;
    END
  END Tile_X0Y10_D_config_C_bit0
  PIN Tile_X0Y10_D_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 774.480 1.120 775.040 ;
    END
  END Tile_X0Y10_D_config_C_bit1
  PIN Tile_X0Y10_D_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 778.960 1.120 779.520 ;
    END
  END Tile_X0Y10_D_config_C_bit2
  PIN Tile_X0Y10_D_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 783.440 1.120 784.000 ;
    END
  END Tile_X0Y10_D_config_C_bit3
  PIN Tile_X0Y11_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 379.680 1.120 380.240 ;
    END
  END Tile_X0Y11_A_I_top
  PIN Tile_X0Y11_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 375.200 1.120 375.760 ;
    END
  END Tile_X0Y11_A_O_top
  PIN Tile_X0Y11_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 384.160 1.120 384.720 ;
    END
  END Tile_X0Y11_A_T_top
  PIN Tile_X0Y11_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 428.960 1.120 429.520 ;
    END
  END Tile_X0Y11_A_config_C_bit0
  PIN Tile_X0Y11_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 433.440 1.120 434.000 ;
    END
  END Tile_X0Y11_A_config_C_bit1
  PIN Tile_X0Y11_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 437.920 1.120 438.480 ;
    END
  END Tile_X0Y11_A_config_C_bit2
  PIN Tile_X0Y11_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 442.400 1.120 442.960 ;
    END
  END Tile_X0Y11_A_config_C_bit3
  PIN Tile_X0Y11_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 393.120 1.120 393.680 ;
    END
  END Tile_X0Y11_B_I_top
  PIN Tile_X0Y11_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 388.640 1.120 389.200 ;
    END
  END Tile_X0Y11_B_O_top
  PIN Tile_X0Y11_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 397.600 1.120 398.160 ;
    END
  END Tile_X0Y11_B_T_top
  PIN Tile_X0Y11_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 446.880 1.120 447.440 ;
    END
  END Tile_X0Y11_B_config_C_bit0
  PIN Tile_X0Y11_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 451.360 1.120 451.920 ;
    END
  END Tile_X0Y11_B_config_C_bit1
  PIN Tile_X0Y11_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 455.840 1.120 456.400 ;
    END
  END Tile_X0Y11_B_config_C_bit2
  PIN Tile_X0Y11_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 460.320 1.120 460.880 ;
    END
  END Tile_X0Y11_B_config_C_bit3
  PIN Tile_X0Y11_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 406.560 1.120 407.120 ;
    END
  END Tile_X0Y11_C_I_top
  PIN Tile_X0Y11_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 402.080 1.120 402.640 ;
    END
  END Tile_X0Y11_C_O_top
  PIN Tile_X0Y11_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 411.040 1.120 411.600 ;
    END
  END Tile_X0Y11_C_T_top
  PIN Tile_X0Y11_C_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 464.800 1.120 465.360 ;
    END
  END Tile_X0Y11_C_config_C_bit0
  PIN Tile_X0Y11_C_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 469.280 1.120 469.840 ;
    END
  END Tile_X0Y11_C_config_C_bit1
  PIN Tile_X0Y11_C_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 473.760 1.120 474.320 ;
    END
  END Tile_X0Y11_C_config_C_bit2
  PIN Tile_X0Y11_C_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 478.240 1.120 478.800 ;
    END
  END Tile_X0Y11_C_config_C_bit3
  PIN Tile_X0Y11_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 420.000 1.120 420.560 ;
    END
  END Tile_X0Y11_D_I_top
  PIN Tile_X0Y11_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 415.520 1.120 416.080 ;
    END
  END Tile_X0Y11_D_O_top
  PIN Tile_X0Y11_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 424.480 1.120 425.040 ;
    END
  END Tile_X0Y11_D_T_top
  PIN Tile_X0Y11_D_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 482.720 1.120 483.280 ;
    END
  END Tile_X0Y11_D_config_C_bit0
  PIN Tile_X0Y11_D_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 487.200 1.120 487.760 ;
    END
  END Tile_X0Y11_D_config_C_bit1
  PIN Tile_X0Y11_D_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 491.680 1.120 492.240 ;
    END
  END Tile_X0Y11_D_config_C_bit2
  PIN Tile_X0Y11_D_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 496.160 1.120 496.720 ;
    END
  END Tile_X0Y11_D_config_C_bit3
  PIN Tile_X0Y12_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 92.400 1.120 92.960 ;
    END
  END Tile_X0Y12_A_I_top
  PIN Tile_X0Y12_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.920 1.120 88.480 ;
    END
  END Tile_X0Y12_A_O_top
  PIN Tile_X0Y12_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.880 1.120 97.440 ;
    END
  END Tile_X0Y12_A_T_top
  PIN Tile_X0Y12_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.680 1.120 142.240 ;
    END
  END Tile_X0Y12_A_config_C_bit0
  PIN Tile_X0Y12_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 146.160 1.120 146.720 ;
    END
  END Tile_X0Y12_A_config_C_bit1
  PIN Tile_X0Y12_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.640 1.120 151.200 ;
    END
  END Tile_X0Y12_A_config_C_bit2
  PIN Tile_X0Y12_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 155.120 1.120 155.680 ;
    END
  END Tile_X0Y12_A_config_C_bit3
  PIN Tile_X0Y12_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 105.840 1.120 106.400 ;
    END
  END Tile_X0Y12_B_I_top
  PIN Tile_X0Y12_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 101.360 1.120 101.920 ;
    END
  END Tile_X0Y12_B_O_top
  PIN Tile_X0Y12_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.320 1.120 110.880 ;
    END
  END Tile_X0Y12_B_T_top
  PIN Tile_X0Y12_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 159.600 1.120 160.160 ;
    END
  END Tile_X0Y12_B_config_C_bit0
  PIN Tile_X0Y12_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.080 1.120 164.640 ;
    END
  END Tile_X0Y12_B_config_C_bit1
  PIN Tile_X0Y12_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.560 1.120 169.120 ;
    END
  END Tile_X0Y12_B_config_C_bit2
  PIN Tile_X0Y12_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 173.040 1.120 173.600 ;
    END
  END Tile_X0Y12_B_config_C_bit3
  PIN Tile_X0Y12_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 119.280 1.120 119.840 ;
    END
  END Tile_X0Y12_C_I_top
  PIN Tile_X0Y12_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.800 1.120 115.360 ;
    END
  END Tile_X0Y12_C_O_top
  PIN Tile_X0Y12_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 123.760 1.120 124.320 ;
    END
  END Tile_X0Y12_C_T_top
  PIN Tile_X0Y12_C_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 177.520 1.120 178.080 ;
    END
  END Tile_X0Y12_C_config_C_bit0
  PIN Tile_X0Y12_C_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.000 1.120 182.560 ;
    END
  END Tile_X0Y12_C_config_C_bit1
  PIN Tile_X0Y12_C_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 186.480 1.120 187.040 ;
    END
  END Tile_X0Y12_C_config_C_bit2
  PIN Tile_X0Y12_C_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 190.960 1.120 191.520 ;
    END
  END Tile_X0Y12_C_config_C_bit3
  PIN Tile_X0Y12_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.720 1.120 133.280 ;
    END
  END Tile_X0Y12_D_I_top
  PIN Tile_X0Y12_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 128.240 1.120 128.800 ;
    END
  END Tile_X0Y12_D_O_top
  PIN Tile_X0Y12_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.200 1.120 137.760 ;
    END
  END Tile_X0Y12_D_T_top
  PIN Tile_X0Y12_D_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 195.440 1.120 196.000 ;
    END
  END Tile_X0Y12_D_config_C_bit0
  PIN Tile_X0Y12_D_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 199.920 1.120 200.480 ;
    END
  END Tile_X0Y12_D_config_C_bit1
  PIN Tile_X0Y12_D_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.400 1.120 204.960 ;
    END
  END Tile_X0Y12_D_config_C_bit2
  PIN Tile_X0Y12_D_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 208.880 1.120 209.440 ;
    END
  END Tile_X0Y12_D_config_C_bit3
  PIN Tile_X0Y1_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3252.480 1.120 3253.040 ;
    END
  END Tile_X0Y1_A_I_top
  PIN Tile_X0Y1_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3248.000 1.120 3248.560 ;
    END
  END Tile_X0Y1_A_O_top
  PIN Tile_X0Y1_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3256.960 1.120 3257.520 ;
    END
  END Tile_X0Y1_A_T_top
  PIN Tile_X0Y1_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3301.760 1.120 3302.320 ;
    END
  END Tile_X0Y1_A_config_C_bit0
  PIN Tile_X0Y1_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3306.240 1.120 3306.800 ;
    END
  END Tile_X0Y1_A_config_C_bit1
  PIN Tile_X0Y1_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3310.720 1.120 3311.280 ;
    END
  END Tile_X0Y1_A_config_C_bit2
  PIN Tile_X0Y1_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3315.200 1.120 3315.760 ;
    END
  END Tile_X0Y1_A_config_C_bit3
  PIN Tile_X0Y1_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3265.920 1.120 3266.480 ;
    END
  END Tile_X0Y1_B_I_top
  PIN Tile_X0Y1_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3261.440 1.120 3262.000 ;
    END
  END Tile_X0Y1_B_O_top
  PIN Tile_X0Y1_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3270.400 1.120 3270.960 ;
    END
  END Tile_X0Y1_B_T_top
  PIN Tile_X0Y1_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3319.680 1.120 3320.240 ;
    END
  END Tile_X0Y1_B_config_C_bit0
  PIN Tile_X0Y1_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3324.160 1.120 3324.720 ;
    END
  END Tile_X0Y1_B_config_C_bit1
  PIN Tile_X0Y1_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3328.640 1.120 3329.200 ;
    END
  END Tile_X0Y1_B_config_C_bit2
  PIN Tile_X0Y1_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3333.120 1.120 3333.680 ;
    END
  END Tile_X0Y1_B_config_C_bit3
  PIN Tile_X0Y1_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3279.360 1.120 3279.920 ;
    END
  END Tile_X0Y1_C_I_top
  PIN Tile_X0Y1_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3274.880 1.120 3275.440 ;
    END
  END Tile_X0Y1_C_O_top
  PIN Tile_X0Y1_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3283.840 1.120 3284.400 ;
    END
  END Tile_X0Y1_C_T_top
  PIN Tile_X0Y1_C_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3337.600 1.120 3338.160 ;
    END
  END Tile_X0Y1_C_config_C_bit0
  PIN Tile_X0Y1_C_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3342.080 1.120 3342.640 ;
    END
  END Tile_X0Y1_C_config_C_bit1
  PIN Tile_X0Y1_C_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3346.560 1.120 3347.120 ;
    END
  END Tile_X0Y1_C_config_C_bit2
  PIN Tile_X0Y1_C_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3351.040 1.120 3351.600 ;
    END
  END Tile_X0Y1_C_config_C_bit3
  PIN Tile_X0Y1_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3292.800 1.120 3293.360 ;
    END
  END Tile_X0Y1_D_I_top
  PIN Tile_X0Y1_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3288.320 1.120 3288.880 ;
    END
  END Tile_X0Y1_D_O_top
  PIN Tile_X0Y1_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3297.280 1.120 3297.840 ;
    END
  END Tile_X0Y1_D_T_top
  PIN Tile_X0Y1_D_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3355.520 1.120 3356.080 ;
    END
  END Tile_X0Y1_D_config_C_bit0
  PIN Tile_X0Y1_D_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3360.000 1.120 3360.560 ;
    END
  END Tile_X0Y1_D_config_C_bit1
  PIN Tile_X0Y1_D_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3364.480 1.120 3365.040 ;
    END
  END Tile_X0Y1_D_config_C_bit2
  PIN Tile_X0Y1_D_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3368.960 1.120 3369.520 ;
    END
  END Tile_X0Y1_D_config_C_bit3
  PIN Tile_X0Y2_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2965.200 1.120 2965.760 ;
    END
  END Tile_X0Y2_A_I_top
  PIN Tile_X0Y2_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2960.720 1.120 2961.280 ;
    END
  END Tile_X0Y2_A_O_top
  PIN Tile_X0Y2_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2969.680 1.120 2970.240 ;
    END
  END Tile_X0Y2_A_T_top
  PIN Tile_X0Y2_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3014.480 1.120 3015.040 ;
    END
  END Tile_X0Y2_A_config_C_bit0
  PIN Tile_X0Y2_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3018.960 1.120 3019.520 ;
    END
  END Tile_X0Y2_A_config_C_bit1
  PIN Tile_X0Y2_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3023.440 1.120 3024.000 ;
    END
  END Tile_X0Y2_A_config_C_bit2
  PIN Tile_X0Y2_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3027.920 1.120 3028.480 ;
    END
  END Tile_X0Y2_A_config_C_bit3
  PIN Tile_X0Y2_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2978.640 1.120 2979.200 ;
    END
  END Tile_X0Y2_B_I_top
  PIN Tile_X0Y2_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2974.160 1.120 2974.720 ;
    END
  END Tile_X0Y2_B_O_top
  PIN Tile_X0Y2_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2983.120 1.120 2983.680 ;
    END
  END Tile_X0Y2_B_T_top
  PIN Tile_X0Y2_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3032.400 1.120 3032.960 ;
    END
  END Tile_X0Y2_B_config_C_bit0
  PIN Tile_X0Y2_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3036.880 1.120 3037.440 ;
    END
  END Tile_X0Y2_B_config_C_bit1
  PIN Tile_X0Y2_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3041.360 1.120 3041.920 ;
    END
  END Tile_X0Y2_B_config_C_bit2
  PIN Tile_X0Y2_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3045.840 1.120 3046.400 ;
    END
  END Tile_X0Y2_B_config_C_bit3
  PIN Tile_X0Y2_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2992.080 1.120 2992.640 ;
    END
  END Tile_X0Y2_C_I_top
  PIN Tile_X0Y2_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2987.600 1.120 2988.160 ;
    END
  END Tile_X0Y2_C_O_top
  PIN Tile_X0Y2_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2996.560 1.120 2997.120 ;
    END
  END Tile_X0Y2_C_T_top
  PIN Tile_X0Y2_C_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3050.320 1.120 3050.880 ;
    END
  END Tile_X0Y2_C_config_C_bit0
  PIN Tile_X0Y2_C_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3054.800 1.120 3055.360 ;
    END
  END Tile_X0Y2_C_config_C_bit1
  PIN Tile_X0Y2_C_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3059.280 1.120 3059.840 ;
    END
  END Tile_X0Y2_C_config_C_bit2
  PIN Tile_X0Y2_C_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3063.760 1.120 3064.320 ;
    END
  END Tile_X0Y2_C_config_C_bit3
  PIN Tile_X0Y2_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3005.520 1.120 3006.080 ;
    END
  END Tile_X0Y2_D_I_top
  PIN Tile_X0Y2_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3001.040 1.120 3001.600 ;
    END
  END Tile_X0Y2_D_O_top
  PIN Tile_X0Y2_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3010.000 1.120 3010.560 ;
    END
  END Tile_X0Y2_D_T_top
  PIN Tile_X0Y2_D_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3068.240 1.120 3068.800 ;
    END
  END Tile_X0Y2_D_config_C_bit0
  PIN Tile_X0Y2_D_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3072.720 1.120 3073.280 ;
    END
  END Tile_X0Y2_D_config_C_bit1
  PIN Tile_X0Y2_D_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3077.200 1.120 3077.760 ;
    END
  END Tile_X0Y2_D_config_C_bit2
  PIN Tile_X0Y2_D_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3081.680 1.120 3082.240 ;
    END
  END Tile_X0Y2_D_config_C_bit3
  PIN Tile_X0Y3_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2677.920 1.120 2678.480 ;
    END
  END Tile_X0Y3_A_I_top
  PIN Tile_X0Y3_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2673.440 1.120 2674.000 ;
    END
  END Tile_X0Y3_A_O_top
  PIN Tile_X0Y3_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2682.400 1.120 2682.960 ;
    END
  END Tile_X0Y3_A_T_top
  PIN Tile_X0Y3_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2727.200 1.120 2727.760 ;
    END
  END Tile_X0Y3_A_config_C_bit0
  PIN Tile_X0Y3_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2731.680 1.120 2732.240 ;
    END
  END Tile_X0Y3_A_config_C_bit1
  PIN Tile_X0Y3_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2736.160 1.120 2736.720 ;
    END
  END Tile_X0Y3_A_config_C_bit2
  PIN Tile_X0Y3_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2740.640 1.120 2741.200 ;
    END
  END Tile_X0Y3_A_config_C_bit3
  PIN Tile_X0Y3_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2691.360 1.120 2691.920 ;
    END
  END Tile_X0Y3_B_I_top
  PIN Tile_X0Y3_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2686.880 1.120 2687.440 ;
    END
  END Tile_X0Y3_B_O_top
  PIN Tile_X0Y3_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2695.840 1.120 2696.400 ;
    END
  END Tile_X0Y3_B_T_top
  PIN Tile_X0Y3_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2745.120 1.120 2745.680 ;
    END
  END Tile_X0Y3_B_config_C_bit0
  PIN Tile_X0Y3_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2749.600 1.120 2750.160 ;
    END
  END Tile_X0Y3_B_config_C_bit1
  PIN Tile_X0Y3_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2754.080 1.120 2754.640 ;
    END
  END Tile_X0Y3_B_config_C_bit2
  PIN Tile_X0Y3_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2758.560 1.120 2759.120 ;
    END
  END Tile_X0Y3_B_config_C_bit3
  PIN Tile_X0Y3_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2704.800 1.120 2705.360 ;
    END
  END Tile_X0Y3_C_I_top
  PIN Tile_X0Y3_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2700.320 1.120 2700.880 ;
    END
  END Tile_X0Y3_C_O_top
  PIN Tile_X0Y3_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2709.280 1.120 2709.840 ;
    END
  END Tile_X0Y3_C_T_top
  PIN Tile_X0Y3_C_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2763.040 1.120 2763.600 ;
    END
  END Tile_X0Y3_C_config_C_bit0
  PIN Tile_X0Y3_C_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2767.520 1.120 2768.080 ;
    END
  END Tile_X0Y3_C_config_C_bit1
  PIN Tile_X0Y3_C_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2772.000 1.120 2772.560 ;
    END
  END Tile_X0Y3_C_config_C_bit2
  PIN Tile_X0Y3_C_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2776.480 1.120 2777.040 ;
    END
  END Tile_X0Y3_C_config_C_bit3
  PIN Tile_X0Y3_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2718.240 1.120 2718.800 ;
    END
  END Tile_X0Y3_D_I_top
  PIN Tile_X0Y3_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2713.760 1.120 2714.320 ;
    END
  END Tile_X0Y3_D_O_top
  PIN Tile_X0Y3_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2722.720 1.120 2723.280 ;
    END
  END Tile_X0Y3_D_T_top
  PIN Tile_X0Y3_D_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2780.960 1.120 2781.520 ;
    END
  END Tile_X0Y3_D_config_C_bit0
  PIN Tile_X0Y3_D_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2785.440 1.120 2786.000 ;
    END
  END Tile_X0Y3_D_config_C_bit1
  PIN Tile_X0Y3_D_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2789.920 1.120 2790.480 ;
    END
  END Tile_X0Y3_D_config_C_bit2
  PIN Tile_X0Y3_D_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2794.400 1.120 2794.960 ;
    END
  END Tile_X0Y3_D_config_C_bit3
  PIN Tile_X0Y4_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2390.640 1.120 2391.200 ;
    END
  END Tile_X0Y4_A_I_top
  PIN Tile_X0Y4_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2386.160 1.120 2386.720 ;
    END
  END Tile_X0Y4_A_O_top
  PIN Tile_X0Y4_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2395.120 1.120 2395.680 ;
    END
  END Tile_X0Y4_A_T_top
  PIN Tile_X0Y4_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2439.920 1.120 2440.480 ;
    END
  END Tile_X0Y4_A_config_C_bit0
  PIN Tile_X0Y4_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2444.400 1.120 2444.960 ;
    END
  END Tile_X0Y4_A_config_C_bit1
  PIN Tile_X0Y4_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2448.880 1.120 2449.440 ;
    END
  END Tile_X0Y4_A_config_C_bit2
  PIN Tile_X0Y4_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2453.360 1.120 2453.920 ;
    END
  END Tile_X0Y4_A_config_C_bit3
  PIN Tile_X0Y4_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2404.080 1.120 2404.640 ;
    END
  END Tile_X0Y4_B_I_top
  PIN Tile_X0Y4_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2399.600 1.120 2400.160 ;
    END
  END Tile_X0Y4_B_O_top
  PIN Tile_X0Y4_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2408.560 1.120 2409.120 ;
    END
  END Tile_X0Y4_B_T_top
  PIN Tile_X0Y4_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2457.840 1.120 2458.400 ;
    END
  END Tile_X0Y4_B_config_C_bit0
  PIN Tile_X0Y4_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2462.320 1.120 2462.880 ;
    END
  END Tile_X0Y4_B_config_C_bit1
  PIN Tile_X0Y4_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2466.800 1.120 2467.360 ;
    END
  END Tile_X0Y4_B_config_C_bit2
  PIN Tile_X0Y4_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2471.280 1.120 2471.840 ;
    END
  END Tile_X0Y4_B_config_C_bit3
  PIN Tile_X0Y4_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2417.520 1.120 2418.080 ;
    END
  END Tile_X0Y4_C_I_top
  PIN Tile_X0Y4_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2413.040 1.120 2413.600 ;
    END
  END Tile_X0Y4_C_O_top
  PIN Tile_X0Y4_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2422.000 1.120 2422.560 ;
    END
  END Tile_X0Y4_C_T_top
  PIN Tile_X0Y4_C_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2475.760 1.120 2476.320 ;
    END
  END Tile_X0Y4_C_config_C_bit0
  PIN Tile_X0Y4_C_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2480.240 1.120 2480.800 ;
    END
  END Tile_X0Y4_C_config_C_bit1
  PIN Tile_X0Y4_C_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2484.720 1.120 2485.280 ;
    END
  END Tile_X0Y4_C_config_C_bit2
  PIN Tile_X0Y4_C_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2489.200 1.120 2489.760 ;
    END
  END Tile_X0Y4_C_config_C_bit3
  PIN Tile_X0Y4_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2430.960 1.120 2431.520 ;
    END
  END Tile_X0Y4_D_I_top
  PIN Tile_X0Y4_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2426.480 1.120 2427.040 ;
    END
  END Tile_X0Y4_D_O_top
  PIN Tile_X0Y4_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2435.440 1.120 2436.000 ;
    END
  END Tile_X0Y4_D_T_top
  PIN Tile_X0Y4_D_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2493.680 1.120 2494.240 ;
    END
  END Tile_X0Y4_D_config_C_bit0
  PIN Tile_X0Y4_D_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2498.160 1.120 2498.720 ;
    END
  END Tile_X0Y4_D_config_C_bit1
  PIN Tile_X0Y4_D_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2502.640 1.120 2503.200 ;
    END
  END Tile_X0Y4_D_config_C_bit2
  PIN Tile_X0Y4_D_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2507.120 1.120 2507.680 ;
    END
  END Tile_X0Y4_D_config_C_bit3
  PIN Tile_X0Y5_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2103.360 1.120 2103.920 ;
    END
  END Tile_X0Y5_A_I_top
  PIN Tile_X0Y5_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2098.880 1.120 2099.440 ;
    END
  END Tile_X0Y5_A_O_top
  PIN Tile_X0Y5_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2107.840 1.120 2108.400 ;
    END
  END Tile_X0Y5_A_T_top
  PIN Tile_X0Y5_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2152.640 1.120 2153.200 ;
    END
  END Tile_X0Y5_A_config_C_bit0
  PIN Tile_X0Y5_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2157.120 1.120 2157.680 ;
    END
  END Tile_X0Y5_A_config_C_bit1
  PIN Tile_X0Y5_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2161.600 1.120 2162.160 ;
    END
  END Tile_X0Y5_A_config_C_bit2
  PIN Tile_X0Y5_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2166.080 1.120 2166.640 ;
    END
  END Tile_X0Y5_A_config_C_bit3
  PIN Tile_X0Y5_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2116.800 1.120 2117.360 ;
    END
  END Tile_X0Y5_B_I_top
  PIN Tile_X0Y5_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2112.320 1.120 2112.880 ;
    END
  END Tile_X0Y5_B_O_top
  PIN Tile_X0Y5_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2121.280 1.120 2121.840 ;
    END
  END Tile_X0Y5_B_T_top
  PIN Tile_X0Y5_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2170.560 1.120 2171.120 ;
    END
  END Tile_X0Y5_B_config_C_bit0
  PIN Tile_X0Y5_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2175.040 1.120 2175.600 ;
    END
  END Tile_X0Y5_B_config_C_bit1
  PIN Tile_X0Y5_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2179.520 1.120 2180.080 ;
    END
  END Tile_X0Y5_B_config_C_bit2
  PIN Tile_X0Y5_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2184.000 1.120 2184.560 ;
    END
  END Tile_X0Y5_B_config_C_bit3
  PIN Tile_X0Y5_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2130.240 1.120 2130.800 ;
    END
  END Tile_X0Y5_C_I_top
  PIN Tile_X0Y5_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2125.760 1.120 2126.320 ;
    END
  END Tile_X0Y5_C_O_top
  PIN Tile_X0Y5_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2134.720 1.120 2135.280 ;
    END
  END Tile_X0Y5_C_T_top
  PIN Tile_X0Y5_C_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2188.480 1.120 2189.040 ;
    END
  END Tile_X0Y5_C_config_C_bit0
  PIN Tile_X0Y5_C_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2192.960 1.120 2193.520 ;
    END
  END Tile_X0Y5_C_config_C_bit1
  PIN Tile_X0Y5_C_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2197.440 1.120 2198.000 ;
    END
  END Tile_X0Y5_C_config_C_bit2
  PIN Tile_X0Y5_C_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2201.920 1.120 2202.480 ;
    END
  END Tile_X0Y5_C_config_C_bit3
  PIN Tile_X0Y5_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2143.680 1.120 2144.240 ;
    END
  END Tile_X0Y5_D_I_top
  PIN Tile_X0Y5_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2139.200 1.120 2139.760 ;
    END
  END Tile_X0Y5_D_O_top
  PIN Tile_X0Y5_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2148.160 1.120 2148.720 ;
    END
  END Tile_X0Y5_D_T_top
  PIN Tile_X0Y5_D_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2206.400 1.120 2206.960 ;
    END
  END Tile_X0Y5_D_config_C_bit0
  PIN Tile_X0Y5_D_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2210.880 1.120 2211.440 ;
    END
  END Tile_X0Y5_D_config_C_bit1
  PIN Tile_X0Y5_D_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2215.360 1.120 2215.920 ;
    END
  END Tile_X0Y5_D_config_C_bit2
  PIN Tile_X0Y5_D_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2219.840 1.120 2220.400 ;
    END
  END Tile_X0Y5_D_config_C_bit3
  PIN Tile_X0Y6_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1816.080 1.120 1816.640 ;
    END
  END Tile_X0Y6_A_I_top
  PIN Tile_X0Y6_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1811.600 1.120 1812.160 ;
    END
  END Tile_X0Y6_A_O_top
  PIN Tile_X0Y6_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1820.560 1.120 1821.120 ;
    END
  END Tile_X0Y6_A_T_top
  PIN Tile_X0Y6_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1865.360 1.120 1865.920 ;
    END
  END Tile_X0Y6_A_config_C_bit0
  PIN Tile_X0Y6_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1869.840 1.120 1870.400 ;
    END
  END Tile_X0Y6_A_config_C_bit1
  PIN Tile_X0Y6_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1874.320 1.120 1874.880 ;
    END
  END Tile_X0Y6_A_config_C_bit2
  PIN Tile_X0Y6_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1878.800 1.120 1879.360 ;
    END
  END Tile_X0Y6_A_config_C_bit3
  PIN Tile_X0Y6_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1829.520 1.120 1830.080 ;
    END
  END Tile_X0Y6_B_I_top
  PIN Tile_X0Y6_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1825.040 1.120 1825.600 ;
    END
  END Tile_X0Y6_B_O_top
  PIN Tile_X0Y6_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1834.000 1.120 1834.560 ;
    END
  END Tile_X0Y6_B_T_top
  PIN Tile_X0Y6_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1883.280 1.120 1883.840 ;
    END
  END Tile_X0Y6_B_config_C_bit0
  PIN Tile_X0Y6_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1887.760 1.120 1888.320 ;
    END
  END Tile_X0Y6_B_config_C_bit1
  PIN Tile_X0Y6_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1892.240 1.120 1892.800 ;
    END
  END Tile_X0Y6_B_config_C_bit2
  PIN Tile_X0Y6_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1896.720 1.120 1897.280 ;
    END
  END Tile_X0Y6_B_config_C_bit3
  PIN Tile_X0Y6_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1842.960 1.120 1843.520 ;
    END
  END Tile_X0Y6_C_I_top
  PIN Tile_X0Y6_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1838.480 1.120 1839.040 ;
    END
  END Tile_X0Y6_C_O_top
  PIN Tile_X0Y6_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1847.440 1.120 1848.000 ;
    END
  END Tile_X0Y6_C_T_top
  PIN Tile_X0Y6_C_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1901.200 1.120 1901.760 ;
    END
  END Tile_X0Y6_C_config_C_bit0
  PIN Tile_X0Y6_C_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1905.680 1.120 1906.240 ;
    END
  END Tile_X0Y6_C_config_C_bit1
  PIN Tile_X0Y6_C_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1910.160 1.120 1910.720 ;
    END
  END Tile_X0Y6_C_config_C_bit2
  PIN Tile_X0Y6_C_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1914.640 1.120 1915.200 ;
    END
  END Tile_X0Y6_C_config_C_bit3
  PIN Tile_X0Y6_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1856.400 1.120 1856.960 ;
    END
  END Tile_X0Y6_D_I_top
  PIN Tile_X0Y6_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1851.920 1.120 1852.480 ;
    END
  END Tile_X0Y6_D_O_top
  PIN Tile_X0Y6_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1860.880 1.120 1861.440 ;
    END
  END Tile_X0Y6_D_T_top
  PIN Tile_X0Y6_D_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1919.120 1.120 1919.680 ;
    END
  END Tile_X0Y6_D_config_C_bit0
  PIN Tile_X0Y6_D_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1923.600 1.120 1924.160 ;
    END
  END Tile_X0Y6_D_config_C_bit1
  PIN Tile_X0Y6_D_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1928.080 1.120 1928.640 ;
    END
  END Tile_X0Y6_D_config_C_bit2
  PIN Tile_X0Y6_D_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1932.560 1.120 1933.120 ;
    END
  END Tile_X0Y6_D_config_C_bit3
  PIN Tile_X0Y7_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1528.800 1.120 1529.360 ;
    END
  END Tile_X0Y7_A_I_top
  PIN Tile_X0Y7_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1524.320 1.120 1524.880 ;
    END
  END Tile_X0Y7_A_O_top
  PIN Tile_X0Y7_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1533.280 1.120 1533.840 ;
    END
  END Tile_X0Y7_A_T_top
  PIN Tile_X0Y7_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1578.080 1.120 1578.640 ;
    END
  END Tile_X0Y7_A_config_C_bit0
  PIN Tile_X0Y7_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1582.560 1.120 1583.120 ;
    END
  END Tile_X0Y7_A_config_C_bit1
  PIN Tile_X0Y7_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1587.040 1.120 1587.600 ;
    END
  END Tile_X0Y7_A_config_C_bit2
  PIN Tile_X0Y7_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1591.520 1.120 1592.080 ;
    END
  END Tile_X0Y7_A_config_C_bit3
  PIN Tile_X0Y7_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1542.240 1.120 1542.800 ;
    END
  END Tile_X0Y7_B_I_top
  PIN Tile_X0Y7_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1537.760 1.120 1538.320 ;
    END
  END Tile_X0Y7_B_O_top
  PIN Tile_X0Y7_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1546.720 1.120 1547.280 ;
    END
  END Tile_X0Y7_B_T_top
  PIN Tile_X0Y7_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1596.000 1.120 1596.560 ;
    END
  END Tile_X0Y7_B_config_C_bit0
  PIN Tile_X0Y7_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1600.480 1.120 1601.040 ;
    END
  END Tile_X0Y7_B_config_C_bit1
  PIN Tile_X0Y7_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1604.960 1.120 1605.520 ;
    END
  END Tile_X0Y7_B_config_C_bit2
  PIN Tile_X0Y7_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1609.440 1.120 1610.000 ;
    END
  END Tile_X0Y7_B_config_C_bit3
  PIN Tile_X0Y7_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1555.680 1.120 1556.240 ;
    END
  END Tile_X0Y7_C_I_top
  PIN Tile_X0Y7_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1551.200 1.120 1551.760 ;
    END
  END Tile_X0Y7_C_O_top
  PIN Tile_X0Y7_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1560.160 1.120 1560.720 ;
    END
  END Tile_X0Y7_C_T_top
  PIN Tile_X0Y7_C_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1613.920 1.120 1614.480 ;
    END
  END Tile_X0Y7_C_config_C_bit0
  PIN Tile_X0Y7_C_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1618.400 1.120 1618.960 ;
    END
  END Tile_X0Y7_C_config_C_bit1
  PIN Tile_X0Y7_C_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1622.880 1.120 1623.440 ;
    END
  END Tile_X0Y7_C_config_C_bit2
  PIN Tile_X0Y7_C_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1627.360 1.120 1627.920 ;
    END
  END Tile_X0Y7_C_config_C_bit3
  PIN Tile_X0Y7_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1569.120 1.120 1569.680 ;
    END
  END Tile_X0Y7_D_I_top
  PIN Tile_X0Y7_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1564.640 1.120 1565.200 ;
    END
  END Tile_X0Y7_D_O_top
  PIN Tile_X0Y7_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1573.600 1.120 1574.160 ;
    END
  END Tile_X0Y7_D_T_top
  PIN Tile_X0Y7_D_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1631.840 1.120 1632.400 ;
    END
  END Tile_X0Y7_D_config_C_bit0
  PIN Tile_X0Y7_D_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1636.320 1.120 1636.880 ;
    END
  END Tile_X0Y7_D_config_C_bit1
  PIN Tile_X0Y7_D_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1640.800 1.120 1641.360 ;
    END
  END Tile_X0Y7_D_config_C_bit2
  PIN Tile_X0Y7_D_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1645.280 1.120 1645.840 ;
    END
  END Tile_X0Y7_D_config_C_bit3
  PIN Tile_X0Y8_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1241.520 1.120 1242.080 ;
    END
  END Tile_X0Y8_A_I_top
  PIN Tile_X0Y8_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1237.040 1.120 1237.600 ;
    END
  END Tile_X0Y8_A_O_top
  PIN Tile_X0Y8_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1246.000 1.120 1246.560 ;
    END
  END Tile_X0Y8_A_T_top
  PIN Tile_X0Y8_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1290.800 1.120 1291.360 ;
    END
  END Tile_X0Y8_A_config_C_bit0
  PIN Tile_X0Y8_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1295.280 1.120 1295.840 ;
    END
  END Tile_X0Y8_A_config_C_bit1
  PIN Tile_X0Y8_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1299.760 1.120 1300.320 ;
    END
  END Tile_X0Y8_A_config_C_bit2
  PIN Tile_X0Y8_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1304.240 1.120 1304.800 ;
    END
  END Tile_X0Y8_A_config_C_bit3
  PIN Tile_X0Y8_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1254.960 1.120 1255.520 ;
    END
  END Tile_X0Y8_B_I_top
  PIN Tile_X0Y8_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1250.480 1.120 1251.040 ;
    END
  END Tile_X0Y8_B_O_top
  PIN Tile_X0Y8_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1259.440 1.120 1260.000 ;
    END
  END Tile_X0Y8_B_T_top
  PIN Tile_X0Y8_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1308.720 1.120 1309.280 ;
    END
  END Tile_X0Y8_B_config_C_bit0
  PIN Tile_X0Y8_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1313.200 1.120 1313.760 ;
    END
  END Tile_X0Y8_B_config_C_bit1
  PIN Tile_X0Y8_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1317.680 1.120 1318.240 ;
    END
  END Tile_X0Y8_B_config_C_bit2
  PIN Tile_X0Y8_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1322.160 1.120 1322.720 ;
    END
  END Tile_X0Y8_B_config_C_bit3
  PIN Tile_X0Y8_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1268.400 1.120 1268.960 ;
    END
  END Tile_X0Y8_C_I_top
  PIN Tile_X0Y8_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1263.920 1.120 1264.480 ;
    END
  END Tile_X0Y8_C_O_top
  PIN Tile_X0Y8_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1272.880 1.120 1273.440 ;
    END
  END Tile_X0Y8_C_T_top
  PIN Tile_X0Y8_C_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1326.640 1.120 1327.200 ;
    END
  END Tile_X0Y8_C_config_C_bit0
  PIN Tile_X0Y8_C_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1331.120 1.120 1331.680 ;
    END
  END Tile_X0Y8_C_config_C_bit1
  PIN Tile_X0Y8_C_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1335.600 1.120 1336.160 ;
    END
  END Tile_X0Y8_C_config_C_bit2
  PIN Tile_X0Y8_C_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1340.080 1.120 1340.640 ;
    END
  END Tile_X0Y8_C_config_C_bit3
  PIN Tile_X0Y8_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1281.840 1.120 1282.400 ;
    END
  END Tile_X0Y8_D_I_top
  PIN Tile_X0Y8_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1277.360 1.120 1277.920 ;
    END
  END Tile_X0Y8_D_O_top
  PIN Tile_X0Y8_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1286.320 1.120 1286.880 ;
    END
  END Tile_X0Y8_D_T_top
  PIN Tile_X0Y8_D_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1344.560 1.120 1345.120 ;
    END
  END Tile_X0Y8_D_config_C_bit0
  PIN Tile_X0Y8_D_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1349.040 1.120 1349.600 ;
    END
  END Tile_X0Y8_D_config_C_bit1
  PIN Tile_X0Y8_D_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1353.520 1.120 1354.080 ;
    END
  END Tile_X0Y8_D_config_C_bit2
  PIN Tile_X0Y8_D_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1358.000 1.120 1358.560 ;
    END
  END Tile_X0Y8_D_config_C_bit3
  PIN Tile_X0Y9_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 954.240 1.120 954.800 ;
    END
  END Tile_X0Y9_A_I_top
  PIN Tile_X0Y9_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 949.760 1.120 950.320 ;
    END
  END Tile_X0Y9_A_O_top
  PIN Tile_X0Y9_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 958.720 1.120 959.280 ;
    END
  END Tile_X0Y9_A_T_top
  PIN Tile_X0Y9_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1003.520 1.120 1004.080 ;
    END
  END Tile_X0Y9_A_config_C_bit0
  PIN Tile_X0Y9_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1008.000 1.120 1008.560 ;
    END
  END Tile_X0Y9_A_config_C_bit1
  PIN Tile_X0Y9_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1012.480 1.120 1013.040 ;
    END
  END Tile_X0Y9_A_config_C_bit2
  PIN Tile_X0Y9_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1016.960 1.120 1017.520 ;
    END
  END Tile_X0Y9_A_config_C_bit3
  PIN Tile_X0Y9_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 967.680 1.120 968.240 ;
    END
  END Tile_X0Y9_B_I_top
  PIN Tile_X0Y9_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 963.200 1.120 963.760 ;
    END
  END Tile_X0Y9_B_O_top
  PIN Tile_X0Y9_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 972.160 1.120 972.720 ;
    END
  END Tile_X0Y9_B_T_top
  PIN Tile_X0Y9_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1021.440 1.120 1022.000 ;
    END
  END Tile_X0Y9_B_config_C_bit0
  PIN Tile_X0Y9_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1025.920 1.120 1026.480 ;
    END
  END Tile_X0Y9_B_config_C_bit1
  PIN Tile_X0Y9_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1030.400 1.120 1030.960 ;
    END
  END Tile_X0Y9_B_config_C_bit2
  PIN Tile_X0Y9_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1034.880 1.120 1035.440 ;
    END
  END Tile_X0Y9_B_config_C_bit3
  PIN Tile_X0Y9_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 981.120 1.120 981.680 ;
    END
  END Tile_X0Y9_C_I_top
  PIN Tile_X0Y9_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 976.640 1.120 977.200 ;
    END
  END Tile_X0Y9_C_O_top
  PIN Tile_X0Y9_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 985.600 1.120 986.160 ;
    END
  END Tile_X0Y9_C_T_top
  PIN Tile_X0Y9_C_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1039.360 1.120 1039.920 ;
    END
  END Tile_X0Y9_C_config_C_bit0
  PIN Tile_X0Y9_C_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1043.840 1.120 1044.400 ;
    END
  END Tile_X0Y9_C_config_C_bit1
  PIN Tile_X0Y9_C_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1048.320 1.120 1048.880 ;
    END
  END Tile_X0Y9_C_config_C_bit2
  PIN Tile_X0Y9_C_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1052.800 1.120 1053.360 ;
    END
  END Tile_X0Y9_C_config_C_bit3
  PIN Tile_X0Y9_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 994.560 1.120 995.120 ;
    END
  END Tile_X0Y9_D_I_top
  PIN Tile_X0Y9_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.405000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 990.080 1.120 990.640 ;
    END
  END Tile_X0Y9_D_O_top
  PIN Tile_X0Y9_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 999.040 1.120 999.600 ;
    END
  END Tile_X0Y9_D_T_top
  PIN Tile_X0Y9_D_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1057.280 1.120 1057.840 ;
    END
  END Tile_X0Y9_D_config_C_bit0
  PIN Tile_X0Y9_D_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1061.760 1.120 1062.320 ;
    END
  END Tile_X0Y9_D_config_C_bit1
  PIN Tile_X0Y9_D_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1066.240 1.120 1066.800 ;
    END
  END Tile_X0Y9_D_config_C_bit2
  PIN Tile_X0Y9_D_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1070.720 1.120 1071.280 ;
    END
  END Tile_X0Y9_D_config_C_bit3
  PIN Tile_X1Y13_BOOT_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 210.560 0.000 211.120 0.560 ;
    END
  END Tile_X1Y13_BOOT_top
  PIN Tile_X1Y13_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 0.000 160.720 0.560 ;
    END
  END Tile_X1Y13_CONFIGURED_top
  PIN Tile_X1Y13_RESET_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 1.641600 ;
    PORT
      LAYER Metal2 ;
        RECT 150.080 0.000 150.640 0.560 ;
    END
  END Tile_X1Y13_RESET_top
  PIN Tile_X1Y13_SLOT_top0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 170.240 0.000 170.800 0.560 ;
    END
  END Tile_X1Y13_SLOT_top0
  PIN Tile_X1Y13_SLOT_top1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 0.000 180.880 0.560 ;
    END
  END Tile_X1Y13_SLOT_top1
  PIN Tile_X1Y13_SLOT_top2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 0.000 190.960 0.560 ;
    END
  END Tile_X1Y13_SLOT_top2
  PIN Tile_X1Y13_SLOT_top3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 200.480 0.000 201.040 0.560 ;
    END
  END Tile_X1Y13_SLOT_top3
  PIN Tile_X8Y10_A_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 750.960 2324.560 751.520 ;
    END
  END Tile_X8Y10_A_SRAM0
  PIN Tile_X8Y10_A_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 755.440 2324.560 756.000 ;
    END
  END Tile_X8Y10_A_SRAM1
  PIN Tile_X8Y10_A_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 759.920 2324.560 760.480 ;
    END
  END Tile_X8Y10_A_SRAM2
  PIN Tile_X8Y10_A_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 764.400 2324.560 764.960 ;
    END
  END Tile_X8Y10_A_SRAM3
  PIN Tile_X8Y10_A_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 768.880 2324.560 769.440 ;
    END
  END Tile_X8Y10_A_SRAM4
  PIN Tile_X8Y10_A_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 773.360 2324.560 773.920 ;
    END
  END Tile_X8Y10_A_SRAM5
  PIN Tile_X8Y10_A_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 777.840 2324.560 778.400 ;
    END
  END Tile_X8Y10_A_SRAM6
  PIN Tile_X8Y10_A_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 782.320 2324.560 782.880 ;
    END
  END Tile_X8Y10_A_SRAM7
  PIN Tile_X8Y10_A_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 786.800 2324.560 787.360 ;
    END
  END Tile_X8Y10_A_SRAM8
  PIN Tile_X8Y10_CEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 706.160 2324.560 706.720 ;
    END
  END Tile_X8Y10_CEN_SRAM
  PIN Tile_X8Y10_CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 827.120 2324.560 827.680 ;
    END
  END Tile_X8Y10_CLK_SRAM
  PIN Tile_X8Y10_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 701.680 2324.560 702.240 ;
    END
  END Tile_X8Y10_CONFIGURED_top
  PIN Tile_X8Y10_D_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 791.280 2324.560 791.840 ;
    END
  END Tile_X8Y10_D_SRAM0
  PIN Tile_X8Y10_D_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 795.760 2324.560 796.320 ;
    END
  END Tile_X8Y10_D_SRAM1
  PIN Tile_X8Y10_D_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 800.240 2324.560 800.800 ;
    END
  END Tile_X8Y10_D_SRAM2
  PIN Tile_X8Y10_D_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 804.720 2324.560 805.280 ;
    END
  END Tile_X8Y10_D_SRAM3
  PIN Tile_X8Y10_D_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 809.200 2324.560 809.760 ;
    END
  END Tile_X8Y10_D_SRAM4
  PIN Tile_X8Y10_D_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 813.680 2324.560 814.240 ;
    END
  END Tile_X8Y10_D_SRAM5
  PIN Tile_X8Y10_D_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 818.160 2324.560 818.720 ;
    END
  END Tile_X8Y10_D_SRAM6
  PIN Tile_X8Y10_D_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 822.640 2324.560 823.200 ;
    END
  END Tile_X8Y10_D_SRAM7
  PIN Tile_X8Y10_GWEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 710.640 2324.560 711.200 ;
    END
  END Tile_X8Y10_GWEN_SRAM
  PIN Tile_X8Y10_Q_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 665.840 2324.560 666.400 ;
    END
  END Tile_X8Y10_Q_SRAM0
  PIN Tile_X8Y10_Q_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 670.320 2324.560 670.880 ;
    END
  END Tile_X8Y10_Q_SRAM1
  PIN Tile_X8Y10_Q_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 674.800 2324.560 675.360 ;
    END
  END Tile_X8Y10_Q_SRAM2
  PIN Tile_X8Y10_Q_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 679.280 2324.560 679.840 ;
    END
  END Tile_X8Y10_Q_SRAM3
  PIN Tile_X8Y10_Q_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.531500 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 683.760 2324.560 684.320 ;
    END
  END Tile_X8Y10_Q_SRAM4
  PIN Tile_X8Y10_Q_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.528500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 688.240 2324.560 688.800 ;
    END
  END Tile_X8Y10_Q_SRAM5
  PIN Tile_X8Y10_Q_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 692.720 2324.560 693.280 ;
    END
  END Tile_X8Y10_Q_SRAM6
  PIN Tile_X8Y10_Q_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 697.200 2324.560 697.760 ;
    END
  END Tile_X8Y10_Q_SRAM7
  PIN Tile_X8Y10_WEN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 715.120 2324.560 715.680 ;
    END
  END Tile_X8Y10_WEN_SRAM0
  PIN Tile_X8Y10_WEN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 719.600 2324.560 720.160 ;
    END
  END Tile_X8Y10_WEN_SRAM1
  PIN Tile_X8Y10_WEN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 724.080 2324.560 724.640 ;
    END
  END Tile_X8Y10_WEN_SRAM2
  PIN Tile_X8Y10_WEN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 728.560 2324.560 729.120 ;
    END
  END Tile_X8Y10_WEN_SRAM3
  PIN Tile_X8Y10_WEN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 733.040 2324.560 733.600 ;
    END
  END Tile_X8Y10_WEN_SRAM4
  PIN Tile_X8Y10_WEN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 737.520 2324.560 738.080 ;
    END
  END Tile_X8Y10_WEN_SRAM5
  PIN Tile_X8Y10_WEN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 742.000 2324.560 742.560 ;
    END
  END Tile_X8Y10_WEN_SRAM6
  PIN Tile_X8Y10_WEN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 746.480 2324.560 747.040 ;
    END
  END Tile_X8Y10_WEN_SRAM7
  PIN Tile_X8Y12_A_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 176.400 2324.560 176.960 ;
    END
  END Tile_X8Y12_A_SRAM0
  PIN Tile_X8Y12_A_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 180.880 2324.560 181.440 ;
    END
  END Tile_X8Y12_A_SRAM1
  PIN Tile_X8Y12_A_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 185.360 2324.560 185.920 ;
    END
  END Tile_X8Y12_A_SRAM2
  PIN Tile_X8Y12_A_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 189.840 2324.560 190.400 ;
    END
  END Tile_X8Y12_A_SRAM3
  PIN Tile_X8Y12_A_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 194.320 2324.560 194.880 ;
    END
  END Tile_X8Y12_A_SRAM4
  PIN Tile_X8Y12_A_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 198.800 2324.560 199.360 ;
    END
  END Tile_X8Y12_A_SRAM5
  PIN Tile_X8Y12_A_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 203.280 2324.560 203.840 ;
    END
  END Tile_X8Y12_A_SRAM6
  PIN Tile_X8Y12_A_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 207.760 2324.560 208.320 ;
    END
  END Tile_X8Y12_A_SRAM7
  PIN Tile_X8Y12_A_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 212.240 2324.560 212.800 ;
    END
  END Tile_X8Y12_A_SRAM8
  PIN Tile_X8Y12_CEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 131.600 2324.560 132.160 ;
    END
  END Tile_X8Y12_CEN_SRAM
  PIN Tile_X8Y12_CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 252.560 2324.560 253.120 ;
    END
  END Tile_X8Y12_CLK_SRAM
  PIN Tile_X8Y12_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 127.120 2324.560 127.680 ;
    END
  END Tile_X8Y12_CONFIGURED_top
  PIN Tile_X8Y12_D_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 216.720 2324.560 217.280 ;
    END
  END Tile_X8Y12_D_SRAM0
  PIN Tile_X8Y12_D_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 221.200 2324.560 221.760 ;
    END
  END Tile_X8Y12_D_SRAM1
  PIN Tile_X8Y12_D_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 225.680 2324.560 226.240 ;
    END
  END Tile_X8Y12_D_SRAM2
  PIN Tile_X8Y12_D_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 230.160 2324.560 230.720 ;
    END
  END Tile_X8Y12_D_SRAM3
  PIN Tile_X8Y12_D_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 234.640 2324.560 235.200 ;
    END
  END Tile_X8Y12_D_SRAM4
  PIN Tile_X8Y12_D_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 239.120 2324.560 239.680 ;
    END
  END Tile_X8Y12_D_SRAM5
  PIN Tile_X8Y12_D_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 243.600 2324.560 244.160 ;
    END
  END Tile_X8Y12_D_SRAM6
  PIN Tile_X8Y12_D_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 248.080 2324.560 248.640 ;
    END
  END Tile_X8Y12_D_SRAM7
  PIN Tile_X8Y12_GWEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 136.080 2324.560 136.640 ;
    END
  END Tile_X8Y12_GWEN_SRAM
  PIN Tile_X8Y12_Q_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 91.280 2324.560 91.840 ;
    END
  END Tile_X8Y12_Q_SRAM0
  PIN Tile_X8Y12_Q_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 95.760 2324.560 96.320 ;
    END
  END Tile_X8Y12_Q_SRAM1
  PIN Tile_X8Y12_Q_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 100.240 2324.560 100.800 ;
    END
  END Tile_X8Y12_Q_SRAM2
  PIN Tile_X8Y12_Q_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 104.720 2324.560 105.280 ;
    END
  END Tile_X8Y12_Q_SRAM3
  PIN Tile_X8Y12_Q_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.531500 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 109.200 2324.560 109.760 ;
    END
  END Tile_X8Y12_Q_SRAM4
  PIN Tile_X8Y12_Q_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.528500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 113.680 2324.560 114.240 ;
    END
  END Tile_X8Y12_Q_SRAM5
  PIN Tile_X8Y12_Q_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 118.160 2324.560 118.720 ;
    END
  END Tile_X8Y12_Q_SRAM6
  PIN Tile_X8Y12_Q_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 122.640 2324.560 123.200 ;
    END
  END Tile_X8Y12_Q_SRAM7
  PIN Tile_X8Y12_WEN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 140.560 2324.560 141.120 ;
    END
  END Tile_X8Y12_WEN_SRAM0
  PIN Tile_X8Y12_WEN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 145.040 2324.560 145.600 ;
    END
  END Tile_X8Y12_WEN_SRAM1
  PIN Tile_X8Y12_WEN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 149.520 2324.560 150.080 ;
    END
  END Tile_X8Y12_WEN_SRAM2
  PIN Tile_X8Y12_WEN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 154.000 2324.560 154.560 ;
    END
  END Tile_X8Y12_WEN_SRAM3
  PIN Tile_X8Y12_WEN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 158.480 2324.560 159.040 ;
    END
  END Tile_X8Y12_WEN_SRAM4
  PIN Tile_X8Y12_WEN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 162.960 2324.560 163.520 ;
    END
  END Tile_X8Y12_WEN_SRAM5
  PIN Tile_X8Y12_WEN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 167.440 2324.560 168.000 ;
    END
  END Tile_X8Y12_WEN_SRAM6
  PIN Tile_X8Y12_WEN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 171.920 2324.560 172.480 ;
    END
  END Tile_X8Y12_WEN_SRAM7
  PIN Tile_X8Y2_A_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3049.200 2324.560 3049.760 ;
    END
  END Tile_X8Y2_A_SRAM0
  PIN Tile_X8Y2_A_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3053.680 2324.560 3054.240 ;
    END
  END Tile_X8Y2_A_SRAM1
  PIN Tile_X8Y2_A_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3058.160 2324.560 3058.720 ;
    END
  END Tile_X8Y2_A_SRAM2
  PIN Tile_X8Y2_A_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3062.640 2324.560 3063.200 ;
    END
  END Tile_X8Y2_A_SRAM3
  PIN Tile_X8Y2_A_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3067.120 2324.560 3067.680 ;
    END
  END Tile_X8Y2_A_SRAM4
  PIN Tile_X8Y2_A_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3071.600 2324.560 3072.160 ;
    END
  END Tile_X8Y2_A_SRAM5
  PIN Tile_X8Y2_A_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3076.080 2324.560 3076.640 ;
    END
  END Tile_X8Y2_A_SRAM6
  PIN Tile_X8Y2_A_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3080.560 2324.560 3081.120 ;
    END
  END Tile_X8Y2_A_SRAM7
  PIN Tile_X8Y2_A_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3085.040 2324.560 3085.600 ;
    END
  END Tile_X8Y2_A_SRAM8
  PIN Tile_X8Y2_CEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3004.400 2324.560 3004.960 ;
    END
  END Tile_X8Y2_CEN_SRAM
  PIN Tile_X8Y2_CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3125.360 2324.560 3125.920 ;
    END
  END Tile_X8Y2_CLK_SRAM
  PIN Tile_X8Y2_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2999.920 2324.560 3000.480 ;
    END
  END Tile_X8Y2_CONFIGURED_top
  PIN Tile_X8Y2_D_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3089.520 2324.560 3090.080 ;
    END
  END Tile_X8Y2_D_SRAM0
  PIN Tile_X8Y2_D_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3094.000 2324.560 3094.560 ;
    END
  END Tile_X8Y2_D_SRAM1
  PIN Tile_X8Y2_D_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3098.480 2324.560 3099.040 ;
    END
  END Tile_X8Y2_D_SRAM2
  PIN Tile_X8Y2_D_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3102.960 2324.560 3103.520 ;
    END
  END Tile_X8Y2_D_SRAM3
  PIN Tile_X8Y2_D_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3107.440 2324.560 3108.000 ;
    END
  END Tile_X8Y2_D_SRAM4
  PIN Tile_X8Y2_D_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3111.920 2324.560 3112.480 ;
    END
  END Tile_X8Y2_D_SRAM5
  PIN Tile_X8Y2_D_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3116.400 2324.560 3116.960 ;
    END
  END Tile_X8Y2_D_SRAM6
  PIN Tile_X8Y2_D_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3120.880 2324.560 3121.440 ;
    END
  END Tile_X8Y2_D_SRAM7
  PIN Tile_X8Y2_GWEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3008.880 2324.560 3009.440 ;
    END
  END Tile_X8Y2_GWEN_SRAM
  PIN Tile_X8Y2_Q_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2964.080 2324.560 2964.640 ;
    END
  END Tile_X8Y2_Q_SRAM0
  PIN Tile_X8Y2_Q_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2968.560 2324.560 2969.120 ;
    END
  END Tile_X8Y2_Q_SRAM1
  PIN Tile_X8Y2_Q_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2973.040 2324.560 2973.600 ;
    END
  END Tile_X8Y2_Q_SRAM2
  PIN Tile_X8Y2_Q_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2977.520 2324.560 2978.080 ;
    END
  END Tile_X8Y2_Q_SRAM3
  PIN Tile_X8Y2_Q_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.531500 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2982.000 2324.560 2982.560 ;
    END
  END Tile_X8Y2_Q_SRAM4
  PIN Tile_X8Y2_Q_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.528500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2986.480 2324.560 2987.040 ;
    END
  END Tile_X8Y2_Q_SRAM5
  PIN Tile_X8Y2_Q_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2990.960 2324.560 2991.520 ;
    END
  END Tile_X8Y2_Q_SRAM6
  PIN Tile_X8Y2_Q_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2995.440 2324.560 2996.000 ;
    END
  END Tile_X8Y2_Q_SRAM7
  PIN Tile_X8Y2_WEN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3013.360 2324.560 3013.920 ;
    END
  END Tile_X8Y2_WEN_SRAM0
  PIN Tile_X8Y2_WEN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3017.840 2324.560 3018.400 ;
    END
  END Tile_X8Y2_WEN_SRAM1
  PIN Tile_X8Y2_WEN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3022.320 2324.560 3022.880 ;
    END
  END Tile_X8Y2_WEN_SRAM2
  PIN Tile_X8Y2_WEN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3026.800 2324.560 3027.360 ;
    END
  END Tile_X8Y2_WEN_SRAM3
  PIN Tile_X8Y2_WEN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3031.280 2324.560 3031.840 ;
    END
  END Tile_X8Y2_WEN_SRAM4
  PIN Tile_X8Y2_WEN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3035.760 2324.560 3036.320 ;
    END
  END Tile_X8Y2_WEN_SRAM5
  PIN Tile_X8Y2_WEN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3040.240 2324.560 3040.800 ;
    END
  END Tile_X8Y2_WEN_SRAM6
  PIN Tile_X8Y2_WEN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 3044.720 2324.560 3045.280 ;
    END
  END Tile_X8Y2_WEN_SRAM7
  PIN Tile_X8Y4_A_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2474.640 2324.560 2475.200 ;
    END
  END Tile_X8Y4_A_SRAM0
  PIN Tile_X8Y4_A_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2479.120 2324.560 2479.680 ;
    END
  END Tile_X8Y4_A_SRAM1
  PIN Tile_X8Y4_A_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2483.600 2324.560 2484.160 ;
    END
  END Tile_X8Y4_A_SRAM2
  PIN Tile_X8Y4_A_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2488.080 2324.560 2488.640 ;
    END
  END Tile_X8Y4_A_SRAM3
  PIN Tile_X8Y4_A_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2492.560 2324.560 2493.120 ;
    END
  END Tile_X8Y4_A_SRAM4
  PIN Tile_X8Y4_A_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2497.040 2324.560 2497.600 ;
    END
  END Tile_X8Y4_A_SRAM5
  PIN Tile_X8Y4_A_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2501.520 2324.560 2502.080 ;
    END
  END Tile_X8Y4_A_SRAM6
  PIN Tile_X8Y4_A_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2506.000 2324.560 2506.560 ;
    END
  END Tile_X8Y4_A_SRAM7
  PIN Tile_X8Y4_A_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2510.480 2324.560 2511.040 ;
    END
  END Tile_X8Y4_A_SRAM8
  PIN Tile_X8Y4_CEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2429.840 2324.560 2430.400 ;
    END
  END Tile_X8Y4_CEN_SRAM
  PIN Tile_X8Y4_CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2550.800 2324.560 2551.360 ;
    END
  END Tile_X8Y4_CLK_SRAM
  PIN Tile_X8Y4_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2425.360 2324.560 2425.920 ;
    END
  END Tile_X8Y4_CONFIGURED_top
  PIN Tile_X8Y4_D_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2514.960 2324.560 2515.520 ;
    END
  END Tile_X8Y4_D_SRAM0
  PIN Tile_X8Y4_D_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2519.440 2324.560 2520.000 ;
    END
  END Tile_X8Y4_D_SRAM1
  PIN Tile_X8Y4_D_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2523.920 2324.560 2524.480 ;
    END
  END Tile_X8Y4_D_SRAM2
  PIN Tile_X8Y4_D_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2528.400 2324.560 2528.960 ;
    END
  END Tile_X8Y4_D_SRAM3
  PIN Tile_X8Y4_D_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2532.880 2324.560 2533.440 ;
    END
  END Tile_X8Y4_D_SRAM4
  PIN Tile_X8Y4_D_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2537.360 2324.560 2537.920 ;
    END
  END Tile_X8Y4_D_SRAM5
  PIN Tile_X8Y4_D_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2541.840 2324.560 2542.400 ;
    END
  END Tile_X8Y4_D_SRAM6
  PIN Tile_X8Y4_D_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2546.320 2324.560 2546.880 ;
    END
  END Tile_X8Y4_D_SRAM7
  PIN Tile_X8Y4_GWEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2434.320 2324.560 2434.880 ;
    END
  END Tile_X8Y4_GWEN_SRAM
  PIN Tile_X8Y4_Q_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2389.520 2324.560 2390.080 ;
    END
  END Tile_X8Y4_Q_SRAM0
  PIN Tile_X8Y4_Q_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2394.000 2324.560 2394.560 ;
    END
  END Tile_X8Y4_Q_SRAM1
  PIN Tile_X8Y4_Q_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2398.480 2324.560 2399.040 ;
    END
  END Tile_X8Y4_Q_SRAM2
  PIN Tile_X8Y4_Q_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2402.960 2324.560 2403.520 ;
    END
  END Tile_X8Y4_Q_SRAM3
  PIN Tile_X8Y4_Q_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.531500 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2407.440 2324.560 2408.000 ;
    END
  END Tile_X8Y4_Q_SRAM4
  PIN Tile_X8Y4_Q_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.528500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2411.920 2324.560 2412.480 ;
    END
  END Tile_X8Y4_Q_SRAM5
  PIN Tile_X8Y4_Q_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2416.400 2324.560 2416.960 ;
    END
  END Tile_X8Y4_Q_SRAM6
  PIN Tile_X8Y4_Q_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2420.880 2324.560 2421.440 ;
    END
  END Tile_X8Y4_Q_SRAM7
  PIN Tile_X8Y4_WEN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2438.800 2324.560 2439.360 ;
    END
  END Tile_X8Y4_WEN_SRAM0
  PIN Tile_X8Y4_WEN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2443.280 2324.560 2443.840 ;
    END
  END Tile_X8Y4_WEN_SRAM1
  PIN Tile_X8Y4_WEN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2447.760 2324.560 2448.320 ;
    END
  END Tile_X8Y4_WEN_SRAM2
  PIN Tile_X8Y4_WEN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2452.240 2324.560 2452.800 ;
    END
  END Tile_X8Y4_WEN_SRAM3
  PIN Tile_X8Y4_WEN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2456.720 2324.560 2457.280 ;
    END
  END Tile_X8Y4_WEN_SRAM4
  PIN Tile_X8Y4_WEN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2461.200 2324.560 2461.760 ;
    END
  END Tile_X8Y4_WEN_SRAM5
  PIN Tile_X8Y4_WEN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2465.680 2324.560 2466.240 ;
    END
  END Tile_X8Y4_WEN_SRAM6
  PIN Tile_X8Y4_WEN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 2470.160 2324.560 2470.720 ;
    END
  END Tile_X8Y4_WEN_SRAM7
  PIN Tile_X8Y6_A_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1900.080 2324.560 1900.640 ;
    END
  END Tile_X8Y6_A_SRAM0
  PIN Tile_X8Y6_A_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1904.560 2324.560 1905.120 ;
    END
  END Tile_X8Y6_A_SRAM1
  PIN Tile_X8Y6_A_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1909.040 2324.560 1909.600 ;
    END
  END Tile_X8Y6_A_SRAM2
  PIN Tile_X8Y6_A_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1913.520 2324.560 1914.080 ;
    END
  END Tile_X8Y6_A_SRAM3
  PIN Tile_X8Y6_A_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1918.000 2324.560 1918.560 ;
    END
  END Tile_X8Y6_A_SRAM4
  PIN Tile_X8Y6_A_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1922.480 2324.560 1923.040 ;
    END
  END Tile_X8Y6_A_SRAM5
  PIN Tile_X8Y6_A_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1926.960 2324.560 1927.520 ;
    END
  END Tile_X8Y6_A_SRAM6
  PIN Tile_X8Y6_A_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1931.440 2324.560 1932.000 ;
    END
  END Tile_X8Y6_A_SRAM7
  PIN Tile_X8Y6_A_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1935.920 2324.560 1936.480 ;
    END
  END Tile_X8Y6_A_SRAM8
  PIN Tile_X8Y6_CEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1855.280 2324.560 1855.840 ;
    END
  END Tile_X8Y6_CEN_SRAM
  PIN Tile_X8Y6_CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1976.240 2324.560 1976.800 ;
    END
  END Tile_X8Y6_CLK_SRAM
  PIN Tile_X8Y6_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1850.800 2324.560 1851.360 ;
    END
  END Tile_X8Y6_CONFIGURED_top
  PIN Tile_X8Y6_D_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1940.400 2324.560 1940.960 ;
    END
  END Tile_X8Y6_D_SRAM0
  PIN Tile_X8Y6_D_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1944.880 2324.560 1945.440 ;
    END
  END Tile_X8Y6_D_SRAM1
  PIN Tile_X8Y6_D_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1949.360 2324.560 1949.920 ;
    END
  END Tile_X8Y6_D_SRAM2
  PIN Tile_X8Y6_D_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1953.840 2324.560 1954.400 ;
    END
  END Tile_X8Y6_D_SRAM3
  PIN Tile_X8Y6_D_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1958.320 2324.560 1958.880 ;
    END
  END Tile_X8Y6_D_SRAM4
  PIN Tile_X8Y6_D_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1962.800 2324.560 1963.360 ;
    END
  END Tile_X8Y6_D_SRAM5
  PIN Tile_X8Y6_D_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1967.280 2324.560 1967.840 ;
    END
  END Tile_X8Y6_D_SRAM6
  PIN Tile_X8Y6_D_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1971.760 2324.560 1972.320 ;
    END
  END Tile_X8Y6_D_SRAM7
  PIN Tile_X8Y6_GWEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1859.760 2324.560 1860.320 ;
    END
  END Tile_X8Y6_GWEN_SRAM
  PIN Tile_X8Y6_Q_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1814.960 2324.560 1815.520 ;
    END
  END Tile_X8Y6_Q_SRAM0
  PIN Tile_X8Y6_Q_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1819.440 2324.560 1820.000 ;
    END
  END Tile_X8Y6_Q_SRAM1
  PIN Tile_X8Y6_Q_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1823.920 2324.560 1824.480 ;
    END
  END Tile_X8Y6_Q_SRAM2
  PIN Tile_X8Y6_Q_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1828.400 2324.560 1828.960 ;
    END
  END Tile_X8Y6_Q_SRAM3
  PIN Tile_X8Y6_Q_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.531500 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1832.880 2324.560 1833.440 ;
    END
  END Tile_X8Y6_Q_SRAM4
  PIN Tile_X8Y6_Q_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.528500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1837.360 2324.560 1837.920 ;
    END
  END Tile_X8Y6_Q_SRAM5
  PIN Tile_X8Y6_Q_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1841.840 2324.560 1842.400 ;
    END
  END Tile_X8Y6_Q_SRAM6
  PIN Tile_X8Y6_Q_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1846.320 2324.560 1846.880 ;
    END
  END Tile_X8Y6_Q_SRAM7
  PIN Tile_X8Y6_WEN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1864.240 2324.560 1864.800 ;
    END
  END Tile_X8Y6_WEN_SRAM0
  PIN Tile_X8Y6_WEN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1868.720 2324.560 1869.280 ;
    END
  END Tile_X8Y6_WEN_SRAM1
  PIN Tile_X8Y6_WEN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1873.200 2324.560 1873.760 ;
    END
  END Tile_X8Y6_WEN_SRAM2
  PIN Tile_X8Y6_WEN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1877.680 2324.560 1878.240 ;
    END
  END Tile_X8Y6_WEN_SRAM3
  PIN Tile_X8Y6_WEN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1882.160 2324.560 1882.720 ;
    END
  END Tile_X8Y6_WEN_SRAM4
  PIN Tile_X8Y6_WEN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1886.640 2324.560 1887.200 ;
    END
  END Tile_X8Y6_WEN_SRAM5
  PIN Tile_X8Y6_WEN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1891.120 2324.560 1891.680 ;
    END
  END Tile_X8Y6_WEN_SRAM6
  PIN Tile_X8Y6_WEN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1895.600 2324.560 1896.160 ;
    END
  END Tile_X8Y6_WEN_SRAM7
  PIN Tile_X8Y8_A_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1325.520 2324.560 1326.080 ;
    END
  END Tile_X8Y8_A_SRAM0
  PIN Tile_X8Y8_A_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1330.000 2324.560 1330.560 ;
    END
  END Tile_X8Y8_A_SRAM1
  PIN Tile_X8Y8_A_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1334.480 2324.560 1335.040 ;
    END
  END Tile_X8Y8_A_SRAM2
  PIN Tile_X8Y8_A_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1338.960 2324.560 1339.520 ;
    END
  END Tile_X8Y8_A_SRAM3
  PIN Tile_X8Y8_A_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1343.440 2324.560 1344.000 ;
    END
  END Tile_X8Y8_A_SRAM4
  PIN Tile_X8Y8_A_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1347.920 2324.560 1348.480 ;
    END
  END Tile_X8Y8_A_SRAM5
  PIN Tile_X8Y8_A_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1352.400 2324.560 1352.960 ;
    END
  END Tile_X8Y8_A_SRAM6
  PIN Tile_X8Y8_A_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1356.880 2324.560 1357.440 ;
    END
  END Tile_X8Y8_A_SRAM7
  PIN Tile_X8Y8_A_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1361.360 2324.560 1361.920 ;
    END
  END Tile_X8Y8_A_SRAM8
  PIN Tile_X8Y8_CEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1280.720 2324.560 1281.280 ;
    END
  END Tile_X8Y8_CEN_SRAM
  PIN Tile_X8Y8_CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1401.680 2324.560 1402.240 ;
    END
  END Tile_X8Y8_CLK_SRAM
  PIN Tile_X8Y8_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1276.240 2324.560 1276.800 ;
    END
  END Tile_X8Y8_CONFIGURED_top
  PIN Tile_X8Y8_D_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1365.840 2324.560 1366.400 ;
    END
  END Tile_X8Y8_D_SRAM0
  PIN Tile_X8Y8_D_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1370.320 2324.560 1370.880 ;
    END
  END Tile_X8Y8_D_SRAM1
  PIN Tile_X8Y8_D_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1374.800 2324.560 1375.360 ;
    END
  END Tile_X8Y8_D_SRAM2
  PIN Tile_X8Y8_D_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1379.280 2324.560 1379.840 ;
    END
  END Tile_X8Y8_D_SRAM3
  PIN Tile_X8Y8_D_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1383.760 2324.560 1384.320 ;
    END
  END Tile_X8Y8_D_SRAM4
  PIN Tile_X8Y8_D_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1388.240 2324.560 1388.800 ;
    END
  END Tile_X8Y8_D_SRAM5
  PIN Tile_X8Y8_D_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1392.720 2324.560 1393.280 ;
    END
  END Tile_X8Y8_D_SRAM6
  PIN Tile_X8Y8_D_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1397.200 2324.560 1397.760 ;
    END
  END Tile_X8Y8_D_SRAM7
  PIN Tile_X8Y8_GWEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1285.200 2324.560 1285.760 ;
    END
  END Tile_X8Y8_GWEN_SRAM
  PIN Tile_X8Y8_Q_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1240.400 2324.560 1240.960 ;
    END
  END Tile_X8Y8_Q_SRAM0
  PIN Tile_X8Y8_Q_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1244.880 2324.560 1245.440 ;
    END
  END Tile_X8Y8_Q_SRAM1
  PIN Tile_X8Y8_Q_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1249.360 2324.560 1249.920 ;
    END
  END Tile_X8Y8_Q_SRAM2
  PIN Tile_X8Y8_Q_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1253.840 2324.560 1254.400 ;
    END
  END Tile_X8Y8_Q_SRAM3
  PIN Tile_X8Y8_Q_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.531500 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1258.320 2324.560 1258.880 ;
    END
  END Tile_X8Y8_Q_SRAM4
  PIN Tile_X8Y8_Q_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.528500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1262.800 2324.560 1263.360 ;
    END
  END Tile_X8Y8_Q_SRAM5
  PIN Tile_X8Y8_Q_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1267.280 2324.560 1267.840 ;
    END
  END Tile_X8Y8_Q_SRAM6
  PIN Tile_X8Y8_Q_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1271.760 2324.560 1272.320 ;
    END
  END Tile_X8Y8_Q_SRAM7
  PIN Tile_X8Y8_WEN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1289.680 2324.560 1290.240 ;
    END
  END Tile_X8Y8_WEN_SRAM0
  PIN Tile_X8Y8_WEN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1294.160 2324.560 1294.720 ;
    END
  END Tile_X8Y8_WEN_SRAM1
  PIN Tile_X8Y8_WEN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1298.640 2324.560 1299.200 ;
    END
  END Tile_X8Y8_WEN_SRAM2
  PIN Tile_X8Y8_WEN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1303.120 2324.560 1303.680 ;
    END
  END Tile_X8Y8_WEN_SRAM3
  PIN Tile_X8Y8_WEN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1307.600 2324.560 1308.160 ;
    END
  END Tile_X8Y8_WEN_SRAM4
  PIN Tile_X8Y8_WEN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1312.080 2324.560 1312.640 ;
    END
  END Tile_X8Y8_WEN_SRAM5
  PIN Tile_X8Y8_WEN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1316.560 2324.560 1317.120 ;
    END
  END Tile_X8Y8_WEN_SRAM6
  PIN Tile_X8Y8_WEN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2323.440 1321.040 2324.560 1321.600 ;
    END
  END Tile_X8Y8_WEN_SRAM7
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.464000 ;
    ANTENNADIFFAREA 3.283200 ;
    PORT
      LAYER Metal2 ;
        RECT 3.920 0.000 4.480 0.560 ;
    END
  END UserCLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 19.440 651.280 21.040 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.440 651.280 121.040 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 19.440 364.000 21.040 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.440 364.000 121.040 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 19.440 76.720 21.040 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.440 76.720 121.040 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 19.440 3236.800 21.040 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.440 3236.800 121.040 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 19.440 2949.520 21.040 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.440 2949.520 121.040 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 19.440 2662.240 21.040 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.440 2662.240 121.040 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 19.440 2374.960 21.040 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.440 2374.960 121.040 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 19.440 2087.680 21.040 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.440 2087.680 121.040 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 19.440 1800.400 21.040 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.440 1800.400 121.040 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 19.440 1513.120 21.040 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.440 1513.120 121.040 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 19.440 1225.840 21.040 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.440 1225.840 121.040 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 19.440 938.560 21.040 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.440 938.560 121.040 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.240 3524.080 163.840 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.240 3524.080 263.840 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.240 3524.080 363.840 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.240 651.280 163.840 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.240 651.280 263.840 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.240 651.280 363.840 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.240 364.000 163.840 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.240 364.000 263.840 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.240 364.000 363.840 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.240 76.720 163.840 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.240 76.720 263.840 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.240 76.720 363.840 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.240 5.600 163.840 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.240 5.600 263.840 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.240 5.600 363.840 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.240 3236.800 163.840 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.240 3236.800 263.840 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.240 3236.800 363.840 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.240 2949.520 163.840 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.240 2949.520 263.840 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.240 2949.520 363.840 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.240 2662.240 163.840 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.240 2662.240 263.840 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.240 2662.240 363.840 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.240 2374.960 163.840 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.240 2374.960 263.840 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.240 2374.960 363.840 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.240 2087.680 163.840 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.240 2087.680 263.840 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.240 2087.680 363.840 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.240 1800.400 163.840 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.240 1800.400 263.840 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.240 1800.400 363.840 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.240 1513.120 163.840 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.240 1513.120 263.840 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.240 1513.120 363.840 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.240 1225.840 163.840 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.240 1225.840 263.840 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.240 1225.840 363.840 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.240 938.560 163.840 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.240 938.560 263.840 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.240 938.560 363.840 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.520 3524.080 451.120 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.520 3524.080 551.120 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 649.520 3524.080 651.120 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.520 651.280 451.120 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.520 651.280 551.120 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 649.520 651.280 651.120 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.520 364.000 451.120 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.520 364.000 551.120 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 649.520 364.000 651.120 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.520 76.720 451.120 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.520 76.720 551.120 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 649.520 76.720 651.120 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.520 5.600 451.120 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.520 5.600 551.120 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 649.520 5.600 651.120 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.520 3236.800 451.120 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.520 3236.800 551.120 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 649.520 3236.800 651.120 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.520 2949.520 451.120 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.520 2949.520 551.120 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 649.520 2949.520 651.120 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.520 2662.240 451.120 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.520 2662.240 551.120 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 649.520 2662.240 651.120 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.520 2374.960 451.120 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.520 2374.960 551.120 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 649.520 2374.960 651.120 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.520 2087.680 451.120 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.520 2087.680 551.120 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 649.520 2087.680 651.120 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.520 1800.400 451.120 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.520 1800.400 551.120 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 649.520 1800.400 651.120 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.520 1513.120 451.120 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.520 1513.120 551.120 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 649.520 1513.120 651.120 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.520 1225.840 451.120 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.520 1225.840 551.120 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 649.520 1225.840 651.120 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.520 938.560 451.120 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 549.520 938.560 551.120 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 649.520 938.560 651.120 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.800 3524.080 738.400 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 836.800 3524.080 838.400 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 936.800 3524.080 938.400 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.800 651.280 738.400 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 836.800 651.280 838.400 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 936.800 651.280 938.400 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.800 364.000 738.400 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 836.800 364.000 838.400 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 936.800 364.000 938.400 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.800 76.720 738.400 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 836.800 76.720 838.400 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 936.800 76.720 938.400 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.800 5.600 738.400 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 836.800 5.600 838.400 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 936.800 5.600 938.400 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.800 3236.800 738.400 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 836.800 3236.800 838.400 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 936.800 3236.800 938.400 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.800 2949.520 738.400 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 836.800 2949.520 838.400 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 936.800 2949.520 938.400 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.800 2662.240 738.400 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 836.800 2662.240 838.400 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 936.800 2662.240 938.400 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.800 2374.960 738.400 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 836.800 2374.960 838.400 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 936.800 2374.960 938.400 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.800 2087.680 738.400 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 836.800 2087.680 838.400 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 936.800 2087.680 938.400 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.800 1800.400 738.400 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 836.800 1800.400 838.400 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 936.800 1800.400 938.400 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.800 1513.120 738.400 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 836.800 1513.120 838.400 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 936.800 1513.120 938.400 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.800 1225.840 738.400 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 836.800 1225.840 838.400 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 936.800 1225.840 938.400 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 736.800 938.560 738.400 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 836.800 938.560 838.400 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 936.800 938.560 938.400 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.080 3524.080 1025.680 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1124.080 3524.080 1125.680 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1224.080 3524.080 1225.680 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.080 651.280 1025.680 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1124.080 651.280 1125.680 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1224.080 651.280 1225.680 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.080 364.000 1025.680 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1124.080 364.000 1125.680 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1224.080 364.000 1225.680 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.080 76.720 1025.680 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1124.080 76.720 1125.680 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1224.080 76.720 1225.680 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.080 5.600 1025.680 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1124.080 5.600 1125.680 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1224.080 5.600 1225.680 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.080 3236.800 1025.680 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1124.080 3236.800 1125.680 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1224.080 3236.800 1225.680 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.080 2949.520 1025.680 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1124.080 2949.520 1125.680 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1224.080 2949.520 1225.680 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.080 2662.240 1025.680 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1124.080 2662.240 1125.680 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1224.080 2662.240 1225.680 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.080 2374.960 1025.680 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1124.080 2374.960 1125.680 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1224.080 2374.960 1225.680 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.080 2087.680 1025.680 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1124.080 2087.680 1125.680 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1224.080 2087.680 1225.680 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.080 1800.400 1025.680 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1124.080 1800.400 1125.680 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1224.080 1800.400 1225.680 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.080 1513.120 1025.680 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1124.080 1513.120 1125.680 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1224.080 1513.120 1225.680 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.080 1225.840 1025.680 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1124.080 1225.840 1125.680 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1224.080 1225.840 1225.680 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.080 938.560 1025.680 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1124.080 938.560 1125.680 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1224.080 938.560 1225.680 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.080 3524.080 1347.680 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1446.080 3524.080 1447.680 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 3524.080 1547.680 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.080 651.280 1347.680 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1446.080 651.280 1447.680 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 651.280 1547.680 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.080 364.000 1347.680 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1446.080 364.000 1447.680 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 364.000 1547.680 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.080 76.720 1347.680 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1446.080 76.720 1447.680 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 76.720 1547.680 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.080 5.600 1347.680 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1446.080 5.600 1447.680 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 5.600 1547.680 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.080 3236.800 1347.680 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1446.080 3236.800 1447.680 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 3236.800 1547.680 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.080 2949.520 1347.680 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1446.080 2949.520 1447.680 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 2949.520 1547.680 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.080 2662.240 1347.680 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1446.080 2662.240 1447.680 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 2662.240 1547.680 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.080 2374.960 1347.680 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1446.080 2374.960 1447.680 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 2374.960 1547.680 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.080 2087.680 1347.680 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1446.080 2087.680 1447.680 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 2087.680 1547.680 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.080 1800.400 1347.680 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1446.080 1800.400 1447.680 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 1800.400 1547.680 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.080 1513.120 1347.680 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1446.080 1513.120 1447.680 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 1513.120 1547.680 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.080 1225.840 1347.680 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1446.080 1225.840 1447.680 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 1225.840 1547.680 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1346.080 938.560 1347.680 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1446.080 938.560 1447.680 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 938.560 1547.680 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1633.360 3524.080 1634.960 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1733.360 3524.080 1734.960 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1833.360 3524.080 1834.960 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1633.360 76.720 1634.960 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1733.360 76.720 1734.960 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1833.360 76.720 1834.960 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1633.360 5.600 1634.960 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1733.360 5.600 1734.960 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1833.360 5.600 1834.960 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1633.360 2949.520 1634.960 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1733.360 2949.520 1734.960 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1833.360 2949.520 1834.960 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1633.360 2374.960 1634.960 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1733.360 2374.960 1734.960 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1833.360 2374.960 1834.960 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1633.360 1800.400 1634.960 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1733.360 1800.400 1734.960 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1833.360 1800.400 1834.960 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1633.360 1225.840 1634.960 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1733.360 1225.840 1734.960 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1833.360 1225.840 1834.960 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1633.360 651.280 1634.960 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1733.360 651.280 1734.960 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1833.360 651.280 1834.960 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1897.120 3524.080 1898.720 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1997.120 3524.080 1998.720 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2097.120 3524.080 2098.720 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1897.120 651.280 1898.720 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1997.120 651.280 1998.720 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2097.120 651.280 2098.720 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1897.120 364.000 1898.720 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1997.120 364.000 1998.720 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2097.120 364.000 2098.720 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1897.120 76.720 1898.720 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1997.120 76.720 1998.720 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2097.120 76.720 2098.720 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1897.120 5.600 1898.720 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1997.120 5.600 1998.720 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2097.120 5.600 2098.720 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1897.120 3236.800 1898.720 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1997.120 3236.800 1998.720 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2097.120 3236.800 2098.720 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1897.120 2949.520 1898.720 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1997.120 2949.520 1998.720 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2097.120 2949.520 2098.720 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1897.120 2662.240 1898.720 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1997.120 2662.240 1998.720 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2097.120 2662.240 2098.720 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1897.120 2374.960 1898.720 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1997.120 2374.960 1998.720 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2097.120 2374.960 2098.720 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1897.120 2087.680 1898.720 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1997.120 2087.680 1998.720 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2097.120 2087.680 2098.720 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1897.120 1800.400 1898.720 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1997.120 1800.400 1998.720 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2097.120 1800.400 2098.720 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1897.120 1513.120 1898.720 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1997.120 1513.120 1998.720 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2097.120 1513.120 2098.720 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1897.120 1225.840 1898.720 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1997.120 1225.840 1998.720 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2097.120 1225.840 2098.720 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1897.120 938.560 1898.720 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1997.120 938.560 1998.720 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2097.120 938.560 2098.720 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2184.400 3524.080 2186.000 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2284.400 3524.080 2286.000 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2184.400 76.720 2186.000 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2284.400 76.720 2286.000 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2184.400 5.600 2186.000 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2284.400 5.600 2286.000 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2184.400 2949.520 2186.000 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2284.400 2949.520 2286.000 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2184.400 2374.960 2186.000 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2284.400 2374.960 2286.000 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2184.400 1800.400 2186.000 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2284.400 1800.400 2286.000 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2184.400 1225.840 2186.000 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2284.400 1225.840 2286.000 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2184.400 651.280 2186.000 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2284.400 651.280 2286.000 1225.840 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.740 651.280 24.340 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.740 651.280 124.340 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 22.740 364.000 24.340 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.740 364.000 124.340 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 22.740 76.720 24.340 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.740 76.720 124.340 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 22.740 3236.800 24.340 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.740 3236.800 124.340 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 22.740 2949.520 24.340 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.740 2949.520 124.340 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 22.740 2662.240 24.340 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.740 2662.240 124.340 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 22.740 2374.960 24.340 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.740 2374.960 124.340 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 22.740 2087.680 24.340 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.740 2087.680 124.340 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 22.740 1800.400 24.340 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.740 1800.400 124.340 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 22.740 1513.120 24.340 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.740 1513.120 124.340 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 22.740 1225.840 24.340 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.740 1225.840 124.340 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 22.740 938.560 24.340 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.740 938.560 124.340 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.540 3524.080 167.140 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 265.540 3524.080 267.140 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.540 3524.080 367.140 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.540 651.280 167.140 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 265.540 651.280 267.140 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.540 651.280 367.140 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.540 364.000 167.140 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 265.540 364.000 267.140 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.540 364.000 367.140 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.540 76.720 167.140 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 265.540 76.720 267.140 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.540 76.720 367.140 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.540 5.600 167.140 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 265.540 5.600 267.140 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.540 5.600 367.140 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.540 3236.800 167.140 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 265.540 3236.800 267.140 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.540 3236.800 367.140 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.540 2949.520 167.140 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 265.540 2949.520 267.140 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.540 2949.520 367.140 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.540 2662.240 167.140 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 265.540 2662.240 267.140 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.540 2662.240 367.140 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.540 2374.960 167.140 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 265.540 2374.960 267.140 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.540 2374.960 367.140 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.540 2087.680 167.140 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 265.540 2087.680 267.140 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.540 2087.680 367.140 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.540 1800.400 167.140 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 265.540 1800.400 267.140 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.540 1800.400 367.140 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.540 1513.120 167.140 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 265.540 1513.120 267.140 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.540 1513.120 367.140 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.540 1225.840 167.140 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 265.540 1225.840 267.140 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.540 1225.840 367.140 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.540 938.560 167.140 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 265.540 938.560 267.140 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.540 938.560 367.140 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 452.820 3524.080 454.420 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 552.820 3524.080 554.420 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 652.820 3524.080 654.420 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 452.820 651.280 454.420 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 552.820 651.280 554.420 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 652.820 651.280 654.420 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 452.820 364.000 454.420 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 552.820 364.000 554.420 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 652.820 364.000 654.420 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 452.820 76.720 454.420 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 552.820 76.720 554.420 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 652.820 76.720 654.420 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 452.820 5.600 454.420 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 552.820 5.600 554.420 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 652.820 5.600 654.420 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 452.820 3236.800 454.420 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 552.820 3236.800 554.420 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 652.820 3236.800 654.420 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 452.820 2949.520 454.420 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 552.820 2949.520 554.420 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 652.820 2949.520 654.420 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 452.820 2662.240 454.420 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 552.820 2662.240 554.420 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 652.820 2662.240 654.420 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 452.820 2374.960 454.420 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 552.820 2374.960 554.420 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 652.820 2374.960 654.420 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 452.820 2087.680 454.420 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 552.820 2087.680 554.420 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 652.820 2087.680 654.420 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 452.820 1800.400 454.420 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 552.820 1800.400 554.420 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 652.820 1800.400 654.420 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 452.820 1513.120 454.420 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 552.820 1513.120 554.420 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 652.820 1513.120 654.420 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 452.820 1225.840 454.420 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 552.820 1225.840 554.420 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 652.820 1225.840 654.420 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 452.820 938.560 454.420 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 552.820 938.560 554.420 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 652.820 938.560 654.420 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 740.100 3524.080 741.700 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 840.100 3524.080 841.700 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.100 3524.080 941.700 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 740.100 651.280 741.700 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 840.100 651.280 841.700 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.100 651.280 941.700 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 740.100 364.000 741.700 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 840.100 364.000 841.700 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.100 364.000 941.700 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 740.100 76.720 741.700 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 840.100 76.720 841.700 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.100 76.720 941.700 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 740.100 5.600 741.700 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 840.100 5.600 841.700 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.100 5.600 941.700 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 740.100 3236.800 741.700 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 840.100 3236.800 841.700 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.100 3236.800 941.700 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 740.100 2949.520 741.700 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 840.100 2949.520 841.700 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.100 2949.520 941.700 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 740.100 2662.240 741.700 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 840.100 2662.240 841.700 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.100 2662.240 941.700 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 740.100 2374.960 741.700 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 840.100 2374.960 841.700 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.100 2374.960 941.700 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 740.100 2087.680 741.700 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 840.100 2087.680 841.700 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.100 2087.680 941.700 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 740.100 1800.400 741.700 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 840.100 1800.400 841.700 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.100 1800.400 941.700 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 740.100 1513.120 741.700 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 840.100 1513.120 841.700 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.100 1513.120 941.700 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 740.100 1225.840 741.700 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 840.100 1225.840 841.700 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.100 1225.840 941.700 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 740.100 938.560 741.700 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 840.100 938.560 841.700 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.100 938.560 941.700 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1027.380 3524.080 1028.980 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.380 3524.080 1128.980 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1227.380 3524.080 1228.980 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1027.380 651.280 1028.980 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.380 651.280 1128.980 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1227.380 651.280 1228.980 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1027.380 364.000 1028.980 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.380 364.000 1128.980 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1227.380 364.000 1228.980 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1027.380 76.720 1028.980 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.380 76.720 1128.980 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1227.380 76.720 1228.980 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1027.380 5.600 1028.980 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.380 5.600 1128.980 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1227.380 5.600 1228.980 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1027.380 3236.800 1028.980 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.380 3236.800 1128.980 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1227.380 3236.800 1228.980 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1027.380 2949.520 1028.980 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.380 2949.520 1128.980 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1227.380 2949.520 1228.980 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1027.380 2662.240 1028.980 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.380 2662.240 1128.980 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1227.380 2662.240 1228.980 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1027.380 2374.960 1028.980 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.380 2374.960 1128.980 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1227.380 2374.960 1228.980 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1027.380 2087.680 1028.980 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.380 2087.680 1128.980 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1227.380 2087.680 1228.980 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1027.380 1800.400 1028.980 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.380 1800.400 1128.980 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1227.380 1800.400 1228.980 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1027.380 1513.120 1028.980 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.380 1513.120 1128.980 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1227.380 1513.120 1228.980 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1027.380 1225.840 1028.980 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.380 1225.840 1128.980 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1227.380 1225.840 1228.980 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1027.380 938.560 1028.980 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1127.380 938.560 1128.980 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1227.380 938.560 1228.980 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1349.380 3524.080 1350.980 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1449.380 3524.080 1450.980 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1549.380 3524.080 1550.980 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1349.380 651.280 1350.980 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1449.380 651.280 1450.980 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1549.380 651.280 1550.980 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1349.380 364.000 1350.980 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1449.380 364.000 1450.980 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1549.380 364.000 1550.980 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1349.380 76.720 1350.980 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1449.380 76.720 1450.980 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1549.380 76.720 1550.980 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1349.380 5.600 1350.980 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1449.380 5.600 1450.980 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1549.380 5.600 1550.980 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1349.380 3236.800 1350.980 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1449.380 3236.800 1450.980 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1549.380 3236.800 1550.980 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1349.380 2949.520 1350.980 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1449.380 2949.520 1450.980 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1549.380 2949.520 1550.980 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1349.380 2662.240 1350.980 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1449.380 2662.240 1450.980 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1549.380 2662.240 1550.980 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1349.380 2374.960 1350.980 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1449.380 2374.960 1450.980 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1549.380 2374.960 1550.980 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1349.380 2087.680 1350.980 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1449.380 2087.680 1450.980 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1549.380 2087.680 1550.980 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1349.380 1800.400 1350.980 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1449.380 1800.400 1450.980 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1549.380 1800.400 1550.980 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1349.380 1513.120 1350.980 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1449.380 1513.120 1450.980 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1549.380 1513.120 1550.980 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1349.380 1225.840 1350.980 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1449.380 1225.840 1450.980 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1549.380 1225.840 1550.980 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1349.380 938.560 1350.980 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1449.380 938.560 1450.980 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1549.380 938.560 1550.980 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1636.660 3524.080 1638.260 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1736.660 3524.080 1738.260 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1836.660 3524.080 1838.260 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1636.660 76.720 1638.260 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1736.660 76.720 1738.260 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1836.660 76.720 1838.260 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1636.660 5.600 1638.260 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1736.660 5.600 1738.260 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1836.660 5.600 1838.260 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1636.660 2949.520 1638.260 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1736.660 2949.520 1738.260 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1836.660 2949.520 1838.260 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1636.660 2374.960 1638.260 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1736.660 2374.960 1738.260 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1836.660 2374.960 1838.260 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1636.660 1800.400 1638.260 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1736.660 1800.400 1738.260 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1836.660 1800.400 1838.260 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1636.660 1225.840 1638.260 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1736.660 1225.840 1738.260 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1836.660 1225.840 1838.260 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1636.660 651.280 1638.260 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1736.660 651.280 1738.260 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1836.660 651.280 1838.260 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1900.420 3524.080 1902.020 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2000.420 3524.080 2002.020 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2100.420 3524.080 2102.020 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1900.420 651.280 1902.020 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2000.420 651.280 2002.020 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2100.420 651.280 2102.020 938.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1900.420 364.000 1902.020 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2000.420 364.000 2002.020 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2100.420 364.000 2102.020 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1900.420 76.720 1902.020 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2000.420 76.720 2002.020 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2100.420 76.720 2102.020 364.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1900.420 5.600 1902.020 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2000.420 5.600 2002.020 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2100.420 5.600 2102.020 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1900.420 3236.800 1902.020 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2000.420 3236.800 2002.020 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2100.420 3236.800 2102.020 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1900.420 2949.520 1902.020 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2000.420 2949.520 2002.020 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2100.420 2949.520 2102.020 3236.800 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1900.420 2662.240 1902.020 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2000.420 2662.240 2002.020 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2100.420 2662.240 2102.020 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1900.420 2374.960 1902.020 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2000.420 2374.960 2002.020 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2100.420 2374.960 2102.020 2662.240 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1900.420 2087.680 1902.020 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2000.420 2087.680 2002.020 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2100.420 2087.680 2102.020 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1900.420 1800.400 1902.020 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2000.420 1800.400 2002.020 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2100.420 1800.400 2102.020 2087.680 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1900.420 1513.120 1902.020 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2000.420 1513.120 2002.020 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2100.420 1513.120 2102.020 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1900.420 1225.840 1902.020 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2000.420 1225.840 2002.020 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2100.420 1225.840 2102.020 1513.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1900.420 938.560 1902.020 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2000.420 938.560 2002.020 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2100.420 938.560 2102.020 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2187.700 3524.080 2189.300 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2287.700 3524.080 2289.300 3595.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2187.700 76.720 2189.300 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2287.700 76.720 2289.300 651.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2187.700 5.600 2189.300 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2287.700 5.600 2289.300 76.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2187.700 2949.520 2189.300 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2287.700 2949.520 2289.300 3524.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2187.700 2374.960 2189.300 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2287.700 2374.960 2289.300 2949.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2187.700 1800.400 2189.300 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2287.700 1800.400 2289.300 2374.960 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2187.700 1225.840 2189.300 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2287.700 1225.840 2289.300 1800.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2187.700 651.280 2189.300 1225.840 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2287.700 651.280 2289.300 1225.840 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 3.490 9.090 2321.070 3591.150 ;
      LAYER Metal1 ;
        RECT 3.920 9.220 2320.640 3591.020 ;
      LAYER Metal2 ;
        RECT 1.820 0.860 2323.300 3595.670 ;
        RECT 1.820 0.090 3.620 0.860 ;
        RECT 4.780 0.090 10.340 0.860 ;
        RECT 11.500 0.090 17.060 0.860 ;
        RECT 18.220 0.090 23.780 0.860 ;
        RECT 24.940 0.090 30.500 0.860 ;
        RECT 31.660 0.090 37.220 0.860 ;
        RECT 38.380 0.090 43.940 0.860 ;
        RECT 45.100 0.090 50.660 0.860 ;
        RECT 51.820 0.090 57.380 0.860 ;
        RECT 58.540 0.090 64.100 0.860 ;
        RECT 65.260 0.090 70.820 0.860 ;
        RECT 71.980 0.090 77.540 0.860 ;
        RECT 78.700 0.090 84.260 0.860 ;
        RECT 85.420 0.090 90.980 0.860 ;
        RECT 92.140 0.090 97.700 0.860 ;
        RECT 98.860 0.090 104.420 0.860 ;
        RECT 105.580 0.090 111.140 0.860 ;
        RECT 112.300 0.090 117.860 0.860 ;
        RECT 119.020 0.090 124.580 0.860 ;
        RECT 125.740 0.090 131.300 0.860 ;
        RECT 132.460 0.090 138.020 0.860 ;
        RECT 139.180 0.090 149.780 0.860 ;
        RECT 150.940 0.090 159.860 0.860 ;
        RECT 161.020 0.090 169.940 0.860 ;
        RECT 171.100 0.090 180.020 0.860 ;
        RECT 181.180 0.090 190.100 0.860 ;
        RECT 191.260 0.090 200.180 0.860 ;
        RECT 201.340 0.090 210.260 0.860 ;
        RECT 211.420 0.090 230.420 0.860 ;
        RECT 231.580 0.090 240.500 0.860 ;
        RECT 241.660 0.090 250.580 0.860 ;
        RECT 251.740 0.090 260.660 0.860 ;
        RECT 261.820 0.090 270.740 0.860 ;
        RECT 271.900 0.090 280.820 0.860 ;
        RECT 281.980 0.090 290.900 0.860 ;
        RECT 292.060 0.090 300.980 0.860 ;
        RECT 302.140 0.090 311.060 0.860 ;
        RECT 312.220 0.090 321.140 0.860 ;
        RECT 322.300 0.090 331.220 0.860 ;
        RECT 332.380 0.090 341.300 0.860 ;
        RECT 342.460 0.090 351.380 0.860 ;
        RECT 352.540 0.090 361.460 0.860 ;
        RECT 362.620 0.090 371.540 0.860 ;
        RECT 372.700 0.090 381.620 0.860 ;
        RECT 382.780 0.090 391.700 0.860 ;
        RECT 392.860 0.090 401.780 0.860 ;
        RECT 402.940 0.090 411.860 0.860 ;
        RECT 413.020 0.090 421.940 0.860 ;
        RECT 423.100 0.090 452.740 0.860 ;
        RECT 453.900 0.090 466.180 0.860 ;
        RECT 467.340 0.090 479.620 0.860 ;
        RECT 480.780 0.090 493.060 0.860 ;
        RECT 494.220 0.090 506.500 0.860 ;
        RECT 507.660 0.090 519.940 0.860 ;
        RECT 521.100 0.090 533.380 0.860 ;
        RECT 534.540 0.090 546.820 0.860 ;
        RECT 547.980 0.090 560.260 0.860 ;
        RECT 561.420 0.090 573.700 0.860 ;
        RECT 574.860 0.090 587.140 0.860 ;
        RECT 588.300 0.090 600.580 0.860 ;
        RECT 601.740 0.090 614.020 0.860 ;
        RECT 615.180 0.090 627.460 0.860 ;
        RECT 628.620 0.090 640.900 0.860 ;
        RECT 642.060 0.090 654.340 0.860 ;
        RECT 655.500 0.090 667.780 0.860 ;
        RECT 668.940 0.090 681.220 0.860 ;
        RECT 682.380 0.090 694.660 0.860 ;
        RECT 695.820 0.090 708.100 0.860 ;
        RECT 709.260 0.090 740.020 0.860 ;
        RECT 741.180 0.090 753.460 0.860 ;
        RECT 754.620 0.090 766.900 0.860 ;
        RECT 768.060 0.090 780.340 0.860 ;
        RECT 781.500 0.090 793.780 0.860 ;
        RECT 794.940 0.090 807.220 0.860 ;
        RECT 808.380 0.090 820.660 0.860 ;
        RECT 821.820 0.090 834.100 0.860 ;
        RECT 835.260 0.090 847.540 0.860 ;
        RECT 848.700 0.090 860.980 0.860 ;
        RECT 862.140 0.090 874.420 0.860 ;
        RECT 875.580 0.090 887.860 0.860 ;
        RECT 889.020 0.090 901.300 0.860 ;
        RECT 902.460 0.090 914.740 0.860 ;
        RECT 915.900 0.090 928.180 0.860 ;
        RECT 929.340 0.090 941.620 0.860 ;
        RECT 942.780 0.090 955.060 0.860 ;
        RECT 956.220 0.090 968.500 0.860 ;
        RECT 969.660 0.090 981.940 0.860 ;
        RECT 983.100 0.090 995.380 0.860 ;
        RECT 996.540 0.090 1034.020 0.860 ;
        RECT 1035.180 0.090 1048.580 0.860 ;
        RECT 1049.740 0.090 1063.140 0.860 ;
        RECT 1064.300 0.090 1077.700 0.860 ;
        RECT 1078.860 0.090 1092.260 0.860 ;
        RECT 1093.420 0.090 1106.820 0.860 ;
        RECT 1107.980 0.090 1121.380 0.860 ;
        RECT 1122.540 0.090 1135.940 0.860 ;
        RECT 1137.100 0.090 1150.500 0.860 ;
        RECT 1151.660 0.090 1165.060 0.860 ;
        RECT 1166.220 0.090 1179.620 0.860 ;
        RECT 1180.780 0.090 1194.180 0.860 ;
        RECT 1195.340 0.090 1208.740 0.860 ;
        RECT 1209.900 0.090 1223.300 0.860 ;
        RECT 1224.460 0.090 1237.860 0.860 ;
        RECT 1239.020 0.090 1252.420 0.860 ;
        RECT 1253.580 0.090 1266.980 0.860 ;
        RECT 1268.140 0.090 1281.540 0.860 ;
        RECT 1282.700 0.090 1296.100 0.860 ;
        RECT 1297.260 0.090 1310.660 0.860 ;
        RECT 1311.820 0.090 1349.300 0.860 ;
        RECT 1350.460 0.090 1362.740 0.860 ;
        RECT 1363.900 0.090 1376.180 0.860 ;
        RECT 1377.340 0.090 1389.620 0.860 ;
        RECT 1390.780 0.090 1403.060 0.860 ;
        RECT 1404.220 0.090 1416.500 0.860 ;
        RECT 1417.660 0.090 1429.940 0.860 ;
        RECT 1431.100 0.090 1443.380 0.860 ;
        RECT 1444.540 0.090 1456.820 0.860 ;
        RECT 1457.980 0.090 1470.260 0.860 ;
        RECT 1471.420 0.090 1483.700 0.860 ;
        RECT 1484.860 0.090 1497.140 0.860 ;
        RECT 1498.300 0.090 1510.580 0.860 ;
        RECT 1511.740 0.090 1524.020 0.860 ;
        RECT 1525.180 0.090 1537.460 0.860 ;
        RECT 1538.620 0.090 1550.900 0.860 ;
        RECT 1552.060 0.090 1564.340 0.860 ;
        RECT 1565.500 0.090 1577.780 0.860 ;
        RECT 1578.940 0.090 1591.220 0.860 ;
        RECT 1592.380 0.090 1604.660 0.860 ;
        RECT 1605.820 0.090 1634.340 0.860 ;
        RECT 1635.500 0.090 1646.660 0.860 ;
        RECT 1647.820 0.090 1658.980 0.860 ;
        RECT 1660.140 0.090 1671.300 0.860 ;
        RECT 1672.460 0.090 1683.620 0.860 ;
        RECT 1684.780 0.090 1695.940 0.860 ;
        RECT 1697.100 0.090 1708.260 0.860 ;
        RECT 1709.420 0.090 1720.580 0.860 ;
        RECT 1721.740 0.090 1732.900 0.860 ;
        RECT 1734.060 0.090 1745.220 0.860 ;
        RECT 1746.380 0.090 1757.540 0.860 ;
        RECT 1758.700 0.090 1769.860 0.860 ;
        RECT 1771.020 0.090 1782.180 0.860 ;
        RECT 1783.340 0.090 1794.500 0.860 ;
        RECT 1795.660 0.090 1806.820 0.860 ;
        RECT 1807.980 0.090 1819.140 0.860 ;
        RECT 1820.300 0.090 1831.460 0.860 ;
        RECT 1832.620 0.090 1843.780 0.860 ;
        RECT 1844.940 0.090 1856.100 0.860 ;
        RECT 1857.260 0.090 1868.420 0.860 ;
        RECT 1869.580 0.090 1900.340 0.860 ;
        RECT 1901.500 0.090 1913.780 0.860 ;
        RECT 1914.940 0.090 1927.220 0.860 ;
        RECT 1928.380 0.090 1940.660 0.860 ;
        RECT 1941.820 0.090 1954.100 0.860 ;
        RECT 1955.260 0.090 1967.540 0.860 ;
        RECT 1968.700 0.090 1980.980 0.860 ;
        RECT 1982.140 0.090 1994.420 0.860 ;
        RECT 1995.580 0.090 2007.860 0.860 ;
        RECT 2009.020 0.090 2021.300 0.860 ;
        RECT 2022.460 0.090 2034.740 0.860 ;
        RECT 2035.900 0.090 2048.180 0.860 ;
        RECT 2049.340 0.090 2061.620 0.860 ;
        RECT 2062.780 0.090 2075.060 0.860 ;
        RECT 2076.220 0.090 2088.500 0.860 ;
        RECT 2089.660 0.090 2101.940 0.860 ;
        RECT 2103.100 0.090 2115.380 0.860 ;
        RECT 2116.540 0.090 2128.820 0.860 ;
        RECT 2129.980 0.090 2142.260 0.860 ;
        RECT 2143.420 0.090 2155.700 0.860 ;
        RECT 2156.860 0.090 2183.140 0.860 ;
        RECT 2184.300 0.090 2189.860 0.860 ;
        RECT 2191.020 0.090 2196.580 0.860 ;
        RECT 2197.740 0.090 2203.300 0.860 ;
        RECT 2204.460 0.090 2210.020 0.860 ;
        RECT 2211.180 0.090 2216.740 0.860 ;
        RECT 2217.900 0.090 2223.460 0.860 ;
        RECT 2224.620 0.090 2230.180 0.860 ;
        RECT 2231.340 0.090 2240.820 0.860 ;
        RECT 2241.980 0.090 2243.620 0.860 ;
        RECT 2244.780 0.090 2250.340 0.860 ;
        RECT 2251.500 0.090 2257.060 0.860 ;
        RECT 2258.220 0.090 2263.780 0.860 ;
        RECT 2264.940 0.090 2270.500 0.860 ;
        RECT 2271.660 0.090 2277.220 0.860 ;
        RECT 2278.380 0.090 2283.940 0.860 ;
        RECT 2285.100 0.090 2290.660 0.860 ;
        RECT 2291.820 0.090 2297.380 0.860 ;
        RECT 2298.540 0.090 2304.100 0.860 ;
        RECT 2305.260 0.090 2310.820 0.860 ;
        RECT 2311.980 0.090 2323.300 0.860 ;
      LAYER Metal3 ;
        RECT 0.560 3594.380 2324.000 3595.620 ;
        RECT 0.860 3593.220 2324.000 3594.380 ;
        RECT 0.560 3592.140 2324.000 3593.220 ;
        RECT 0.860 3590.980 2324.000 3592.140 ;
        RECT 0.560 3589.900 2324.000 3590.980 ;
        RECT 0.860 3588.740 2324.000 3589.900 ;
        RECT 0.560 3587.660 2324.000 3588.740 ;
        RECT 0.860 3586.500 2324.000 3587.660 ;
        RECT 0.560 3585.420 2324.000 3586.500 ;
        RECT 0.860 3584.260 2324.000 3585.420 ;
        RECT 0.560 3583.180 2324.000 3584.260 ;
        RECT 0.860 3582.020 2324.000 3583.180 ;
        RECT 0.560 3580.940 2324.000 3582.020 ;
        RECT 0.860 3579.780 2324.000 3580.940 ;
        RECT 0.560 3578.700 2324.000 3579.780 ;
        RECT 0.860 3577.540 2324.000 3578.700 ;
        RECT 0.560 3576.460 2324.000 3577.540 ;
        RECT 0.860 3575.300 2324.000 3576.460 ;
        RECT 0.560 3574.220 2324.000 3575.300 ;
        RECT 0.860 3573.060 2324.000 3574.220 ;
        RECT 0.560 3571.980 2324.000 3573.060 ;
        RECT 0.860 3570.820 2324.000 3571.980 ;
        RECT 0.560 3569.740 2324.000 3570.820 ;
        RECT 0.860 3568.580 2324.000 3569.740 ;
        RECT 0.560 3567.500 2324.000 3568.580 ;
        RECT 0.860 3566.340 2324.000 3567.500 ;
        RECT 0.560 3565.260 2324.000 3566.340 ;
        RECT 0.860 3564.100 2324.000 3565.260 ;
        RECT 0.560 3563.020 2324.000 3564.100 ;
        RECT 0.860 3561.860 2324.000 3563.020 ;
        RECT 0.560 3560.780 2324.000 3561.860 ;
        RECT 0.860 3559.620 2324.000 3560.780 ;
        RECT 0.560 3558.540 2324.000 3559.620 ;
        RECT 0.860 3557.380 2324.000 3558.540 ;
        RECT 0.560 3556.300 2324.000 3557.380 ;
        RECT 0.860 3555.140 2324.000 3556.300 ;
        RECT 0.560 3554.060 2324.000 3555.140 ;
        RECT 0.860 3552.900 2324.000 3554.060 ;
        RECT 0.560 3551.820 2324.000 3552.900 ;
        RECT 0.860 3550.660 2324.000 3551.820 ;
        RECT 0.560 3549.580 2324.000 3550.660 ;
        RECT 0.860 3548.420 2324.000 3549.580 ;
        RECT 0.560 3547.340 2324.000 3548.420 ;
        RECT 0.860 3546.180 2324.000 3547.340 ;
        RECT 0.560 3545.100 2324.000 3546.180 ;
        RECT 0.860 3543.940 2324.000 3545.100 ;
        RECT 0.560 3542.860 2324.000 3543.940 ;
        RECT 0.860 3541.700 2324.000 3542.860 ;
        RECT 0.560 3540.620 2324.000 3541.700 ;
        RECT 0.860 3539.460 2324.000 3540.620 ;
        RECT 0.560 3538.380 2324.000 3539.460 ;
        RECT 0.860 3537.220 2324.000 3538.380 ;
        RECT 0.560 3536.140 2324.000 3537.220 ;
        RECT 0.860 3534.980 2324.000 3536.140 ;
        RECT 0.560 3533.900 2324.000 3534.980 ;
        RECT 0.860 3532.740 2324.000 3533.900 ;
        RECT 0.560 3531.660 2324.000 3532.740 ;
        RECT 0.860 3530.500 2324.000 3531.660 ;
        RECT 0.560 3529.420 2324.000 3530.500 ;
        RECT 0.860 3528.260 2324.000 3529.420 ;
        RECT 0.560 3527.180 2324.000 3528.260 ;
        RECT 0.860 3526.020 2324.000 3527.180 ;
        RECT 0.560 3524.940 2324.000 3526.020 ;
        RECT 0.860 3523.780 2324.000 3524.940 ;
        RECT 0.560 3513.180 2324.000 3523.780 ;
        RECT 1.420 3512.020 2324.000 3513.180 ;
        RECT 0.560 3508.700 2324.000 3512.020 ;
        RECT 1.420 3507.540 2324.000 3508.700 ;
        RECT 0.560 3504.220 2324.000 3507.540 ;
        RECT 1.420 3503.060 2324.000 3504.220 ;
        RECT 0.560 3499.740 2324.000 3503.060 ;
        RECT 1.420 3498.580 2324.000 3499.740 ;
        RECT 0.560 3495.260 2324.000 3498.580 ;
        RECT 1.420 3494.100 2324.000 3495.260 ;
        RECT 0.560 3490.780 2324.000 3494.100 ;
        RECT 1.420 3489.620 2324.000 3490.780 ;
        RECT 0.560 3486.300 2324.000 3489.620 ;
        RECT 1.420 3485.140 2324.000 3486.300 ;
        RECT 0.560 3481.820 2324.000 3485.140 ;
        RECT 1.420 3480.660 2324.000 3481.820 ;
        RECT 0.560 3477.340 2324.000 3480.660 ;
        RECT 1.420 3476.180 2324.000 3477.340 ;
        RECT 0.560 3472.860 2324.000 3476.180 ;
        RECT 1.420 3471.700 2324.000 3472.860 ;
        RECT 0.560 3468.380 2324.000 3471.700 ;
        RECT 1.420 3467.220 2324.000 3468.380 ;
        RECT 0.560 3463.900 2324.000 3467.220 ;
        RECT 1.420 3462.740 2324.000 3463.900 ;
        RECT 0.560 3459.420 2324.000 3462.740 ;
        RECT 1.420 3458.260 2324.000 3459.420 ;
        RECT 0.560 3454.940 2324.000 3458.260 ;
        RECT 1.420 3453.780 2324.000 3454.940 ;
        RECT 0.560 3450.460 2324.000 3453.780 ;
        RECT 1.420 3449.300 2324.000 3450.460 ;
        RECT 0.560 3445.980 2324.000 3449.300 ;
        RECT 1.420 3444.820 2324.000 3445.980 ;
        RECT 0.560 3441.500 2324.000 3444.820 ;
        RECT 1.420 3440.340 2324.000 3441.500 ;
        RECT 0.560 3437.020 2324.000 3440.340 ;
        RECT 1.420 3435.860 2324.000 3437.020 ;
        RECT 0.560 3432.540 2324.000 3435.860 ;
        RECT 1.420 3431.380 2324.000 3432.540 ;
        RECT 0.560 3428.060 2324.000 3431.380 ;
        RECT 1.420 3426.900 2324.000 3428.060 ;
        RECT 0.560 3423.580 2324.000 3426.900 ;
        RECT 1.420 3422.420 2324.000 3423.580 ;
        RECT 0.560 3419.100 2324.000 3422.420 ;
        RECT 1.420 3417.940 2324.000 3419.100 ;
        RECT 0.560 3414.620 2324.000 3417.940 ;
        RECT 1.420 3413.460 2324.000 3414.620 ;
        RECT 0.560 3410.140 2324.000 3413.460 ;
        RECT 1.420 3408.980 2324.000 3410.140 ;
        RECT 0.560 3405.660 2324.000 3408.980 ;
        RECT 1.420 3404.500 2324.000 3405.660 ;
        RECT 0.560 3401.180 2324.000 3404.500 ;
        RECT 1.420 3400.020 2324.000 3401.180 ;
        RECT 0.560 3396.700 2324.000 3400.020 ;
        RECT 1.420 3395.540 2324.000 3396.700 ;
        RECT 0.560 3392.220 2324.000 3395.540 ;
        RECT 1.420 3391.060 2324.000 3392.220 ;
        RECT 0.560 3387.740 2324.000 3391.060 ;
        RECT 1.420 3386.580 2324.000 3387.740 ;
        RECT 0.560 3383.260 2324.000 3386.580 ;
        RECT 1.420 3382.100 2324.000 3383.260 ;
        RECT 0.560 3378.780 2324.000 3382.100 ;
        RECT 1.420 3377.620 2324.000 3378.780 ;
        RECT 0.560 3374.300 2324.000 3377.620 ;
        RECT 1.420 3373.140 2324.000 3374.300 ;
        RECT 0.560 3369.820 2324.000 3373.140 ;
        RECT 1.420 3368.660 2324.000 3369.820 ;
        RECT 0.560 3365.340 2324.000 3368.660 ;
        RECT 1.420 3364.180 2324.000 3365.340 ;
        RECT 0.560 3360.860 2324.000 3364.180 ;
        RECT 1.420 3359.700 2324.000 3360.860 ;
        RECT 0.560 3356.380 2324.000 3359.700 ;
        RECT 1.420 3355.220 2324.000 3356.380 ;
        RECT 0.560 3351.900 2324.000 3355.220 ;
        RECT 1.420 3350.740 2324.000 3351.900 ;
        RECT 0.560 3347.420 2324.000 3350.740 ;
        RECT 1.420 3346.260 2324.000 3347.420 ;
        RECT 0.560 3342.940 2324.000 3346.260 ;
        RECT 1.420 3341.780 2324.000 3342.940 ;
        RECT 0.560 3338.460 2324.000 3341.780 ;
        RECT 1.420 3337.300 2324.000 3338.460 ;
        RECT 0.560 3333.980 2324.000 3337.300 ;
        RECT 1.420 3332.820 2324.000 3333.980 ;
        RECT 0.560 3329.500 2324.000 3332.820 ;
        RECT 1.420 3328.340 2324.000 3329.500 ;
        RECT 0.560 3325.020 2324.000 3328.340 ;
        RECT 1.420 3323.860 2324.000 3325.020 ;
        RECT 0.560 3320.540 2324.000 3323.860 ;
        RECT 1.420 3319.380 2324.000 3320.540 ;
        RECT 0.560 3316.060 2324.000 3319.380 ;
        RECT 1.420 3314.900 2324.000 3316.060 ;
        RECT 0.560 3311.580 2324.000 3314.900 ;
        RECT 1.420 3310.420 2324.000 3311.580 ;
        RECT 0.560 3307.100 2324.000 3310.420 ;
        RECT 1.420 3305.940 2324.000 3307.100 ;
        RECT 0.560 3302.620 2324.000 3305.940 ;
        RECT 1.420 3301.460 2324.000 3302.620 ;
        RECT 0.560 3298.140 2324.000 3301.460 ;
        RECT 1.420 3296.980 2324.000 3298.140 ;
        RECT 0.560 3293.660 2324.000 3296.980 ;
        RECT 1.420 3292.500 2324.000 3293.660 ;
        RECT 0.560 3289.180 2324.000 3292.500 ;
        RECT 1.420 3288.020 2324.000 3289.180 ;
        RECT 0.560 3284.700 2324.000 3288.020 ;
        RECT 1.420 3283.540 2324.000 3284.700 ;
        RECT 0.560 3280.220 2324.000 3283.540 ;
        RECT 1.420 3279.060 2324.000 3280.220 ;
        RECT 0.560 3275.740 2324.000 3279.060 ;
        RECT 1.420 3274.580 2324.000 3275.740 ;
        RECT 0.560 3271.260 2324.000 3274.580 ;
        RECT 1.420 3270.100 2324.000 3271.260 ;
        RECT 0.560 3266.780 2324.000 3270.100 ;
        RECT 1.420 3265.620 2324.000 3266.780 ;
        RECT 0.560 3262.300 2324.000 3265.620 ;
        RECT 1.420 3261.140 2324.000 3262.300 ;
        RECT 0.560 3257.820 2324.000 3261.140 ;
        RECT 1.420 3256.660 2324.000 3257.820 ;
        RECT 0.560 3253.340 2324.000 3256.660 ;
        RECT 1.420 3252.180 2324.000 3253.340 ;
        RECT 0.560 3248.860 2324.000 3252.180 ;
        RECT 1.420 3247.700 2324.000 3248.860 ;
        RECT 0.560 3225.900 2324.000 3247.700 ;
        RECT 1.420 3224.740 2324.000 3225.900 ;
        RECT 0.560 3221.420 2324.000 3224.740 ;
        RECT 1.420 3220.260 2324.000 3221.420 ;
        RECT 0.560 3216.940 2324.000 3220.260 ;
        RECT 1.420 3215.780 2324.000 3216.940 ;
        RECT 0.560 3212.460 2324.000 3215.780 ;
        RECT 1.420 3211.300 2324.000 3212.460 ;
        RECT 0.560 3207.980 2324.000 3211.300 ;
        RECT 1.420 3206.820 2324.000 3207.980 ;
        RECT 0.560 3203.500 2324.000 3206.820 ;
        RECT 1.420 3202.340 2324.000 3203.500 ;
        RECT 0.560 3199.020 2324.000 3202.340 ;
        RECT 1.420 3197.860 2324.000 3199.020 ;
        RECT 0.560 3194.540 2324.000 3197.860 ;
        RECT 1.420 3193.380 2324.000 3194.540 ;
        RECT 0.560 3190.060 2324.000 3193.380 ;
        RECT 1.420 3188.900 2324.000 3190.060 ;
        RECT 0.560 3185.580 2324.000 3188.900 ;
        RECT 1.420 3184.420 2324.000 3185.580 ;
        RECT 0.560 3181.100 2324.000 3184.420 ;
        RECT 1.420 3179.940 2324.000 3181.100 ;
        RECT 0.560 3176.620 2324.000 3179.940 ;
        RECT 1.420 3175.460 2324.000 3176.620 ;
        RECT 0.560 3172.140 2324.000 3175.460 ;
        RECT 1.420 3170.980 2324.000 3172.140 ;
        RECT 0.560 3167.660 2324.000 3170.980 ;
        RECT 1.420 3166.500 2324.000 3167.660 ;
        RECT 0.560 3163.180 2324.000 3166.500 ;
        RECT 1.420 3162.020 2324.000 3163.180 ;
        RECT 0.560 3158.700 2324.000 3162.020 ;
        RECT 1.420 3157.540 2324.000 3158.700 ;
        RECT 0.560 3154.220 2324.000 3157.540 ;
        RECT 1.420 3153.060 2324.000 3154.220 ;
        RECT 0.560 3149.740 2324.000 3153.060 ;
        RECT 1.420 3148.580 2324.000 3149.740 ;
        RECT 0.560 3145.260 2324.000 3148.580 ;
        RECT 1.420 3144.100 2324.000 3145.260 ;
        RECT 0.560 3140.780 2324.000 3144.100 ;
        RECT 1.420 3139.620 2324.000 3140.780 ;
        RECT 0.560 3136.300 2324.000 3139.620 ;
        RECT 1.420 3135.140 2324.000 3136.300 ;
        RECT 0.560 3131.820 2324.000 3135.140 ;
        RECT 1.420 3130.660 2324.000 3131.820 ;
        RECT 0.560 3127.340 2324.000 3130.660 ;
        RECT 1.420 3126.220 2324.000 3127.340 ;
        RECT 1.420 3126.180 2323.140 3126.220 ;
        RECT 0.560 3125.060 2323.140 3126.180 ;
        RECT 0.560 3122.860 2324.000 3125.060 ;
        RECT 1.420 3121.740 2324.000 3122.860 ;
        RECT 1.420 3121.700 2323.140 3121.740 ;
        RECT 0.560 3120.580 2323.140 3121.700 ;
        RECT 0.560 3118.380 2324.000 3120.580 ;
        RECT 1.420 3117.260 2324.000 3118.380 ;
        RECT 1.420 3117.220 2323.140 3117.260 ;
        RECT 0.560 3116.100 2323.140 3117.220 ;
        RECT 0.560 3113.900 2324.000 3116.100 ;
        RECT 1.420 3112.780 2324.000 3113.900 ;
        RECT 1.420 3112.740 2323.140 3112.780 ;
        RECT 0.560 3111.620 2323.140 3112.740 ;
        RECT 0.560 3109.420 2324.000 3111.620 ;
        RECT 1.420 3108.300 2324.000 3109.420 ;
        RECT 1.420 3108.260 2323.140 3108.300 ;
        RECT 0.560 3107.140 2323.140 3108.260 ;
        RECT 0.560 3104.940 2324.000 3107.140 ;
        RECT 1.420 3103.820 2324.000 3104.940 ;
        RECT 1.420 3103.780 2323.140 3103.820 ;
        RECT 0.560 3102.660 2323.140 3103.780 ;
        RECT 0.560 3100.460 2324.000 3102.660 ;
        RECT 1.420 3099.340 2324.000 3100.460 ;
        RECT 1.420 3099.300 2323.140 3099.340 ;
        RECT 0.560 3098.180 2323.140 3099.300 ;
        RECT 0.560 3095.980 2324.000 3098.180 ;
        RECT 1.420 3094.860 2324.000 3095.980 ;
        RECT 1.420 3094.820 2323.140 3094.860 ;
        RECT 0.560 3093.700 2323.140 3094.820 ;
        RECT 0.560 3091.500 2324.000 3093.700 ;
        RECT 1.420 3090.380 2324.000 3091.500 ;
        RECT 1.420 3090.340 2323.140 3090.380 ;
        RECT 0.560 3089.220 2323.140 3090.340 ;
        RECT 0.560 3087.020 2324.000 3089.220 ;
        RECT 1.420 3085.900 2324.000 3087.020 ;
        RECT 1.420 3085.860 2323.140 3085.900 ;
        RECT 0.560 3084.740 2323.140 3085.860 ;
        RECT 0.560 3082.540 2324.000 3084.740 ;
        RECT 1.420 3081.420 2324.000 3082.540 ;
        RECT 1.420 3081.380 2323.140 3081.420 ;
        RECT 0.560 3080.260 2323.140 3081.380 ;
        RECT 0.560 3078.060 2324.000 3080.260 ;
        RECT 1.420 3076.940 2324.000 3078.060 ;
        RECT 1.420 3076.900 2323.140 3076.940 ;
        RECT 0.560 3075.780 2323.140 3076.900 ;
        RECT 0.560 3073.580 2324.000 3075.780 ;
        RECT 1.420 3072.460 2324.000 3073.580 ;
        RECT 1.420 3072.420 2323.140 3072.460 ;
        RECT 0.560 3071.300 2323.140 3072.420 ;
        RECT 0.560 3069.100 2324.000 3071.300 ;
        RECT 1.420 3067.980 2324.000 3069.100 ;
        RECT 1.420 3067.940 2323.140 3067.980 ;
        RECT 0.560 3066.820 2323.140 3067.940 ;
        RECT 0.560 3064.620 2324.000 3066.820 ;
        RECT 1.420 3063.500 2324.000 3064.620 ;
        RECT 1.420 3063.460 2323.140 3063.500 ;
        RECT 0.560 3062.340 2323.140 3063.460 ;
        RECT 0.560 3060.140 2324.000 3062.340 ;
        RECT 1.420 3059.020 2324.000 3060.140 ;
        RECT 1.420 3058.980 2323.140 3059.020 ;
        RECT 0.560 3057.860 2323.140 3058.980 ;
        RECT 0.560 3055.660 2324.000 3057.860 ;
        RECT 1.420 3054.540 2324.000 3055.660 ;
        RECT 1.420 3054.500 2323.140 3054.540 ;
        RECT 0.560 3053.380 2323.140 3054.500 ;
        RECT 0.560 3051.180 2324.000 3053.380 ;
        RECT 1.420 3050.060 2324.000 3051.180 ;
        RECT 1.420 3050.020 2323.140 3050.060 ;
        RECT 0.560 3048.900 2323.140 3050.020 ;
        RECT 0.560 3046.700 2324.000 3048.900 ;
        RECT 1.420 3045.580 2324.000 3046.700 ;
        RECT 1.420 3045.540 2323.140 3045.580 ;
        RECT 0.560 3044.420 2323.140 3045.540 ;
        RECT 0.560 3042.220 2324.000 3044.420 ;
        RECT 1.420 3041.100 2324.000 3042.220 ;
        RECT 1.420 3041.060 2323.140 3041.100 ;
        RECT 0.560 3039.940 2323.140 3041.060 ;
        RECT 0.560 3037.740 2324.000 3039.940 ;
        RECT 1.420 3036.620 2324.000 3037.740 ;
        RECT 1.420 3036.580 2323.140 3036.620 ;
        RECT 0.560 3035.460 2323.140 3036.580 ;
        RECT 0.560 3033.260 2324.000 3035.460 ;
        RECT 1.420 3032.140 2324.000 3033.260 ;
        RECT 1.420 3032.100 2323.140 3032.140 ;
        RECT 0.560 3030.980 2323.140 3032.100 ;
        RECT 0.560 3028.780 2324.000 3030.980 ;
        RECT 1.420 3027.660 2324.000 3028.780 ;
        RECT 1.420 3027.620 2323.140 3027.660 ;
        RECT 0.560 3026.500 2323.140 3027.620 ;
        RECT 0.560 3024.300 2324.000 3026.500 ;
        RECT 1.420 3023.180 2324.000 3024.300 ;
        RECT 1.420 3023.140 2323.140 3023.180 ;
        RECT 0.560 3022.020 2323.140 3023.140 ;
        RECT 0.560 3019.820 2324.000 3022.020 ;
        RECT 1.420 3018.700 2324.000 3019.820 ;
        RECT 1.420 3018.660 2323.140 3018.700 ;
        RECT 0.560 3017.540 2323.140 3018.660 ;
        RECT 0.560 3015.340 2324.000 3017.540 ;
        RECT 1.420 3014.220 2324.000 3015.340 ;
        RECT 1.420 3014.180 2323.140 3014.220 ;
        RECT 0.560 3013.060 2323.140 3014.180 ;
        RECT 0.560 3010.860 2324.000 3013.060 ;
        RECT 1.420 3009.740 2324.000 3010.860 ;
        RECT 1.420 3009.700 2323.140 3009.740 ;
        RECT 0.560 3008.580 2323.140 3009.700 ;
        RECT 0.560 3006.380 2324.000 3008.580 ;
        RECT 1.420 3005.260 2324.000 3006.380 ;
        RECT 1.420 3005.220 2323.140 3005.260 ;
        RECT 0.560 3004.100 2323.140 3005.220 ;
        RECT 0.560 3001.900 2324.000 3004.100 ;
        RECT 1.420 3000.780 2324.000 3001.900 ;
        RECT 1.420 3000.740 2323.140 3000.780 ;
        RECT 0.560 2999.620 2323.140 3000.740 ;
        RECT 0.560 2997.420 2324.000 2999.620 ;
        RECT 1.420 2996.300 2324.000 2997.420 ;
        RECT 1.420 2996.260 2323.140 2996.300 ;
        RECT 0.560 2995.140 2323.140 2996.260 ;
        RECT 0.560 2992.940 2324.000 2995.140 ;
        RECT 1.420 2991.820 2324.000 2992.940 ;
        RECT 1.420 2991.780 2323.140 2991.820 ;
        RECT 0.560 2990.660 2323.140 2991.780 ;
        RECT 0.560 2988.460 2324.000 2990.660 ;
        RECT 1.420 2987.340 2324.000 2988.460 ;
        RECT 1.420 2987.300 2323.140 2987.340 ;
        RECT 0.560 2986.180 2323.140 2987.300 ;
        RECT 0.560 2983.980 2324.000 2986.180 ;
        RECT 1.420 2982.860 2324.000 2983.980 ;
        RECT 1.420 2982.820 2323.140 2982.860 ;
        RECT 0.560 2981.700 2323.140 2982.820 ;
        RECT 0.560 2979.500 2324.000 2981.700 ;
        RECT 1.420 2978.380 2324.000 2979.500 ;
        RECT 1.420 2978.340 2323.140 2978.380 ;
        RECT 0.560 2977.220 2323.140 2978.340 ;
        RECT 0.560 2975.020 2324.000 2977.220 ;
        RECT 1.420 2973.900 2324.000 2975.020 ;
        RECT 1.420 2973.860 2323.140 2973.900 ;
        RECT 0.560 2972.740 2323.140 2973.860 ;
        RECT 0.560 2970.540 2324.000 2972.740 ;
        RECT 1.420 2969.420 2324.000 2970.540 ;
        RECT 1.420 2969.380 2323.140 2969.420 ;
        RECT 0.560 2968.260 2323.140 2969.380 ;
        RECT 0.560 2966.060 2324.000 2968.260 ;
        RECT 1.420 2964.940 2324.000 2966.060 ;
        RECT 1.420 2964.900 2323.140 2964.940 ;
        RECT 0.560 2963.780 2323.140 2964.900 ;
        RECT 0.560 2961.580 2324.000 2963.780 ;
        RECT 1.420 2960.420 2324.000 2961.580 ;
        RECT 0.560 2938.620 2324.000 2960.420 ;
        RECT 1.420 2937.460 2324.000 2938.620 ;
        RECT 0.560 2934.140 2324.000 2937.460 ;
        RECT 1.420 2932.980 2324.000 2934.140 ;
        RECT 0.560 2929.660 2324.000 2932.980 ;
        RECT 1.420 2928.500 2324.000 2929.660 ;
        RECT 0.560 2925.180 2324.000 2928.500 ;
        RECT 1.420 2924.020 2324.000 2925.180 ;
        RECT 0.560 2920.700 2324.000 2924.020 ;
        RECT 1.420 2919.540 2324.000 2920.700 ;
        RECT 0.560 2916.220 2324.000 2919.540 ;
        RECT 1.420 2915.060 2324.000 2916.220 ;
        RECT 0.560 2911.740 2324.000 2915.060 ;
        RECT 1.420 2910.580 2324.000 2911.740 ;
        RECT 0.560 2907.260 2324.000 2910.580 ;
        RECT 1.420 2906.100 2324.000 2907.260 ;
        RECT 0.560 2902.780 2324.000 2906.100 ;
        RECT 1.420 2901.620 2324.000 2902.780 ;
        RECT 0.560 2898.300 2324.000 2901.620 ;
        RECT 1.420 2897.140 2324.000 2898.300 ;
        RECT 0.560 2893.820 2324.000 2897.140 ;
        RECT 1.420 2892.660 2324.000 2893.820 ;
        RECT 0.560 2889.340 2324.000 2892.660 ;
        RECT 1.420 2888.180 2324.000 2889.340 ;
        RECT 0.560 2884.860 2324.000 2888.180 ;
        RECT 1.420 2883.700 2324.000 2884.860 ;
        RECT 0.560 2880.380 2324.000 2883.700 ;
        RECT 1.420 2879.220 2324.000 2880.380 ;
        RECT 0.560 2875.900 2324.000 2879.220 ;
        RECT 1.420 2874.740 2324.000 2875.900 ;
        RECT 0.560 2871.420 2324.000 2874.740 ;
        RECT 1.420 2870.260 2324.000 2871.420 ;
        RECT 0.560 2866.940 2324.000 2870.260 ;
        RECT 1.420 2865.780 2324.000 2866.940 ;
        RECT 0.560 2862.460 2324.000 2865.780 ;
        RECT 1.420 2861.300 2324.000 2862.460 ;
        RECT 0.560 2857.980 2324.000 2861.300 ;
        RECT 1.420 2856.820 2324.000 2857.980 ;
        RECT 0.560 2853.500 2324.000 2856.820 ;
        RECT 1.420 2852.340 2324.000 2853.500 ;
        RECT 0.560 2849.020 2324.000 2852.340 ;
        RECT 1.420 2847.860 2324.000 2849.020 ;
        RECT 0.560 2844.540 2324.000 2847.860 ;
        RECT 1.420 2843.380 2324.000 2844.540 ;
        RECT 0.560 2840.060 2324.000 2843.380 ;
        RECT 1.420 2838.900 2324.000 2840.060 ;
        RECT 0.560 2835.580 2324.000 2838.900 ;
        RECT 1.420 2834.420 2324.000 2835.580 ;
        RECT 0.560 2831.100 2324.000 2834.420 ;
        RECT 1.420 2829.940 2324.000 2831.100 ;
        RECT 0.560 2826.620 2324.000 2829.940 ;
        RECT 1.420 2825.460 2324.000 2826.620 ;
        RECT 0.560 2822.140 2324.000 2825.460 ;
        RECT 1.420 2820.980 2324.000 2822.140 ;
        RECT 0.560 2817.660 2324.000 2820.980 ;
        RECT 1.420 2816.500 2324.000 2817.660 ;
        RECT 0.560 2813.180 2324.000 2816.500 ;
        RECT 1.420 2812.020 2324.000 2813.180 ;
        RECT 0.560 2808.700 2324.000 2812.020 ;
        RECT 1.420 2807.540 2324.000 2808.700 ;
        RECT 0.560 2804.220 2324.000 2807.540 ;
        RECT 1.420 2803.060 2324.000 2804.220 ;
        RECT 0.560 2799.740 2324.000 2803.060 ;
        RECT 1.420 2798.580 2324.000 2799.740 ;
        RECT 0.560 2795.260 2324.000 2798.580 ;
        RECT 1.420 2794.100 2324.000 2795.260 ;
        RECT 0.560 2790.780 2324.000 2794.100 ;
        RECT 1.420 2789.620 2324.000 2790.780 ;
        RECT 0.560 2786.300 2324.000 2789.620 ;
        RECT 1.420 2785.140 2324.000 2786.300 ;
        RECT 0.560 2781.820 2324.000 2785.140 ;
        RECT 1.420 2780.660 2324.000 2781.820 ;
        RECT 0.560 2777.340 2324.000 2780.660 ;
        RECT 1.420 2776.180 2324.000 2777.340 ;
        RECT 0.560 2772.860 2324.000 2776.180 ;
        RECT 1.420 2771.700 2324.000 2772.860 ;
        RECT 0.560 2768.380 2324.000 2771.700 ;
        RECT 1.420 2767.220 2324.000 2768.380 ;
        RECT 0.560 2763.900 2324.000 2767.220 ;
        RECT 1.420 2762.740 2324.000 2763.900 ;
        RECT 0.560 2759.420 2324.000 2762.740 ;
        RECT 1.420 2758.260 2324.000 2759.420 ;
        RECT 0.560 2754.940 2324.000 2758.260 ;
        RECT 1.420 2753.780 2324.000 2754.940 ;
        RECT 0.560 2750.460 2324.000 2753.780 ;
        RECT 1.420 2749.300 2324.000 2750.460 ;
        RECT 0.560 2745.980 2324.000 2749.300 ;
        RECT 1.420 2744.820 2324.000 2745.980 ;
        RECT 0.560 2741.500 2324.000 2744.820 ;
        RECT 1.420 2740.340 2324.000 2741.500 ;
        RECT 0.560 2737.020 2324.000 2740.340 ;
        RECT 1.420 2735.860 2324.000 2737.020 ;
        RECT 0.560 2732.540 2324.000 2735.860 ;
        RECT 1.420 2731.380 2324.000 2732.540 ;
        RECT 0.560 2728.060 2324.000 2731.380 ;
        RECT 1.420 2726.900 2324.000 2728.060 ;
        RECT 0.560 2723.580 2324.000 2726.900 ;
        RECT 1.420 2722.420 2324.000 2723.580 ;
        RECT 0.560 2719.100 2324.000 2722.420 ;
        RECT 1.420 2717.940 2324.000 2719.100 ;
        RECT 0.560 2714.620 2324.000 2717.940 ;
        RECT 1.420 2713.460 2324.000 2714.620 ;
        RECT 0.560 2710.140 2324.000 2713.460 ;
        RECT 1.420 2708.980 2324.000 2710.140 ;
        RECT 0.560 2705.660 2324.000 2708.980 ;
        RECT 1.420 2704.500 2324.000 2705.660 ;
        RECT 0.560 2701.180 2324.000 2704.500 ;
        RECT 1.420 2700.020 2324.000 2701.180 ;
        RECT 0.560 2696.700 2324.000 2700.020 ;
        RECT 1.420 2695.540 2324.000 2696.700 ;
        RECT 0.560 2692.220 2324.000 2695.540 ;
        RECT 1.420 2691.060 2324.000 2692.220 ;
        RECT 0.560 2687.740 2324.000 2691.060 ;
        RECT 1.420 2686.580 2324.000 2687.740 ;
        RECT 0.560 2683.260 2324.000 2686.580 ;
        RECT 1.420 2682.100 2324.000 2683.260 ;
        RECT 0.560 2678.780 2324.000 2682.100 ;
        RECT 1.420 2677.620 2324.000 2678.780 ;
        RECT 0.560 2674.300 2324.000 2677.620 ;
        RECT 1.420 2673.140 2324.000 2674.300 ;
        RECT 0.560 2651.340 2324.000 2673.140 ;
        RECT 1.420 2650.180 2324.000 2651.340 ;
        RECT 0.560 2646.860 2324.000 2650.180 ;
        RECT 1.420 2645.700 2324.000 2646.860 ;
        RECT 0.560 2642.380 2324.000 2645.700 ;
        RECT 1.420 2641.220 2324.000 2642.380 ;
        RECT 0.560 2637.900 2324.000 2641.220 ;
        RECT 1.420 2636.740 2324.000 2637.900 ;
        RECT 0.560 2633.420 2324.000 2636.740 ;
        RECT 1.420 2632.260 2324.000 2633.420 ;
        RECT 0.560 2628.940 2324.000 2632.260 ;
        RECT 1.420 2627.780 2324.000 2628.940 ;
        RECT 0.560 2624.460 2324.000 2627.780 ;
        RECT 1.420 2623.300 2324.000 2624.460 ;
        RECT 0.560 2619.980 2324.000 2623.300 ;
        RECT 1.420 2618.820 2324.000 2619.980 ;
        RECT 0.560 2615.500 2324.000 2618.820 ;
        RECT 1.420 2614.340 2324.000 2615.500 ;
        RECT 0.560 2611.020 2324.000 2614.340 ;
        RECT 1.420 2609.860 2324.000 2611.020 ;
        RECT 0.560 2606.540 2324.000 2609.860 ;
        RECT 1.420 2605.380 2324.000 2606.540 ;
        RECT 0.560 2602.060 2324.000 2605.380 ;
        RECT 1.420 2600.900 2324.000 2602.060 ;
        RECT 0.560 2597.580 2324.000 2600.900 ;
        RECT 1.420 2596.420 2324.000 2597.580 ;
        RECT 0.560 2593.100 2324.000 2596.420 ;
        RECT 1.420 2591.940 2324.000 2593.100 ;
        RECT 0.560 2588.620 2324.000 2591.940 ;
        RECT 1.420 2587.460 2324.000 2588.620 ;
        RECT 0.560 2584.140 2324.000 2587.460 ;
        RECT 1.420 2582.980 2324.000 2584.140 ;
        RECT 0.560 2579.660 2324.000 2582.980 ;
        RECT 1.420 2578.500 2324.000 2579.660 ;
        RECT 0.560 2575.180 2324.000 2578.500 ;
        RECT 1.420 2574.020 2324.000 2575.180 ;
        RECT 0.560 2570.700 2324.000 2574.020 ;
        RECT 1.420 2569.540 2324.000 2570.700 ;
        RECT 0.560 2566.220 2324.000 2569.540 ;
        RECT 1.420 2565.060 2324.000 2566.220 ;
        RECT 0.560 2561.740 2324.000 2565.060 ;
        RECT 1.420 2560.580 2324.000 2561.740 ;
        RECT 0.560 2557.260 2324.000 2560.580 ;
        RECT 1.420 2556.100 2324.000 2557.260 ;
        RECT 0.560 2552.780 2324.000 2556.100 ;
        RECT 1.420 2551.660 2324.000 2552.780 ;
        RECT 1.420 2551.620 2323.140 2551.660 ;
        RECT 0.560 2550.500 2323.140 2551.620 ;
        RECT 0.560 2548.300 2324.000 2550.500 ;
        RECT 1.420 2547.180 2324.000 2548.300 ;
        RECT 1.420 2547.140 2323.140 2547.180 ;
        RECT 0.560 2546.020 2323.140 2547.140 ;
        RECT 0.560 2543.820 2324.000 2546.020 ;
        RECT 1.420 2542.700 2324.000 2543.820 ;
        RECT 1.420 2542.660 2323.140 2542.700 ;
        RECT 0.560 2541.540 2323.140 2542.660 ;
        RECT 0.560 2539.340 2324.000 2541.540 ;
        RECT 1.420 2538.220 2324.000 2539.340 ;
        RECT 1.420 2538.180 2323.140 2538.220 ;
        RECT 0.560 2537.060 2323.140 2538.180 ;
        RECT 0.560 2534.860 2324.000 2537.060 ;
        RECT 1.420 2533.740 2324.000 2534.860 ;
        RECT 1.420 2533.700 2323.140 2533.740 ;
        RECT 0.560 2532.580 2323.140 2533.700 ;
        RECT 0.560 2530.380 2324.000 2532.580 ;
        RECT 1.420 2529.260 2324.000 2530.380 ;
        RECT 1.420 2529.220 2323.140 2529.260 ;
        RECT 0.560 2528.100 2323.140 2529.220 ;
        RECT 0.560 2525.900 2324.000 2528.100 ;
        RECT 1.420 2524.780 2324.000 2525.900 ;
        RECT 1.420 2524.740 2323.140 2524.780 ;
        RECT 0.560 2523.620 2323.140 2524.740 ;
        RECT 0.560 2521.420 2324.000 2523.620 ;
        RECT 1.420 2520.300 2324.000 2521.420 ;
        RECT 1.420 2520.260 2323.140 2520.300 ;
        RECT 0.560 2519.140 2323.140 2520.260 ;
        RECT 0.560 2516.940 2324.000 2519.140 ;
        RECT 1.420 2515.820 2324.000 2516.940 ;
        RECT 1.420 2515.780 2323.140 2515.820 ;
        RECT 0.560 2514.660 2323.140 2515.780 ;
        RECT 0.560 2512.460 2324.000 2514.660 ;
        RECT 1.420 2511.340 2324.000 2512.460 ;
        RECT 1.420 2511.300 2323.140 2511.340 ;
        RECT 0.560 2510.180 2323.140 2511.300 ;
        RECT 0.560 2507.980 2324.000 2510.180 ;
        RECT 1.420 2506.860 2324.000 2507.980 ;
        RECT 1.420 2506.820 2323.140 2506.860 ;
        RECT 0.560 2505.700 2323.140 2506.820 ;
        RECT 0.560 2503.500 2324.000 2505.700 ;
        RECT 1.420 2502.380 2324.000 2503.500 ;
        RECT 1.420 2502.340 2323.140 2502.380 ;
        RECT 0.560 2501.220 2323.140 2502.340 ;
        RECT 0.560 2499.020 2324.000 2501.220 ;
        RECT 1.420 2497.900 2324.000 2499.020 ;
        RECT 1.420 2497.860 2323.140 2497.900 ;
        RECT 0.560 2496.740 2323.140 2497.860 ;
        RECT 0.560 2494.540 2324.000 2496.740 ;
        RECT 1.420 2493.420 2324.000 2494.540 ;
        RECT 1.420 2493.380 2323.140 2493.420 ;
        RECT 0.560 2492.260 2323.140 2493.380 ;
        RECT 0.560 2490.060 2324.000 2492.260 ;
        RECT 1.420 2488.940 2324.000 2490.060 ;
        RECT 1.420 2488.900 2323.140 2488.940 ;
        RECT 0.560 2487.780 2323.140 2488.900 ;
        RECT 0.560 2485.580 2324.000 2487.780 ;
        RECT 1.420 2484.460 2324.000 2485.580 ;
        RECT 1.420 2484.420 2323.140 2484.460 ;
        RECT 0.560 2483.300 2323.140 2484.420 ;
        RECT 0.560 2481.100 2324.000 2483.300 ;
        RECT 1.420 2479.980 2324.000 2481.100 ;
        RECT 1.420 2479.940 2323.140 2479.980 ;
        RECT 0.560 2478.820 2323.140 2479.940 ;
        RECT 0.560 2476.620 2324.000 2478.820 ;
        RECT 1.420 2475.500 2324.000 2476.620 ;
        RECT 1.420 2475.460 2323.140 2475.500 ;
        RECT 0.560 2474.340 2323.140 2475.460 ;
        RECT 0.560 2472.140 2324.000 2474.340 ;
        RECT 1.420 2471.020 2324.000 2472.140 ;
        RECT 1.420 2470.980 2323.140 2471.020 ;
        RECT 0.560 2469.860 2323.140 2470.980 ;
        RECT 0.560 2467.660 2324.000 2469.860 ;
        RECT 1.420 2466.540 2324.000 2467.660 ;
        RECT 1.420 2466.500 2323.140 2466.540 ;
        RECT 0.560 2465.380 2323.140 2466.500 ;
        RECT 0.560 2463.180 2324.000 2465.380 ;
        RECT 1.420 2462.060 2324.000 2463.180 ;
        RECT 1.420 2462.020 2323.140 2462.060 ;
        RECT 0.560 2460.900 2323.140 2462.020 ;
        RECT 0.560 2458.700 2324.000 2460.900 ;
        RECT 1.420 2457.580 2324.000 2458.700 ;
        RECT 1.420 2457.540 2323.140 2457.580 ;
        RECT 0.560 2456.420 2323.140 2457.540 ;
        RECT 0.560 2454.220 2324.000 2456.420 ;
        RECT 1.420 2453.100 2324.000 2454.220 ;
        RECT 1.420 2453.060 2323.140 2453.100 ;
        RECT 0.560 2451.940 2323.140 2453.060 ;
        RECT 0.560 2449.740 2324.000 2451.940 ;
        RECT 1.420 2448.620 2324.000 2449.740 ;
        RECT 1.420 2448.580 2323.140 2448.620 ;
        RECT 0.560 2447.460 2323.140 2448.580 ;
        RECT 0.560 2445.260 2324.000 2447.460 ;
        RECT 1.420 2444.140 2324.000 2445.260 ;
        RECT 1.420 2444.100 2323.140 2444.140 ;
        RECT 0.560 2442.980 2323.140 2444.100 ;
        RECT 0.560 2440.780 2324.000 2442.980 ;
        RECT 1.420 2439.660 2324.000 2440.780 ;
        RECT 1.420 2439.620 2323.140 2439.660 ;
        RECT 0.560 2438.500 2323.140 2439.620 ;
        RECT 0.560 2436.300 2324.000 2438.500 ;
        RECT 1.420 2435.180 2324.000 2436.300 ;
        RECT 1.420 2435.140 2323.140 2435.180 ;
        RECT 0.560 2434.020 2323.140 2435.140 ;
        RECT 0.560 2431.820 2324.000 2434.020 ;
        RECT 1.420 2430.700 2324.000 2431.820 ;
        RECT 1.420 2430.660 2323.140 2430.700 ;
        RECT 0.560 2429.540 2323.140 2430.660 ;
        RECT 0.560 2427.340 2324.000 2429.540 ;
        RECT 1.420 2426.220 2324.000 2427.340 ;
        RECT 1.420 2426.180 2323.140 2426.220 ;
        RECT 0.560 2425.060 2323.140 2426.180 ;
        RECT 0.560 2422.860 2324.000 2425.060 ;
        RECT 1.420 2421.740 2324.000 2422.860 ;
        RECT 1.420 2421.700 2323.140 2421.740 ;
        RECT 0.560 2420.580 2323.140 2421.700 ;
        RECT 0.560 2418.380 2324.000 2420.580 ;
        RECT 1.420 2417.260 2324.000 2418.380 ;
        RECT 1.420 2417.220 2323.140 2417.260 ;
        RECT 0.560 2416.100 2323.140 2417.220 ;
        RECT 0.560 2413.900 2324.000 2416.100 ;
        RECT 1.420 2412.780 2324.000 2413.900 ;
        RECT 1.420 2412.740 2323.140 2412.780 ;
        RECT 0.560 2411.620 2323.140 2412.740 ;
        RECT 0.560 2409.420 2324.000 2411.620 ;
        RECT 1.420 2408.300 2324.000 2409.420 ;
        RECT 1.420 2408.260 2323.140 2408.300 ;
        RECT 0.560 2407.140 2323.140 2408.260 ;
        RECT 0.560 2404.940 2324.000 2407.140 ;
        RECT 1.420 2403.820 2324.000 2404.940 ;
        RECT 1.420 2403.780 2323.140 2403.820 ;
        RECT 0.560 2402.660 2323.140 2403.780 ;
        RECT 0.560 2400.460 2324.000 2402.660 ;
        RECT 1.420 2399.340 2324.000 2400.460 ;
        RECT 1.420 2399.300 2323.140 2399.340 ;
        RECT 0.560 2398.180 2323.140 2399.300 ;
        RECT 0.560 2395.980 2324.000 2398.180 ;
        RECT 1.420 2394.860 2324.000 2395.980 ;
        RECT 1.420 2394.820 2323.140 2394.860 ;
        RECT 0.560 2393.700 2323.140 2394.820 ;
        RECT 0.560 2391.500 2324.000 2393.700 ;
        RECT 1.420 2390.380 2324.000 2391.500 ;
        RECT 1.420 2390.340 2323.140 2390.380 ;
        RECT 0.560 2389.220 2323.140 2390.340 ;
        RECT 0.560 2387.020 2324.000 2389.220 ;
        RECT 1.420 2385.860 2324.000 2387.020 ;
        RECT 0.560 2364.060 2324.000 2385.860 ;
        RECT 1.420 2362.900 2324.000 2364.060 ;
        RECT 0.560 2359.580 2324.000 2362.900 ;
        RECT 1.420 2358.420 2324.000 2359.580 ;
        RECT 0.560 2355.100 2324.000 2358.420 ;
        RECT 1.420 2353.940 2324.000 2355.100 ;
        RECT 0.560 2350.620 2324.000 2353.940 ;
        RECT 1.420 2349.460 2324.000 2350.620 ;
        RECT 0.560 2346.140 2324.000 2349.460 ;
        RECT 1.420 2344.980 2324.000 2346.140 ;
        RECT 0.560 2341.660 2324.000 2344.980 ;
        RECT 1.420 2340.500 2324.000 2341.660 ;
        RECT 0.560 2337.180 2324.000 2340.500 ;
        RECT 1.420 2336.020 2324.000 2337.180 ;
        RECT 0.560 2332.700 2324.000 2336.020 ;
        RECT 1.420 2331.540 2324.000 2332.700 ;
        RECT 0.560 2328.220 2324.000 2331.540 ;
        RECT 1.420 2327.060 2324.000 2328.220 ;
        RECT 0.560 2323.740 2324.000 2327.060 ;
        RECT 1.420 2322.580 2324.000 2323.740 ;
        RECT 0.560 2319.260 2324.000 2322.580 ;
        RECT 1.420 2318.100 2324.000 2319.260 ;
        RECT 0.560 2314.780 2324.000 2318.100 ;
        RECT 1.420 2313.620 2324.000 2314.780 ;
        RECT 0.560 2310.300 2324.000 2313.620 ;
        RECT 1.420 2309.140 2324.000 2310.300 ;
        RECT 0.560 2305.820 2324.000 2309.140 ;
        RECT 1.420 2304.660 2324.000 2305.820 ;
        RECT 0.560 2301.340 2324.000 2304.660 ;
        RECT 1.420 2300.180 2324.000 2301.340 ;
        RECT 0.560 2296.860 2324.000 2300.180 ;
        RECT 1.420 2295.700 2324.000 2296.860 ;
        RECT 0.560 2292.380 2324.000 2295.700 ;
        RECT 1.420 2291.220 2324.000 2292.380 ;
        RECT 0.560 2287.900 2324.000 2291.220 ;
        RECT 1.420 2286.740 2324.000 2287.900 ;
        RECT 0.560 2283.420 2324.000 2286.740 ;
        RECT 1.420 2282.260 2324.000 2283.420 ;
        RECT 0.560 2278.940 2324.000 2282.260 ;
        RECT 1.420 2277.780 2324.000 2278.940 ;
        RECT 0.560 2274.460 2324.000 2277.780 ;
        RECT 1.420 2273.300 2324.000 2274.460 ;
        RECT 0.560 2269.980 2324.000 2273.300 ;
        RECT 1.420 2268.820 2324.000 2269.980 ;
        RECT 0.560 2265.500 2324.000 2268.820 ;
        RECT 1.420 2264.340 2324.000 2265.500 ;
        RECT 0.560 2261.020 2324.000 2264.340 ;
        RECT 1.420 2259.860 2324.000 2261.020 ;
        RECT 0.560 2256.540 2324.000 2259.860 ;
        RECT 1.420 2255.380 2324.000 2256.540 ;
        RECT 0.560 2252.060 2324.000 2255.380 ;
        RECT 1.420 2250.900 2324.000 2252.060 ;
        RECT 0.560 2247.580 2324.000 2250.900 ;
        RECT 1.420 2246.420 2324.000 2247.580 ;
        RECT 0.560 2243.100 2324.000 2246.420 ;
        RECT 1.420 2241.940 2324.000 2243.100 ;
        RECT 0.560 2238.620 2324.000 2241.940 ;
        RECT 1.420 2237.460 2324.000 2238.620 ;
        RECT 0.560 2234.140 2324.000 2237.460 ;
        RECT 1.420 2232.980 2324.000 2234.140 ;
        RECT 0.560 2229.660 2324.000 2232.980 ;
        RECT 1.420 2228.500 2324.000 2229.660 ;
        RECT 0.560 2225.180 2324.000 2228.500 ;
        RECT 1.420 2224.020 2324.000 2225.180 ;
        RECT 0.560 2220.700 2324.000 2224.020 ;
        RECT 1.420 2219.540 2324.000 2220.700 ;
        RECT 0.560 2216.220 2324.000 2219.540 ;
        RECT 1.420 2215.060 2324.000 2216.220 ;
        RECT 0.560 2211.740 2324.000 2215.060 ;
        RECT 1.420 2210.580 2324.000 2211.740 ;
        RECT 0.560 2207.260 2324.000 2210.580 ;
        RECT 1.420 2206.100 2324.000 2207.260 ;
        RECT 0.560 2202.780 2324.000 2206.100 ;
        RECT 1.420 2201.620 2324.000 2202.780 ;
        RECT 0.560 2198.300 2324.000 2201.620 ;
        RECT 1.420 2197.140 2324.000 2198.300 ;
        RECT 0.560 2193.820 2324.000 2197.140 ;
        RECT 1.420 2192.660 2324.000 2193.820 ;
        RECT 0.560 2189.340 2324.000 2192.660 ;
        RECT 1.420 2188.180 2324.000 2189.340 ;
        RECT 0.560 2184.860 2324.000 2188.180 ;
        RECT 1.420 2183.700 2324.000 2184.860 ;
        RECT 0.560 2180.380 2324.000 2183.700 ;
        RECT 1.420 2179.220 2324.000 2180.380 ;
        RECT 0.560 2175.900 2324.000 2179.220 ;
        RECT 1.420 2174.740 2324.000 2175.900 ;
        RECT 0.560 2171.420 2324.000 2174.740 ;
        RECT 1.420 2170.260 2324.000 2171.420 ;
        RECT 0.560 2166.940 2324.000 2170.260 ;
        RECT 1.420 2165.780 2324.000 2166.940 ;
        RECT 0.560 2162.460 2324.000 2165.780 ;
        RECT 1.420 2161.300 2324.000 2162.460 ;
        RECT 0.560 2157.980 2324.000 2161.300 ;
        RECT 1.420 2156.820 2324.000 2157.980 ;
        RECT 0.560 2153.500 2324.000 2156.820 ;
        RECT 1.420 2152.340 2324.000 2153.500 ;
        RECT 0.560 2149.020 2324.000 2152.340 ;
        RECT 1.420 2147.860 2324.000 2149.020 ;
        RECT 0.560 2144.540 2324.000 2147.860 ;
        RECT 1.420 2143.380 2324.000 2144.540 ;
        RECT 0.560 2140.060 2324.000 2143.380 ;
        RECT 1.420 2138.900 2324.000 2140.060 ;
        RECT 0.560 2135.580 2324.000 2138.900 ;
        RECT 1.420 2134.420 2324.000 2135.580 ;
        RECT 0.560 2131.100 2324.000 2134.420 ;
        RECT 1.420 2129.940 2324.000 2131.100 ;
        RECT 0.560 2126.620 2324.000 2129.940 ;
        RECT 1.420 2125.460 2324.000 2126.620 ;
        RECT 0.560 2122.140 2324.000 2125.460 ;
        RECT 1.420 2120.980 2324.000 2122.140 ;
        RECT 0.560 2117.660 2324.000 2120.980 ;
        RECT 1.420 2116.500 2324.000 2117.660 ;
        RECT 0.560 2113.180 2324.000 2116.500 ;
        RECT 1.420 2112.020 2324.000 2113.180 ;
        RECT 0.560 2108.700 2324.000 2112.020 ;
        RECT 1.420 2107.540 2324.000 2108.700 ;
        RECT 0.560 2104.220 2324.000 2107.540 ;
        RECT 1.420 2103.060 2324.000 2104.220 ;
        RECT 0.560 2099.740 2324.000 2103.060 ;
        RECT 1.420 2098.580 2324.000 2099.740 ;
        RECT 0.560 2076.780 2324.000 2098.580 ;
        RECT 1.420 2075.620 2324.000 2076.780 ;
        RECT 0.560 2072.300 2324.000 2075.620 ;
        RECT 1.420 2071.140 2324.000 2072.300 ;
        RECT 0.560 2067.820 2324.000 2071.140 ;
        RECT 1.420 2066.660 2324.000 2067.820 ;
        RECT 0.560 2063.340 2324.000 2066.660 ;
        RECT 1.420 2062.180 2324.000 2063.340 ;
        RECT 0.560 2058.860 2324.000 2062.180 ;
        RECT 1.420 2057.700 2324.000 2058.860 ;
        RECT 0.560 2054.380 2324.000 2057.700 ;
        RECT 1.420 2053.220 2324.000 2054.380 ;
        RECT 0.560 2049.900 2324.000 2053.220 ;
        RECT 1.420 2048.740 2324.000 2049.900 ;
        RECT 0.560 2045.420 2324.000 2048.740 ;
        RECT 1.420 2044.260 2324.000 2045.420 ;
        RECT 0.560 2040.940 2324.000 2044.260 ;
        RECT 1.420 2039.780 2324.000 2040.940 ;
        RECT 0.560 2036.460 2324.000 2039.780 ;
        RECT 1.420 2035.300 2324.000 2036.460 ;
        RECT 0.560 2031.980 2324.000 2035.300 ;
        RECT 1.420 2030.820 2324.000 2031.980 ;
        RECT 0.560 2027.500 2324.000 2030.820 ;
        RECT 1.420 2026.340 2324.000 2027.500 ;
        RECT 0.560 2023.020 2324.000 2026.340 ;
        RECT 1.420 2021.860 2324.000 2023.020 ;
        RECT 0.560 2018.540 2324.000 2021.860 ;
        RECT 1.420 2017.380 2324.000 2018.540 ;
        RECT 0.560 2014.060 2324.000 2017.380 ;
        RECT 1.420 2012.900 2324.000 2014.060 ;
        RECT 0.560 2009.580 2324.000 2012.900 ;
        RECT 1.420 2008.420 2324.000 2009.580 ;
        RECT 0.560 2005.100 2324.000 2008.420 ;
        RECT 1.420 2003.940 2324.000 2005.100 ;
        RECT 0.560 2000.620 2324.000 2003.940 ;
        RECT 1.420 1999.460 2324.000 2000.620 ;
        RECT 0.560 1996.140 2324.000 1999.460 ;
        RECT 1.420 1994.980 2324.000 1996.140 ;
        RECT 0.560 1991.660 2324.000 1994.980 ;
        RECT 1.420 1990.500 2324.000 1991.660 ;
        RECT 0.560 1987.180 2324.000 1990.500 ;
        RECT 1.420 1986.020 2324.000 1987.180 ;
        RECT 0.560 1982.700 2324.000 1986.020 ;
        RECT 1.420 1981.540 2324.000 1982.700 ;
        RECT 0.560 1978.220 2324.000 1981.540 ;
        RECT 1.420 1977.100 2324.000 1978.220 ;
        RECT 1.420 1977.060 2323.140 1977.100 ;
        RECT 0.560 1975.940 2323.140 1977.060 ;
        RECT 0.560 1973.740 2324.000 1975.940 ;
        RECT 1.420 1972.620 2324.000 1973.740 ;
        RECT 1.420 1972.580 2323.140 1972.620 ;
        RECT 0.560 1971.460 2323.140 1972.580 ;
        RECT 0.560 1969.260 2324.000 1971.460 ;
        RECT 1.420 1968.140 2324.000 1969.260 ;
        RECT 1.420 1968.100 2323.140 1968.140 ;
        RECT 0.560 1966.980 2323.140 1968.100 ;
        RECT 0.560 1964.780 2324.000 1966.980 ;
        RECT 1.420 1963.660 2324.000 1964.780 ;
        RECT 1.420 1963.620 2323.140 1963.660 ;
        RECT 0.560 1962.500 2323.140 1963.620 ;
        RECT 0.560 1960.300 2324.000 1962.500 ;
        RECT 1.420 1959.180 2324.000 1960.300 ;
        RECT 1.420 1959.140 2323.140 1959.180 ;
        RECT 0.560 1958.020 2323.140 1959.140 ;
        RECT 0.560 1955.820 2324.000 1958.020 ;
        RECT 1.420 1954.700 2324.000 1955.820 ;
        RECT 1.420 1954.660 2323.140 1954.700 ;
        RECT 0.560 1953.540 2323.140 1954.660 ;
        RECT 0.560 1951.340 2324.000 1953.540 ;
        RECT 1.420 1950.220 2324.000 1951.340 ;
        RECT 1.420 1950.180 2323.140 1950.220 ;
        RECT 0.560 1949.060 2323.140 1950.180 ;
        RECT 0.560 1946.860 2324.000 1949.060 ;
        RECT 1.420 1945.740 2324.000 1946.860 ;
        RECT 1.420 1945.700 2323.140 1945.740 ;
        RECT 0.560 1944.580 2323.140 1945.700 ;
        RECT 0.560 1942.380 2324.000 1944.580 ;
        RECT 1.420 1941.260 2324.000 1942.380 ;
        RECT 1.420 1941.220 2323.140 1941.260 ;
        RECT 0.560 1940.100 2323.140 1941.220 ;
        RECT 0.560 1937.900 2324.000 1940.100 ;
        RECT 1.420 1936.780 2324.000 1937.900 ;
        RECT 1.420 1936.740 2323.140 1936.780 ;
        RECT 0.560 1935.620 2323.140 1936.740 ;
        RECT 0.560 1933.420 2324.000 1935.620 ;
        RECT 1.420 1932.300 2324.000 1933.420 ;
        RECT 1.420 1932.260 2323.140 1932.300 ;
        RECT 0.560 1931.140 2323.140 1932.260 ;
        RECT 0.560 1928.940 2324.000 1931.140 ;
        RECT 1.420 1927.820 2324.000 1928.940 ;
        RECT 1.420 1927.780 2323.140 1927.820 ;
        RECT 0.560 1926.660 2323.140 1927.780 ;
        RECT 0.560 1924.460 2324.000 1926.660 ;
        RECT 1.420 1923.340 2324.000 1924.460 ;
        RECT 1.420 1923.300 2323.140 1923.340 ;
        RECT 0.560 1922.180 2323.140 1923.300 ;
        RECT 0.560 1919.980 2324.000 1922.180 ;
        RECT 1.420 1918.860 2324.000 1919.980 ;
        RECT 1.420 1918.820 2323.140 1918.860 ;
        RECT 0.560 1917.700 2323.140 1918.820 ;
        RECT 0.560 1915.500 2324.000 1917.700 ;
        RECT 1.420 1914.380 2324.000 1915.500 ;
        RECT 1.420 1914.340 2323.140 1914.380 ;
        RECT 0.560 1913.220 2323.140 1914.340 ;
        RECT 0.560 1911.020 2324.000 1913.220 ;
        RECT 1.420 1909.900 2324.000 1911.020 ;
        RECT 1.420 1909.860 2323.140 1909.900 ;
        RECT 0.560 1908.740 2323.140 1909.860 ;
        RECT 0.560 1906.540 2324.000 1908.740 ;
        RECT 1.420 1905.420 2324.000 1906.540 ;
        RECT 1.420 1905.380 2323.140 1905.420 ;
        RECT 0.560 1904.260 2323.140 1905.380 ;
        RECT 0.560 1902.060 2324.000 1904.260 ;
        RECT 1.420 1900.940 2324.000 1902.060 ;
        RECT 1.420 1900.900 2323.140 1900.940 ;
        RECT 0.560 1899.780 2323.140 1900.900 ;
        RECT 0.560 1897.580 2324.000 1899.780 ;
        RECT 1.420 1896.460 2324.000 1897.580 ;
        RECT 1.420 1896.420 2323.140 1896.460 ;
        RECT 0.560 1895.300 2323.140 1896.420 ;
        RECT 0.560 1893.100 2324.000 1895.300 ;
        RECT 1.420 1891.980 2324.000 1893.100 ;
        RECT 1.420 1891.940 2323.140 1891.980 ;
        RECT 0.560 1890.820 2323.140 1891.940 ;
        RECT 0.560 1888.620 2324.000 1890.820 ;
        RECT 1.420 1887.500 2324.000 1888.620 ;
        RECT 1.420 1887.460 2323.140 1887.500 ;
        RECT 0.560 1886.340 2323.140 1887.460 ;
        RECT 0.560 1884.140 2324.000 1886.340 ;
        RECT 1.420 1883.020 2324.000 1884.140 ;
        RECT 1.420 1882.980 2323.140 1883.020 ;
        RECT 0.560 1881.860 2323.140 1882.980 ;
        RECT 0.560 1879.660 2324.000 1881.860 ;
        RECT 1.420 1878.540 2324.000 1879.660 ;
        RECT 1.420 1878.500 2323.140 1878.540 ;
        RECT 0.560 1877.380 2323.140 1878.500 ;
        RECT 0.560 1875.180 2324.000 1877.380 ;
        RECT 1.420 1874.060 2324.000 1875.180 ;
        RECT 1.420 1874.020 2323.140 1874.060 ;
        RECT 0.560 1872.900 2323.140 1874.020 ;
        RECT 0.560 1870.700 2324.000 1872.900 ;
        RECT 1.420 1869.580 2324.000 1870.700 ;
        RECT 1.420 1869.540 2323.140 1869.580 ;
        RECT 0.560 1868.420 2323.140 1869.540 ;
        RECT 0.560 1866.220 2324.000 1868.420 ;
        RECT 1.420 1865.100 2324.000 1866.220 ;
        RECT 1.420 1865.060 2323.140 1865.100 ;
        RECT 0.560 1863.940 2323.140 1865.060 ;
        RECT 0.560 1861.740 2324.000 1863.940 ;
        RECT 1.420 1860.620 2324.000 1861.740 ;
        RECT 1.420 1860.580 2323.140 1860.620 ;
        RECT 0.560 1859.460 2323.140 1860.580 ;
        RECT 0.560 1857.260 2324.000 1859.460 ;
        RECT 1.420 1856.140 2324.000 1857.260 ;
        RECT 1.420 1856.100 2323.140 1856.140 ;
        RECT 0.560 1854.980 2323.140 1856.100 ;
        RECT 0.560 1852.780 2324.000 1854.980 ;
        RECT 1.420 1851.660 2324.000 1852.780 ;
        RECT 1.420 1851.620 2323.140 1851.660 ;
        RECT 0.560 1850.500 2323.140 1851.620 ;
        RECT 0.560 1848.300 2324.000 1850.500 ;
        RECT 1.420 1847.180 2324.000 1848.300 ;
        RECT 1.420 1847.140 2323.140 1847.180 ;
        RECT 0.560 1846.020 2323.140 1847.140 ;
        RECT 0.560 1843.820 2324.000 1846.020 ;
        RECT 1.420 1842.700 2324.000 1843.820 ;
        RECT 1.420 1842.660 2323.140 1842.700 ;
        RECT 0.560 1841.540 2323.140 1842.660 ;
        RECT 0.560 1839.340 2324.000 1841.540 ;
        RECT 1.420 1838.220 2324.000 1839.340 ;
        RECT 1.420 1838.180 2323.140 1838.220 ;
        RECT 0.560 1837.060 2323.140 1838.180 ;
        RECT 0.560 1834.860 2324.000 1837.060 ;
        RECT 1.420 1833.740 2324.000 1834.860 ;
        RECT 1.420 1833.700 2323.140 1833.740 ;
        RECT 0.560 1832.580 2323.140 1833.700 ;
        RECT 0.560 1830.380 2324.000 1832.580 ;
        RECT 1.420 1829.260 2324.000 1830.380 ;
        RECT 1.420 1829.220 2323.140 1829.260 ;
        RECT 0.560 1828.100 2323.140 1829.220 ;
        RECT 0.560 1825.900 2324.000 1828.100 ;
        RECT 1.420 1824.780 2324.000 1825.900 ;
        RECT 1.420 1824.740 2323.140 1824.780 ;
        RECT 0.560 1823.620 2323.140 1824.740 ;
        RECT 0.560 1821.420 2324.000 1823.620 ;
        RECT 1.420 1820.300 2324.000 1821.420 ;
        RECT 1.420 1820.260 2323.140 1820.300 ;
        RECT 0.560 1819.140 2323.140 1820.260 ;
        RECT 0.560 1816.940 2324.000 1819.140 ;
        RECT 1.420 1815.820 2324.000 1816.940 ;
        RECT 1.420 1815.780 2323.140 1815.820 ;
        RECT 0.560 1814.660 2323.140 1815.780 ;
        RECT 0.560 1812.460 2324.000 1814.660 ;
        RECT 1.420 1811.300 2324.000 1812.460 ;
        RECT 0.560 1789.500 2324.000 1811.300 ;
        RECT 1.420 1788.340 2324.000 1789.500 ;
        RECT 0.560 1785.020 2324.000 1788.340 ;
        RECT 1.420 1783.860 2324.000 1785.020 ;
        RECT 0.560 1780.540 2324.000 1783.860 ;
        RECT 1.420 1779.380 2324.000 1780.540 ;
        RECT 0.560 1776.060 2324.000 1779.380 ;
        RECT 1.420 1774.900 2324.000 1776.060 ;
        RECT 0.560 1771.580 2324.000 1774.900 ;
        RECT 1.420 1770.420 2324.000 1771.580 ;
        RECT 0.560 1767.100 2324.000 1770.420 ;
        RECT 1.420 1765.940 2324.000 1767.100 ;
        RECT 0.560 1762.620 2324.000 1765.940 ;
        RECT 1.420 1761.460 2324.000 1762.620 ;
        RECT 0.560 1758.140 2324.000 1761.460 ;
        RECT 1.420 1756.980 2324.000 1758.140 ;
        RECT 0.560 1753.660 2324.000 1756.980 ;
        RECT 1.420 1752.500 2324.000 1753.660 ;
        RECT 0.560 1749.180 2324.000 1752.500 ;
        RECT 1.420 1748.020 2324.000 1749.180 ;
        RECT 0.560 1744.700 2324.000 1748.020 ;
        RECT 1.420 1743.540 2324.000 1744.700 ;
        RECT 0.560 1740.220 2324.000 1743.540 ;
        RECT 1.420 1739.060 2324.000 1740.220 ;
        RECT 0.560 1735.740 2324.000 1739.060 ;
        RECT 1.420 1734.580 2324.000 1735.740 ;
        RECT 0.560 1731.260 2324.000 1734.580 ;
        RECT 1.420 1730.100 2324.000 1731.260 ;
        RECT 0.560 1726.780 2324.000 1730.100 ;
        RECT 1.420 1725.620 2324.000 1726.780 ;
        RECT 0.560 1722.300 2324.000 1725.620 ;
        RECT 1.420 1721.140 2324.000 1722.300 ;
        RECT 0.560 1717.820 2324.000 1721.140 ;
        RECT 1.420 1716.660 2324.000 1717.820 ;
        RECT 0.560 1713.340 2324.000 1716.660 ;
        RECT 1.420 1712.180 2324.000 1713.340 ;
        RECT 0.560 1708.860 2324.000 1712.180 ;
        RECT 1.420 1707.700 2324.000 1708.860 ;
        RECT 0.560 1704.380 2324.000 1707.700 ;
        RECT 1.420 1703.220 2324.000 1704.380 ;
        RECT 0.560 1699.900 2324.000 1703.220 ;
        RECT 1.420 1698.740 2324.000 1699.900 ;
        RECT 0.560 1695.420 2324.000 1698.740 ;
        RECT 1.420 1694.260 2324.000 1695.420 ;
        RECT 0.560 1690.940 2324.000 1694.260 ;
        RECT 1.420 1689.780 2324.000 1690.940 ;
        RECT 0.560 1686.460 2324.000 1689.780 ;
        RECT 1.420 1685.300 2324.000 1686.460 ;
        RECT 0.560 1681.980 2324.000 1685.300 ;
        RECT 1.420 1680.820 2324.000 1681.980 ;
        RECT 0.560 1677.500 2324.000 1680.820 ;
        RECT 1.420 1676.340 2324.000 1677.500 ;
        RECT 0.560 1673.020 2324.000 1676.340 ;
        RECT 1.420 1671.860 2324.000 1673.020 ;
        RECT 0.560 1668.540 2324.000 1671.860 ;
        RECT 1.420 1667.380 2324.000 1668.540 ;
        RECT 0.560 1664.060 2324.000 1667.380 ;
        RECT 1.420 1662.900 2324.000 1664.060 ;
        RECT 0.560 1659.580 2324.000 1662.900 ;
        RECT 1.420 1658.420 2324.000 1659.580 ;
        RECT 0.560 1655.100 2324.000 1658.420 ;
        RECT 1.420 1653.940 2324.000 1655.100 ;
        RECT 0.560 1650.620 2324.000 1653.940 ;
        RECT 1.420 1649.460 2324.000 1650.620 ;
        RECT 0.560 1646.140 2324.000 1649.460 ;
        RECT 1.420 1644.980 2324.000 1646.140 ;
        RECT 0.560 1641.660 2324.000 1644.980 ;
        RECT 1.420 1640.500 2324.000 1641.660 ;
        RECT 0.560 1637.180 2324.000 1640.500 ;
        RECT 1.420 1636.020 2324.000 1637.180 ;
        RECT 0.560 1632.700 2324.000 1636.020 ;
        RECT 1.420 1631.540 2324.000 1632.700 ;
        RECT 0.560 1628.220 2324.000 1631.540 ;
        RECT 1.420 1627.060 2324.000 1628.220 ;
        RECT 0.560 1623.740 2324.000 1627.060 ;
        RECT 1.420 1622.580 2324.000 1623.740 ;
        RECT 0.560 1619.260 2324.000 1622.580 ;
        RECT 1.420 1618.100 2324.000 1619.260 ;
        RECT 0.560 1614.780 2324.000 1618.100 ;
        RECT 1.420 1613.620 2324.000 1614.780 ;
        RECT 0.560 1610.300 2324.000 1613.620 ;
        RECT 1.420 1609.140 2324.000 1610.300 ;
        RECT 0.560 1605.820 2324.000 1609.140 ;
        RECT 1.420 1604.660 2324.000 1605.820 ;
        RECT 0.560 1601.340 2324.000 1604.660 ;
        RECT 1.420 1600.180 2324.000 1601.340 ;
        RECT 0.560 1596.860 2324.000 1600.180 ;
        RECT 1.420 1595.700 2324.000 1596.860 ;
        RECT 0.560 1592.380 2324.000 1595.700 ;
        RECT 1.420 1591.220 2324.000 1592.380 ;
        RECT 0.560 1587.900 2324.000 1591.220 ;
        RECT 1.420 1586.740 2324.000 1587.900 ;
        RECT 0.560 1583.420 2324.000 1586.740 ;
        RECT 1.420 1582.260 2324.000 1583.420 ;
        RECT 0.560 1578.940 2324.000 1582.260 ;
        RECT 1.420 1577.780 2324.000 1578.940 ;
        RECT 0.560 1574.460 2324.000 1577.780 ;
        RECT 1.420 1573.300 2324.000 1574.460 ;
        RECT 0.560 1569.980 2324.000 1573.300 ;
        RECT 1.420 1568.820 2324.000 1569.980 ;
        RECT 0.560 1565.500 2324.000 1568.820 ;
        RECT 1.420 1564.340 2324.000 1565.500 ;
        RECT 0.560 1561.020 2324.000 1564.340 ;
        RECT 1.420 1559.860 2324.000 1561.020 ;
        RECT 0.560 1556.540 2324.000 1559.860 ;
        RECT 1.420 1555.380 2324.000 1556.540 ;
        RECT 0.560 1552.060 2324.000 1555.380 ;
        RECT 1.420 1550.900 2324.000 1552.060 ;
        RECT 0.560 1547.580 2324.000 1550.900 ;
        RECT 1.420 1546.420 2324.000 1547.580 ;
        RECT 0.560 1543.100 2324.000 1546.420 ;
        RECT 1.420 1541.940 2324.000 1543.100 ;
        RECT 0.560 1538.620 2324.000 1541.940 ;
        RECT 1.420 1537.460 2324.000 1538.620 ;
        RECT 0.560 1534.140 2324.000 1537.460 ;
        RECT 1.420 1532.980 2324.000 1534.140 ;
        RECT 0.560 1529.660 2324.000 1532.980 ;
        RECT 1.420 1528.500 2324.000 1529.660 ;
        RECT 0.560 1525.180 2324.000 1528.500 ;
        RECT 1.420 1524.020 2324.000 1525.180 ;
        RECT 0.560 1502.220 2324.000 1524.020 ;
        RECT 1.420 1501.060 2324.000 1502.220 ;
        RECT 0.560 1497.740 2324.000 1501.060 ;
        RECT 1.420 1496.580 2324.000 1497.740 ;
        RECT 0.560 1493.260 2324.000 1496.580 ;
        RECT 1.420 1492.100 2324.000 1493.260 ;
        RECT 0.560 1488.780 2324.000 1492.100 ;
        RECT 1.420 1487.620 2324.000 1488.780 ;
        RECT 0.560 1484.300 2324.000 1487.620 ;
        RECT 1.420 1483.140 2324.000 1484.300 ;
        RECT 0.560 1479.820 2324.000 1483.140 ;
        RECT 1.420 1478.660 2324.000 1479.820 ;
        RECT 0.560 1475.340 2324.000 1478.660 ;
        RECT 1.420 1474.180 2324.000 1475.340 ;
        RECT 0.560 1470.860 2324.000 1474.180 ;
        RECT 1.420 1469.700 2324.000 1470.860 ;
        RECT 0.560 1466.380 2324.000 1469.700 ;
        RECT 1.420 1465.220 2324.000 1466.380 ;
        RECT 0.560 1461.900 2324.000 1465.220 ;
        RECT 1.420 1460.740 2324.000 1461.900 ;
        RECT 0.560 1457.420 2324.000 1460.740 ;
        RECT 1.420 1456.260 2324.000 1457.420 ;
        RECT 0.560 1452.940 2324.000 1456.260 ;
        RECT 1.420 1451.780 2324.000 1452.940 ;
        RECT 0.560 1448.460 2324.000 1451.780 ;
        RECT 1.420 1447.300 2324.000 1448.460 ;
        RECT 0.560 1443.980 2324.000 1447.300 ;
        RECT 1.420 1442.820 2324.000 1443.980 ;
        RECT 0.560 1439.500 2324.000 1442.820 ;
        RECT 1.420 1438.340 2324.000 1439.500 ;
        RECT 0.560 1435.020 2324.000 1438.340 ;
        RECT 1.420 1433.860 2324.000 1435.020 ;
        RECT 0.560 1430.540 2324.000 1433.860 ;
        RECT 1.420 1429.380 2324.000 1430.540 ;
        RECT 0.560 1426.060 2324.000 1429.380 ;
        RECT 1.420 1424.900 2324.000 1426.060 ;
        RECT 0.560 1421.580 2324.000 1424.900 ;
        RECT 1.420 1420.420 2324.000 1421.580 ;
        RECT 0.560 1417.100 2324.000 1420.420 ;
        RECT 1.420 1415.940 2324.000 1417.100 ;
        RECT 0.560 1412.620 2324.000 1415.940 ;
        RECT 1.420 1411.460 2324.000 1412.620 ;
        RECT 0.560 1408.140 2324.000 1411.460 ;
        RECT 1.420 1406.980 2324.000 1408.140 ;
        RECT 0.560 1403.660 2324.000 1406.980 ;
        RECT 1.420 1402.540 2324.000 1403.660 ;
        RECT 1.420 1402.500 2323.140 1402.540 ;
        RECT 0.560 1401.380 2323.140 1402.500 ;
        RECT 0.560 1399.180 2324.000 1401.380 ;
        RECT 1.420 1398.060 2324.000 1399.180 ;
        RECT 1.420 1398.020 2323.140 1398.060 ;
        RECT 0.560 1396.900 2323.140 1398.020 ;
        RECT 0.560 1394.700 2324.000 1396.900 ;
        RECT 1.420 1393.580 2324.000 1394.700 ;
        RECT 1.420 1393.540 2323.140 1393.580 ;
        RECT 0.560 1392.420 2323.140 1393.540 ;
        RECT 0.560 1390.220 2324.000 1392.420 ;
        RECT 1.420 1389.100 2324.000 1390.220 ;
        RECT 1.420 1389.060 2323.140 1389.100 ;
        RECT 0.560 1387.940 2323.140 1389.060 ;
        RECT 0.560 1385.740 2324.000 1387.940 ;
        RECT 1.420 1384.620 2324.000 1385.740 ;
        RECT 1.420 1384.580 2323.140 1384.620 ;
        RECT 0.560 1383.460 2323.140 1384.580 ;
        RECT 0.560 1381.260 2324.000 1383.460 ;
        RECT 1.420 1380.140 2324.000 1381.260 ;
        RECT 1.420 1380.100 2323.140 1380.140 ;
        RECT 0.560 1378.980 2323.140 1380.100 ;
        RECT 0.560 1376.780 2324.000 1378.980 ;
        RECT 1.420 1375.660 2324.000 1376.780 ;
        RECT 1.420 1375.620 2323.140 1375.660 ;
        RECT 0.560 1374.500 2323.140 1375.620 ;
        RECT 0.560 1372.300 2324.000 1374.500 ;
        RECT 1.420 1371.180 2324.000 1372.300 ;
        RECT 1.420 1371.140 2323.140 1371.180 ;
        RECT 0.560 1370.020 2323.140 1371.140 ;
        RECT 0.560 1367.820 2324.000 1370.020 ;
        RECT 1.420 1366.700 2324.000 1367.820 ;
        RECT 1.420 1366.660 2323.140 1366.700 ;
        RECT 0.560 1365.540 2323.140 1366.660 ;
        RECT 0.560 1363.340 2324.000 1365.540 ;
        RECT 1.420 1362.220 2324.000 1363.340 ;
        RECT 1.420 1362.180 2323.140 1362.220 ;
        RECT 0.560 1361.060 2323.140 1362.180 ;
        RECT 0.560 1358.860 2324.000 1361.060 ;
        RECT 1.420 1357.740 2324.000 1358.860 ;
        RECT 1.420 1357.700 2323.140 1357.740 ;
        RECT 0.560 1356.580 2323.140 1357.700 ;
        RECT 0.560 1354.380 2324.000 1356.580 ;
        RECT 1.420 1353.260 2324.000 1354.380 ;
        RECT 1.420 1353.220 2323.140 1353.260 ;
        RECT 0.560 1352.100 2323.140 1353.220 ;
        RECT 0.560 1349.900 2324.000 1352.100 ;
        RECT 1.420 1348.780 2324.000 1349.900 ;
        RECT 1.420 1348.740 2323.140 1348.780 ;
        RECT 0.560 1347.620 2323.140 1348.740 ;
        RECT 0.560 1345.420 2324.000 1347.620 ;
        RECT 1.420 1344.300 2324.000 1345.420 ;
        RECT 1.420 1344.260 2323.140 1344.300 ;
        RECT 0.560 1343.140 2323.140 1344.260 ;
        RECT 0.560 1340.940 2324.000 1343.140 ;
        RECT 1.420 1339.820 2324.000 1340.940 ;
        RECT 1.420 1339.780 2323.140 1339.820 ;
        RECT 0.560 1338.660 2323.140 1339.780 ;
        RECT 0.560 1336.460 2324.000 1338.660 ;
        RECT 1.420 1335.340 2324.000 1336.460 ;
        RECT 1.420 1335.300 2323.140 1335.340 ;
        RECT 0.560 1334.180 2323.140 1335.300 ;
        RECT 0.560 1331.980 2324.000 1334.180 ;
        RECT 1.420 1330.860 2324.000 1331.980 ;
        RECT 1.420 1330.820 2323.140 1330.860 ;
        RECT 0.560 1329.700 2323.140 1330.820 ;
        RECT 0.560 1327.500 2324.000 1329.700 ;
        RECT 1.420 1326.380 2324.000 1327.500 ;
        RECT 1.420 1326.340 2323.140 1326.380 ;
        RECT 0.560 1325.220 2323.140 1326.340 ;
        RECT 0.560 1323.020 2324.000 1325.220 ;
        RECT 1.420 1321.900 2324.000 1323.020 ;
        RECT 1.420 1321.860 2323.140 1321.900 ;
        RECT 0.560 1320.740 2323.140 1321.860 ;
        RECT 0.560 1318.540 2324.000 1320.740 ;
        RECT 1.420 1317.420 2324.000 1318.540 ;
        RECT 1.420 1317.380 2323.140 1317.420 ;
        RECT 0.560 1316.260 2323.140 1317.380 ;
        RECT 0.560 1314.060 2324.000 1316.260 ;
        RECT 1.420 1312.940 2324.000 1314.060 ;
        RECT 1.420 1312.900 2323.140 1312.940 ;
        RECT 0.560 1311.780 2323.140 1312.900 ;
        RECT 0.560 1309.580 2324.000 1311.780 ;
        RECT 1.420 1308.460 2324.000 1309.580 ;
        RECT 1.420 1308.420 2323.140 1308.460 ;
        RECT 0.560 1307.300 2323.140 1308.420 ;
        RECT 0.560 1305.100 2324.000 1307.300 ;
        RECT 1.420 1303.980 2324.000 1305.100 ;
        RECT 1.420 1303.940 2323.140 1303.980 ;
        RECT 0.560 1302.820 2323.140 1303.940 ;
        RECT 0.560 1300.620 2324.000 1302.820 ;
        RECT 1.420 1299.500 2324.000 1300.620 ;
        RECT 1.420 1299.460 2323.140 1299.500 ;
        RECT 0.560 1298.340 2323.140 1299.460 ;
        RECT 0.560 1296.140 2324.000 1298.340 ;
        RECT 1.420 1295.020 2324.000 1296.140 ;
        RECT 1.420 1294.980 2323.140 1295.020 ;
        RECT 0.560 1293.860 2323.140 1294.980 ;
        RECT 0.560 1291.660 2324.000 1293.860 ;
        RECT 1.420 1290.540 2324.000 1291.660 ;
        RECT 1.420 1290.500 2323.140 1290.540 ;
        RECT 0.560 1289.380 2323.140 1290.500 ;
        RECT 0.560 1287.180 2324.000 1289.380 ;
        RECT 1.420 1286.060 2324.000 1287.180 ;
        RECT 1.420 1286.020 2323.140 1286.060 ;
        RECT 0.560 1284.900 2323.140 1286.020 ;
        RECT 0.560 1282.700 2324.000 1284.900 ;
        RECT 1.420 1281.580 2324.000 1282.700 ;
        RECT 1.420 1281.540 2323.140 1281.580 ;
        RECT 0.560 1280.420 2323.140 1281.540 ;
        RECT 0.560 1278.220 2324.000 1280.420 ;
        RECT 1.420 1277.100 2324.000 1278.220 ;
        RECT 1.420 1277.060 2323.140 1277.100 ;
        RECT 0.560 1275.940 2323.140 1277.060 ;
        RECT 0.560 1273.740 2324.000 1275.940 ;
        RECT 1.420 1272.620 2324.000 1273.740 ;
        RECT 1.420 1272.580 2323.140 1272.620 ;
        RECT 0.560 1271.460 2323.140 1272.580 ;
        RECT 0.560 1269.260 2324.000 1271.460 ;
        RECT 1.420 1268.140 2324.000 1269.260 ;
        RECT 1.420 1268.100 2323.140 1268.140 ;
        RECT 0.560 1266.980 2323.140 1268.100 ;
        RECT 0.560 1264.780 2324.000 1266.980 ;
        RECT 1.420 1263.660 2324.000 1264.780 ;
        RECT 1.420 1263.620 2323.140 1263.660 ;
        RECT 0.560 1262.500 2323.140 1263.620 ;
        RECT 0.560 1260.300 2324.000 1262.500 ;
        RECT 1.420 1259.180 2324.000 1260.300 ;
        RECT 1.420 1259.140 2323.140 1259.180 ;
        RECT 0.560 1258.020 2323.140 1259.140 ;
        RECT 0.560 1255.820 2324.000 1258.020 ;
        RECT 1.420 1254.700 2324.000 1255.820 ;
        RECT 1.420 1254.660 2323.140 1254.700 ;
        RECT 0.560 1253.540 2323.140 1254.660 ;
        RECT 0.560 1251.340 2324.000 1253.540 ;
        RECT 1.420 1250.220 2324.000 1251.340 ;
        RECT 1.420 1250.180 2323.140 1250.220 ;
        RECT 0.560 1249.060 2323.140 1250.180 ;
        RECT 0.560 1246.860 2324.000 1249.060 ;
        RECT 1.420 1245.740 2324.000 1246.860 ;
        RECT 1.420 1245.700 2323.140 1245.740 ;
        RECT 0.560 1244.580 2323.140 1245.700 ;
        RECT 0.560 1242.380 2324.000 1244.580 ;
        RECT 1.420 1241.260 2324.000 1242.380 ;
        RECT 1.420 1241.220 2323.140 1241.260 ;
        RECT 0.560 1240.100 2323.140 1241.220 ;
        RECT 0.560 1237.900 2324.000 1240.100 ;
        RECT 1.420 1236.740 2324.000 1237.900 ;
        RECT 0.560 1214.940 2324.000 1236.740 ;
        RECT 1.420 1213.780 2324.000 1214.940 ;
        RECT 0.560 1210.460 2324.000 1213.780 ;
        RECT 1.420 1209.300 2324.000 1210.460 ;
        RECT 0.560 1205.980 2324.000 1209.300 ;
        RECT 1.420 1204.820 2324.000 1205.980 ;
        RECT 0.560 1201.500 2324.000 1204.820 ;
        RECT 1.420 1200.340 2324.000 1201.500 ;
        RECT 0.560 1197.020 2324.000 1200.340 ;
        RECT 1.420 1195.860 2324.000 1197.020 ;
        RECT 0.560 1192.540 2324.000 1195.860 ;
        RECT 1.420 1191.380 2324.000 1192.540 ;
        RECT 0.560 1188.060 2324.000 1191.380 ;
        RECT 1.420 1186.900 2324.000 1188.060 ;
        RECT 0.560 1183.580 2324.000 1186.900 ;
        RECT 1.420 1182.420 2324.000 1183.580 ;
        RECT 0.560 1179.100 2324.000 1182.420 ;
        RECT 1.420 1177.940 2324.000 1179.100 ;
        RECT 0.560 1174.620 2324.000 1177.940 ;
        RECT 1.420 1173.460 2324.000 1174.620 ;
        RECT 0.560 1170.140 2324.000 1173.460 ;
        RECT 1.420 1168.980 2324.000 1170.140 ;
        RECT 0.560 1165.660 2324.000 1168.980 ;
        RECT 1.420 1164.500 2324.000 1165.660 ;
        RECT 0.560 1161.180 2324.000 1164.500 ;
        RECT 1.420 1160.020 2324.000 1161.180 ;
        RECT 0.560 1156.700 2324.000 1160.020 ;
        RECT 1.420 1155.540 2324.000 1156.700 ;
        RECT 0.560 1152.220 2324.000 1155.540 ;
        RECT 1.420 1151.060 2324.000 1152.220 ;
        RECT 0.560 1147.740 2324.000 1151.060 ;
        RECT 1.420 1146.580 2324.000 1147.740 ;
        RECT 0.560 1143.260 2324.000 1146.580 ;
        RECT 1.420 1142.100 2324.000 1143.260 ;
        RECT 0.560 1138.780 2324.000 1142.100 ;
        RECT 1.420 1137.620 2324.000 1138.780 ;
        RECT 0.560 1134.300 2324.000 1137.620 ;
        RECT 1.420 1133.140 2324.000 1134.300 ;
        RECT 0.560 1129.820 2324.000 1133.140 ;
        RECT 1.420 1128.660 2324.000 1129.820 ;
        RECT 0.560 1125.340 2324.000 1128.660 ;
        RECT 1.420 1124.180 2324.000 1125.340 ;
        RECT 0.560 1120.860 2324.000 1124.180 ;
        RECT 1.420 1119.700 2324.000 1120.860 ;
        RECT 0.560 1116.380 2324.000 1119.700 ;
        RECT 1.420 1115.220 2324.000 1116.380 ;
        RECT 0.560 1111.900 2324.000 1115.220 ;
        RECT 1.420 1110.740 2324.000 1111.900 ;
        RECT 0.560 1107.420 2324.000 1110.740 ;
        RECT 1.420 1106.260 2324.000 1107.420 ;
        RECT 0.560 1102.940 2324.000 1106.260 ;
        RECT 1.420 1101.780 2324.000 1102.940 ;
        RECT 0.560 1098.460 2324.000 1101.780 ;
        RECT 1.420 1097.300 2324.000 1098.460 ;
        RECT 0.560 1093.980 2324.000 1097.300 ;
        RECT 1.420 1092.820 2324.000 1093.980 ;
        RECT 0.560 1089.500 2324.000 1092.820 ;
        RECT 1.420 1088.340 2324.000 1089.500 ;
        RECT 0.560 1085.020 2324.000 1088.340 ;
        RECT 1.420 1083.860 2324.000 1085.020 ;
        RECT 0.560 1080.540 2324.000 1083.860 ;
        RECT 1.420 1079.380 2324.000 1080.540 ;
        RECT 0.560 1076.060 2324.000 1079.380 ;
        RECT 1.420 1074.900 2324.000 1076.060 ;
        RECT 0.560 1071.580 2324.000 1074.900 ;
        RECT 1.420 1070.420 2324.000 1071.580 ;
        RECT 0.560 1067.100 2324.000 1070.420 ;
        RECT 1.420 1065.940 2324.000 1067.100 ;
        RECT 0.560 1062.620 2324.000 1065.940 ;
        RECT 1.420 1061.460 2324.000 1062.620 ;
        RECT 0.560 1058.140 2324.000 1061.460 ;
        RECT 1.420 1056.980 2324.000 1058.140 ;
        RECT 0.560 1053.660 2324.000 1056.980 ;
        RECT 1.420 1052.500 2324.000 1053.660 ;
        RECT 0.560 1049.180 2324.000 1052.500 ;
        RECT 1.420 1048.020 2324.000 1049.180 ;
        RECT 0.560 1044.700 2324.000 1048.020 ;
        RECT 1.420 1043.540 2324.000 1044.700 ;
        RECT 0.560 1040.220 2324.000 1043.540 ;
        RECT 1.420 1039.060 2324.000 1040.220 ;
        RECT 0.560 1035.740 2324.000 1039.060 ;
        RECT 1.420 1034.580 2324.000 1035.740 ;
        RECT 0.560 1031.260 2324.000 1034.580 ;
        RECT 1.420 1030.100 2324.000 1031.260 ;
        RECT 0.560 1026.780 2324.000 1030.100 ;
        RECT 1.420 1025.620 2324.000 1026.780 ;
        RECT 0.560 1022.300 2324.000 1025.620 ;
        RECT 1.420 1021.140 2324.000 1022.300 ;
        RECT 0.560 1017.820 2324.000 1021.140 ;
        RECT 1.420 1016.660 2324.000 1017.820 ;
        RECT 0.560 1013.340 2324.000 1016.660 ;
        RECT 1.420 1012.180 2324.000 1013.340 ;
        RECT 0.560 1008.860 2324.000 1012.180 ;
        RECT 1.420 1007.700 2324.000 1008.860 ;
        RECT 0.560 1004.380 2324.000 1007.700 ;
        RECT 1.420 1003.220 2324.000 1004.380 ;
        RECT 0.560 999.900 2324.000 1003.220 ;
        RECT 1.420 998.740 2324.000 999.900 ;
        RECT 0.560 995.420 2324.000 998.740 ;
        RECT 1.420 994.260 2324.000 995.420 ;
        RECT 0.560 990.940 2324.000 994.260 ;
        RECT 1.420 989.780 2324.000 990.940 ;
        RECT 0.560 986.460 2324.000 989.780 ;
        RECT 1.420 985.300 2324.000 986.460 ;
        RECT 0.560 981.980 2324.000 985.300 ;
        RECT 1.420 980.820 2324.000 981.980 ;
        RECT 0.560 977.500 2324.000 980.820 ;
        RECT 1.420 976.340 2324.000 977.500 ;
        RECT 0.560 973.020 2324.000 976.340 ;
        RECT 1.420 971.860 2324.000 973.020 ;
        RECT 0.560 968.540 2324.000 971.860 ;
        RECT 1.420 967.380 2324.000 968.540 ;
        RECT 0.560 964.060 2324.000 967.380 ;
        RECT 1.420 962.900 2324.000 964.060 ;
        RECT 0.560 959.580 2324.000 962.900 ;
        RECT 1.420 958.420 2324.000 959.580 ;
        RECT 0.560 955.100 2324.000 958.420 ;
        RECT 1.420 953.940 2324.000 955.100 ;
        RECT 0.560 950.620 2324.000 953.940 ;
        RECT 1.420 949.460 2324.000 950.620 ;
        RECT 0.560 927.660 2324.000 949.460 ;
        RECT 1.420 926.500 2324.000 927.660 ;
        RECT 0.560 923.180 2324.000 926.500 ;
        RECT 1.420 922.020 2324.000 923.180 ;
        RECT 0.560 918.700 2324.000 922.020 ;
        RECT 1.420 917.540 2324.000 918.700 ;
        RECT 0.560 914.220 2324.000 917.540 ;
        RECT 1.420 913.060 2324.000 914.220 ;
        RECT 0.560 909.740 2324.000 913.060 ;
        RECT 1.420 908.580 2324.000 909.740 ;
        RECT 0.560 905.260 2324.000 908.580 ;
        RECT 1.420 904.100 2324.000 905.260 ;
        RECT 0.560 900.780 2324.000 904.100 ;
        RECT 1.420 899.620 2324.000 900.780 ;
        RECT 0.560 896.300 2324.000 899.620 ;
        RECT 1.420 895.140 2324.000 896.300 ;
        RECT 0.560 891.820 2324.000 895.140 ;
        RECT 1.420 890.660 2324.000 891.820 ;
        RECT 0.560 887.340 2324.000 890.660 ;
        RECT 1.420 886.180 2324.000 887.340 ;
        RECT 0.560 882.860 2324.000 886.180 ;
        RECT 1.420 881.700 2324.000 882.860 ;
        RECT 0.560 878.380 2324.000 881.700 ;
        RECT 1.420 877.220 2324.000 878.380 ;
        RECT 0.560 873.900 2324.000 877.220 ;
        RECT 1.420 872.740 2324.000 873.900 ;
        RECT 0.560 869.420 2324.000 872.740 ;
        RECT 1.420 868.260 2324.000 869.420 ;
        RECT 0.560 864.940 2324.000 868.260 ;
        RECT 1.420 863.780 2324.000 864.940 ;
        RECT 0.560 860.460 2324.000 863.780 ;
        RECT 1.420 859.300 2324.000 860.460 ;
        RECT 0.560 855.980 2324.000 859.300 ;
        RECT 1.420 854.820 2324.000 855.980 ;
        RECT 0.560 851.500 2324.000 854.820 ;
        RECT 1.420 850.340 2324.000 851.500 ;
        RECT 0.560 847.020 2324.000 850.340 ;
        RECT 1.420 845.860 2324.000 847.020 ;
        RECT 0.560 842.540 2324.000 845.860 ;
        RECT 1.420 841.380 2324.000 842.540 ;
        RECT 0.560 838.060 2324.000 841.380 ;
        RECT 1.420 836.900 2324.000 838.060 ;
        RECT 0.560 833.580 2324.000 836.900 ;
        RECT 1.420 832.420 2324.000 833.580 ;
        RECT 0.560 829.100 2324.000 832.420 ;
        RECT 1.420 827.980 2324.000 829.100 ;
        RECT 1.420 827.940 2323.140 827.980 ;
        RECT 0.560 826.820 2323.140 827.940 ;
        RECT 0.560 824.620 2324.000 826.820 ;
        RECT 1.420 823.500 2324.000 824.620 ;
        RECT 1.420 823.460 2323.140 823.500 ;
        RECT 0.560 822.340 2323.140 823.460 ;
        RECT 0.560 820.140 2324.000 822.340 ;
        RECT 1.420 819.020 2324.000 820.140 ;
        RECT 1.420 818.980 2323.140 819.020 ;
        RECT 0.560 817.860 2323.140 818.980 ;
        RECT 0.560 815.660 2324.000 817.860 ;
        RECT 1.420 814.540 2324.000 815.660 ;
        RECT 1.420 814.500 2323.140 814.540 ;
        RECT 0.560 813.380 2323.140 814.500 ;
        RECT 0.560 811.180 2324.000 813.380 ;
        RECT 1.420 810.060 2324.000 811.180 ;
        RECT 1.420 810.020 2323.140 810.060 ;
        RECT 0.560 808.900 2323.140 810.020 ;
        RECT 0.560 806.700 2324.000 808.900 ;
        RECT 1.420 805.580 2324.000 806.700 ;
        RECT 1.420 805.540 2323.140 805.580 ;
        RECT 0.560 804.420 2323.140 805.540 ;
        RECT 0.560 802.220 2324.000 804.420 ;
        RECT 1.420 801.100 2324.000 802.220 ;
        RECT 1.420 801.060 2323.140 801.100 ;
        RECT 0.560 799.940 2323.140 801.060 ;
        RECT 0.560 797.740 2324.000 799.940 ;
        RECT 1.420 796.620 2324.000 797.740 ;
        RECT 1.420 796.580 2323.140 796.620 ;
        RECT 0.560 795.460 2323.140 796.580 ;
        RECT 0.560 793.260 2324.000 795.460 ;
        RECT 1.420 792.140 2324.000 793.260 ;
        RECT 1.420 792.100 2323.140 792.140 ;
        RECT 0.560 790.980 2323.140 792.100 ;
        RECT 0.560 788.780 2324.000 790.980 ;
        RECT 1.420 787.660 2324.000 788.780 ;
        RECT 1.420 787.620 2323.140 787.660 ;
        RECT 0.560 786.500 2323.140 787.620 ;
        RECT 0.560 784.300 2324.000 786.500 ;
        RECT 1.420 783.180 2324.000 784.300 ;
        RECT 1.420 783.140 2323.140 783.180 ;
        RECT 0.560 782.020 2323.140 783.140 ;
        RECT 0.560 779.820 2324.000 782.020 ;
        RECT 1.420 778.700 2324.000 779.820 ;
        RECT 1.420 778.660 2323.140 778.700 ;
        RECT 0.560 777.540 2323.140 778.660 ;
        RECT 0.560 775.340 2324.000 777.540 ;
        RECT 1.420 774.220 2324.000 775.340 ;
        RECT 1.420 774.180 2323.140 774.220 ;
        RECT 0.560 773.060 2323.140 774.180 ;
        RECT 0.560 770.860 2324.000 773.060 ;
        RECT 1.420 769.740 2324.000 770.860 ;
        RECT 1.420 769.700 2323.140 769.740 ;
        RECT 0.560 768.580 2323.140 769.700 ;
        RECT 0.560 766.380 2324.000 768.580 ;
        RECT 1.420 765.260 2324.000 766.380 ;
        RECT 1.420 765.220 2323.140 765.260 ;
        RECT 0.560 764.100 2323.140 765.220 ;
        RECT 0.560 761.900 2324.000 764.100 ;
        RECT 1.420 760.780 2324.000 761.900 ;
        RECT 1.420 760.740 2323.140 760.780 ;
        RECT 0.560 759.620 2323.140 760.740 ;
        RECT 0.560 757.420 2324.000 759.620 ;
        RECT 1.420 756.300 2324.000 757.420 ;
        RECT 1.420 756.260 2323.140 756.300 ;
        RECT 0.560 755.140 2323.140 756.260 ;
        RECT 0.560 752.940 2324.000 755.140 ;
        RECT 1.420 751.820 2324.000 752.940 ;
        RECT 1.420 751.780 2323.140 751.820 ;
        RECT 0.560 750.660 2323.140 751.780 ;
        RECT 0.560 748.460 2324.000 750.660 ;
        RECT 1.420 747.340 2324.000 748.460 ;
        RECT 1.420 747.300 2323.140 747.340 ;
        RECT 0.560 746.180 2323.140 747.300 ;
        RECT 0.560 743.980 2324.000 746.180 ;
        RECT 1.420 742.860 2324.000 743.980 ;
        RECT 1.420 742.820 2323.140 742.860 ;
        RECT 0.560 741.700 2323.140 742.820 ;
        RECT 0.560 739.500 2324.000 741.700 ;
        RECT 1.420 738.380 2324.000 739.500 ;
        RECT 1.420 738.340 2323.140 738.380 ;
        RECT 0.560 737.220 2323.140 738.340 ;
        RECT 0.560 735.020 2324.000 737.220 ;
        RECT 1.420 733.900 2324.000 735.020 ;
        RECT 1.420 733.860 2323.140 733.900 ;
        RECT 0.560 732.740 2323.140 733.860 ;
        RECT 0.560 730.540 2324.000 732.740 ;
        RECT 1.420 729.420 2324.000 730.540 ;
        RECT 1.420 729.380 2323.140 729.420 ;
        RECT 0.560 728.260 2323.140 729.380 ;
        RECT 0.560 726.060 2324.000 728.260 ;
        RECT 1.420 724.940 2324.000 726.060 ;
        RECT 1.420 724.900 2323.140 724.940 ;
        RECT 0.560 723.780 2323.140 724.900 ;
        RECT 0.560 721.580 2324.000 723.780 ;
        RECT 1.420 720.460 2324.000 721.580 ;
        RECT 1.420 720.420 2323.140 720.460 ;
        RECT 0.560 719.300 2323.140 720.420 ;
        RECT 0.560 717.100 2324.000 719.300 ;
        RECT 1.420 715.980 2324.000 717.100 ;
        RECT 1.420 715.940 2323.140 715.980 ;
        RECT 0.560 714.820 2323.140 715.940 ;
        RECT 0.560 712.620 2324.000 714.820 ;
        RECT 1.420 711.500 2324.000 712.620 ;
        RECT 1.420 711.460 2323.140 711.500 ;
        RECT 0.560 710.340 2323.140 711.460 ;
        RECT 0.560 708.140 2324.000 710.340 ;
        RECT 1.420 707.020 2324.000 708.140 ;
        RECT 1.420 706.980 2323.140 707.020 ;
        RECT 0.560 705.860 2323.140 706.980 ;
        RECT 0.560 703.660 2324.000 705.860 ;
        RECT 1.420 702.540 2324.000 703.660 ;
        RECT 1.420 702.500 2323.140 702.540 ;
        RECT 0.560 701.380 2323.140 702.500 ;
        RECT 0.560 699.180 2324.000 701.380 ;
        RECT 1.420 698.060 2324.000 699.180 ;
        RECT 1.420 698.020 2323.140 698.060 ;
        RECT 0.560 696.900 2323.140 698.020 ;
        RECT 0.560 694.700 2324.000 696.900 ;
        RECT 1.420 693.580 2324.000 694.700 ;
        RECT 1.420 693.540 2323.140 693.580 ;
        RECT 0.560 692.420 2323.140 693.540 ;
        RECT 0.560 690.220 2324.000 692.420 ;
        RECT 1.420 689.100 2324.000 690.220 ;
        RECT 1.420 689.060 2323.140 689.100 ;
        RECT 0.560 687.940 2323.140 689.060 ;
        RECT 0.560 685.740 2324.000 687.940 ;
        RECT 1.420 684.620 2324.000 685.740 ;
        RECT 1.420 684.580 2323.140 684.620 ;
        RECT 0.560 683.460 2323.140 684.580 ;
        RECT 0.560 681.260 2324.000 683.460 ;
        RECT 1.420 680.140 2324.000 681.260 ;
        RECT 1.420 680.100 2323.140 680.140 ;
        RECT 0.560 678.980 2323.140 680.100 ;
        RECT 0.560 676.780 2324.000 678.980 ;
        RECT 1.420 675.660 2324.000 676.780 ;
        RECT 1.420 675.620 2323.140 675.660 ;
        RECT 0.560 674.500 2323.140 675.620 ;
        RECT 0.560 672.300 2324.000 674.500 ;
        RECT 1.420 671.180 2324.000 672.300 ;
        RECT 1.420 671.140 2323.140 671.180 ;
        RECT 0.560 670.020 2323.140 671.140 ;
        RECT 0.560 667.820 2324.000 670.020 ;
        RECT 1.420 666.700 2324.000 667.820 ;
        RECT 1.420 666.660 2323.140 666.700 ;
        RECT 0.560 665.540 2323.140 666.660 ;
        RECT 0.560 663.340 2324.000 665.540 ;
        RECT 1.420 662.180 2324.000 663.340 ;
        RECT 0.560 640.380 2324.000 662.180 ;
        RECT 1.420 639.220 2324.000 640.380 ;
        RECT 0.560 635.900 2324.000 639.220 ;
        RECT 1.420 634.740 2324.000 635.900 ;
        RECT 0.560 631.420 2324.000 634.740 ;
        RECT 1.420 630.260 2324.000 631.420 ;
        RECT 0.560 626.940 2324.000 630.260 ;
        RECT 1.420 625.780 2324.000 626.940 ;
        RECT 0.560 622.460 2324.000 625.780 ;
        RECT 1.420 621.300 2324.000 622.460 ;
        RECT 0.560 617.980 2324.000 621.300 ;
        RECT 1.420 616.820 2324.000 617.980 ;
        RECT 0.560 613.500 2324.000 616.820 ;
        RECT 1.420 612.340 2324.000 613.500 ;
        RECT 0.560 609.020 2324.000 612.340 ;
        RECT 1.420 607.860 2324.000 609.020 ;
        RECT 0.560 604.540 2324.000 607.860 ;
        RECT 1.420 603.380 2324.000 604.540 ;
        RECT 0.560 600.060 2324.000 603.380 ;
        RECT 1.420 598.900 2324.000 600.060 ;
        RECT 0.560 595.580 2324.000 598.900 ;
        RECT 1.420 594.420 2324.000 595.580 ;
        RECT 0.560 591.100 2324.000 594.420 ;
        RECT 1.420 589.940 2324.000 591.100 ;
        RECT 0.560 586.620 2324.000 589.940 ;
        RECT 1.420 585.460 2324.000 586.620 ;
        RECT 0.560 582.140 2324.000 585.460 ;
        RECT 1.420 580.980 2324.000 582.140 ;
        RECT 0.560 577.660 2324.000 580.980 ;
        RECT 1.420 576.500 2324.000 577.660 ;
        RECT 0.560 573.180 2324.000 576.500 ;
        RECT 1.420 572.020 2324.000 573.180 ;
        RECT 0.560 568.700 2324.000 572.020 ;
        RECT 1.420 567.540 2324.000 568.700 ;
        RECT 0.560 564.220 2324.000 567.540 ;
        RECT 1.420 563.060 2324.000 564.220 ;
        RECT 0.560 559.740 2324.000 563.060 ;
        RECT 1.420 558.580 2324.000 559.740 ;
        RECT 0.560 555.260 2324.000 558.580 ;
        RECT 1.420 554.100 2324.000 555.260 ;
        RECT 0.560 550.780 2324.000 554.100 ;
        RECT 1.420 549.620 2324.000 550.780 ;
        RECT 0.560 546.300 2324.000 549.620 ;
        RECT 1.420 545.140 2324.000 546.300 ;
        RECT 0.560 541.820 2324.000 545.140 ;
        RECT 1.420 540.660 2324.000 541.820 ;
        RECT 0.560 537.340 2324.000 540.660 ;
        RECT 1.420 536.180 2324.000 537.340 ;
        RECT 0.560 532.860 2324.000 536.180 ;
        RECT 1.420 531.700 2324.000 532.860 ;
        RECT 0.560 528.380 2324.000 531.700 ;
        RECT 1.420 527.220 2324.000 528.380 ;
        RECT 0.560 523.900 2324.000 527.220 ;
        RECT 1.420 522.740 2324.000 523.900 ;
        RECT 0.560 519.420 2324.000 522.740 ;
        RECT 1.420 518.260 2324.000 519.420 ;
        RECT 0.560 514.940 2324.000 518.260 ;
        RECT 1.420 513.780 2324.000 514.940 ;
        RECT 0.560 510.460 2324.000 513.780 ;
        RECT 1.420 509.300 2324.000 510.460 ;
        RECT 0.560 505.980 2324.000 509.300 ;
        RECT 1.420 504.820 2324.000 505.980 ;
        RECT 0.560 501.500 2324.000 504.820 ;
        RECT 1.420 500.340 2324.000 501.500 ;
        RECT 0.560 497.020 2324.000 500.340 ;
        RECT 1.420 495.860 2324.000 497.020 ;
        RECT 0.560 492.540 2324.000 495.860 ;
        RECT 1.420 491.380 2324.000 492.540 ;
        RECT 0.560 488.060 2324.000 491.380 ;
        RECT 1.420 486.900 2324.000 488.060 ;
        RECT 0.560 483.580 2324.000 486.900 ;
        RECT 1.420 482.420 2324.000 483.580 ;
        RECT 0.560 479.100 2324.000 482.420 ;
        RECT 1.420 477.940 2324.000 479.100 ;
        RECT 0.560 474.620 2324.000 477.940 ;
        RECT 1.420 473.460 2324.000 474.620 ;
        RECT 0.560 470.140 2324.000 473.460 ;
        RECT 1.420 468.980 2324.000 470.140 ;
        RECT 0.560 465.660 2324.000 468.980 ;
        RECT 1.420 464.500 2324.000 465.660 ;
        RECT 0.560 461.180 2324.000 464.500 ;
        RECT 1.420 460.020 2324.000 461.180 ;
        RECT 0.560 456.700 2324.000 460.020 ;
        RECT 1.420 455.540 2324.000 456.700 ;
        RECT 0.560 452.220 2324.000 455.540 ;
        RECT 1.420 451.060 2324.000 452.220 ;
        RECT 0.560 447.740 2324.000 451.060 ;
        RECT 1.420 446.580 2324.000 447.740 ;
        RECT 0.560 443.260 2324.000 446.580 ;
        RECT 1.420 442.100 2324.000 443.260 ;
        RECT 0.560 438.780 2324.000 442.100 ;
        RECT 1.420 437.620 2324.000 438.780 ;
        RECT 0.560 434.300 2324.000 437.620 ;
        RECT 1.420 433.140 2324.000 434.300 ;
        RECT 0.560 429.820 2324.000 433.140 ;
        RECT 1.420 428.660 2324.000 429.820 ;
        RECT 0.560 425.340 2324.000 428.660 ;
        RECT 1.420 424.180 2324.000 425.340 ;
        RECT 0.560 420.860 2324.000 424.180 ;
        RECT 1.420 419.700 2324.000 420.860 ;
        RECT 0.560 416.380 2324.000 419.700 ;
        RECT 1.420 415.220 2324.000 416.380 ;
        RECT 0.560 411.900 2324.000 415.220 ;
        RECT 1.420 410.740 2324.000 411.900 ;
        RECT 0.560 407.420 2324.000 410.740 ;
        RECT 1.420 406.260 2324.000 407.420 ;
        RECT 0.560 402.940 2324.000 406.260 ;
        RECT 1.420 401.780 2324.000 402.940 ;
        RECT 0.560 398.460 2324.000 401.780 ;
        RECT 1.420 397.300 2324.000 398.460 ;
        RECT 0.560 393.980 2324.000 397.300 ;
        RECT 1.420 392.820 2324.000 393.980 ;
        RECT 0.560 389.500 2324.000 392.820 ;
        RECT 1.420 388.340 2324.000 389.500 ;
        RECT 0.560 385.020 2324.000 388.340 ;
        RECT 1.420 383.860 2324.000 385.020 ;
        RECT 0.560 380.540 2324.000 383.860 ;
        RECT 1.420 379.380 2324.000 380.540 ;
        RECT 0.560 376.060 2324.000 379.380 ;
        RECT 1.420 374.900 2324.000 376.060 ;
        RECT 0.560 353.100 2324.000 374.900 ;
        RECT 1.420 351.940 2324.000 353.100 ;
        RECT 0.560 348.620 2324.000 351.940 ;
        RECT 1.420 347.460 2324.000 348.620 ;
        RECT 0.560 344.140 2324.000 347.460 ;
        RECT 1.420 342.980 2324.000 344.140 ;
        RECT 0.560 339.660 2324.000 342.980 ;
        RECT 1.420 338.500 2324.000 339.660 ;
        RECT 0.560 335.180 2324.000 338.500 ;
        RECT 1.420 334.020 2324.000 335.180 ;
        RECT 0.560 330.700 2324.000 334.020 ;
        RECT 1.420 329.540 2324.000 330.700 ;
        RECT 0.560 326.220 2324.000 329.540 ;
        RECT 1.420 325.060 2324.000 326.220 ;
        RECT 0.560 321.740 2324.000 325.060 ;
        RECT 1.420 320.580 2324.000 321.740 ;
        RECT 0.560 317.260 2324.000 320.580 ;
        RECT 1.420 316.100 2324.000 317.260 ;
        RECT 0.560 312.780 2324.000 316.100 ;
        RECT 1.420 311.620 2324.000 312.780 ;
        RECT 0.560 308.300 2324.000 311.620 ;
        RECT 1.420 307.140 2324.000 308.300 ;
        RECT 0.560 303.820 2324.000 307.140 ;
        RECT 1.420 302.660 2324.000 303.820 ;
        RECT 0.560 299.340 2324.000 302.660 ;
        RECT 1.420 298.180 2324.000 299.340 ;
        RECT 0.560 294.860 2324.000 298.180 ;
        RECT 1.420 293.700 2324.000 294.860 ;
        RECT 0.560 290.380 2324.000 293.700 ;
        RECT 1.420 289.220 2324.000 290.380 ;
        RECT 0.560 285.900 2324.000 289.220 ;
        RECT 1.420 284.740 2324.000 285.900 ;
        RECT 0.560 281.420 2324.000 284.740 ;
        RECT 1.420 280.260 2324.000 281.420 ;
        RECT 0.560 276.940 2324.000 280.260 ;
        RECT 1.420 275.780 2324.000 276.940 ;
        RECT 0.560 272.460 2324.000 275.780 ;
        RECT 1.420 271.300 2324.000 272.460 ;
        RECT 0.560 267.980 2324.000 271.300 ;
        RECT 1.420 266.820 2324.000 267.980 ;
        RECT 0.560 263.500 2324.000 266.820 ;
        RECT 1.420 262.340 2324.000 263.500 ;
        RECT 0.560 259.020 2324.000 262.340 ;
        RECT 1.420 257.860 2324.000 259.020 ;
        RECT 0.560 254.540 2324.000 257.860 ;
        RECT 1.420 253.420 2324.000 254.540 ;
        RECT 1.420 253.380 2323.140 253.420 ;
        RECT 0.560 252.260 2323.140 253.380 ;
        RECT 0.560 250.060 2324.000 252.260 ;
        RECT 1.420 248.940 2324.000 250.060 ;
        RECT 1.420 248.900 2323.140 248.940 ;
        RECT 0.560 247.780 2323.140 248.900 ;
        RECT 0.560 245.580 2324.000 247.780 ;
        RECT 1.420 244.460 2324.000 245.580 ;
        RECT 1.420 244.420 2323.140 244.460 ;
        RECT 0.560 243.300 2323.140 244.420 ;
        RECT 0.560 241.100 2324.000 243.300 ;
        RECT 1.420 239.980 2324.000 241.100 ;
        RECT 1.420 239.940 2323.140 239.980 ;
        RECT 0.560 238.820 2323.140 239.940 ;
        RECT 0.560 236.620 2324.000 238.820 ;
        RECT 1.420 235.500 2324.000 236.620 ;
        RECT 1.420 235.460 2323.140 235.500 ;
        RECT 0.560 234.340 2323.140 235.460 ;
        RECT 0.560 232.140 2324.000 234.340 ;
        RECT 1.420 231.020 2324.000 232.140 ;
        RECT 1.420 230.980 2323.140 231.020 ;
        RECT 0.560 229.860 2323.140 230.980 ;
        RECT 0.560 227.660 2324.000 229.860 ;
        RECT 1.420 226.540 2324.000 227.660 ;
        RECT 1.420 226.500 2323.140 226.540 ;
        RECT 0.560 225.380 2323.140 226.500 ;
        RECT 0.560 223.180 2324.000 225.380 ;
        RECT 1.420 222.060 2324.000 223.180 ;
        RECT 1.420 222.020 2323.140 222.060 ;
        RECT 0.560 220.900 2323.140 222.020 ;
        RECT 0.560 218.700 2324.000 220.900 ;
        RECT 1.420 217.580 2324.000 218.700 ;
        RECT 1.420 217.540 2323.140 217.580 ;
        RECT 0.560 216.420 2323.140 217.540 ;
        RECT 0.560 214.220 2324.000 216.420 ;
        RECT 1.420 213.100 2324.000 214.220 ;
        RECT 1.420 213.060 2323.140 213.100 ;
        RECT 0.560 211.940 2323.140 213.060 ;
        RECT 0.560 209.740 2324.000 211.940 ;
        RECT 1.420 208.620 2324.000 209.740 ;
        RECT 1.420 208.580 2323.140 208.620 ;
        RECT 0.560 207.460 2323.140 208.580 ;
        RECT 0.560 205.260 2324.000 207.460 ;
        RECT 1.420 204.140 2324.000 205.260 ;
        RECT 1.420 204.100 2323.140 204.140 ;
        RECT 0.560 202.980 2323.140 204.100 ;
        RECT 0.560 200.780 2324.000 202.980 ;
        RECT 1.420 199.660 2324.000 200.780 ;
        RECT 1.420 199.620 2323.140 199.660 ;
        RECT 0.560 198.500 2323.140 199.620 ;
        RECT 0.560 196.300 2324.000 198.500 ;
        RECT 1.420 195.180 2324.000 196.300 ;
        RECT 1.420 195.140 2323.140 195.180 ;
        RECT 0.560 194.020 2323.140 195.140 ;
        RECT 0.560 191.820 2324.000 194.020 ;
        RECT 1.420 190.700 2324.000 191.820 ;
        RECT 1.420 190.660 2323.140 190.700 ;
        RECT 0.560 189.540 2323.140 190.660 ;
        RECT 0.560 187.340 2324.000 189.540 ;
        RECT 1.420 186.220 2324.000 187.340 ;
        RECT 1.420 186.180 2323.140 186.220 ;
        RECT 0.560 185.060 2323.140 186.180 ;
        RECT 0.560 182.860 2324.000 185.060 ;
        RECT 1.420 181.740 2324.000 182.860 ;
        RECT 1.420 181.700 2323.140 181.740 ;
        RECT 0.560 180.580 2323.140 181.700 ;
        RECT 0.560 178.380 2324.000 180.580 ;
        RECT 1.420 177.260 2324.000 178.380 ;
        RECT 1.420 177.220 2323.140 177.260 ;
        RECT 0.560 176.100 2323.140 177.220 ;
        RECT 0.560 173.900 2324.000 176.100 ;
        RECT 1.420 172.780 2324.000 173.900 ;
        RECT 1.420 172.740 2323.140 172.780 ;
        RECT 0.560 171.620 2323.140 172.740 ;
        RECT 0.560 169.420 2324.000 171.620 ;
        RECT 1.420 168.300 2324.000 169.420 ;
        RECT 1.420 168.260 2323.140 168.300 ;
        RECT 0.560 167.140 2323.140 168.260 ;
        RECT 0.560 164.940 2324.000 167.140 ;
        RECT 1.420 163.820 2324.000 164.940 ;
        RECT 1.420 163.780 2323.140 163.820 ;
        RECT 0.560 162.660 2323.140 163.780 ;
        RECT 0.560 160.460 2324.000 162.660 ;
        RECT 1.420 159.340 2324.000 160.460 ;
        RECT 1.420 159.300 2323.140 159.340 ;
        RECT 0.560 158.180 2323.140 159.300 ;
        RECT 0.560 155.980 2324.000 158.180 ;
        RECT 1.420 154.860 2324.000 155.980 ;
        RECT 1.420 154.820 2323.140 154.860 ;
        RECT 0.560 153.700 2323.140 154.820 ;
        RECT 0.560 151.500 2324.000 153.700 ;
        RECT 1.420 150.380 2324.000 151.500 ;
        RECT 1.420 150.340 2323.140 150.380 ;
        RECT 0.560 149.220 2323.140 150.340 ;
        RECT 0.560 147.020 2324.000 149.220 ;
        RECT 1.420 145.900 2324.000 147.020 ;
        RECT 1.420 145.860 2323.140 145.900 ;
        RECT 0.560 144.740 2323.140 145.860 ;
        RECT 0.560 142.540 2324.000 144.740 ;
        RECT 1.420 141.420 2324.000 142.540 ;
        RECT 1.420 141.380 2323.140 141.420 ;
        RECT 0.560 140.260 2323.140 141.380 ;
        RECT 0.560 138.060 2324.000 140.260 ;
        RECT 1.420 136.940 2324.000 138.060 ;
        RECT 1.420 136.900 2323.140 136.940 ;
        RECT 0.560 135.780 2323.140 136.900 ;
        RECT 0.560 133.580 2324.000 135.780 ;
        RECT 1.420 132.460 2324.000 133.580 ;
        RECT 1.420 132.420 2323.140 132.460 ;
        RECT 0.560 131.300 2323.140 132.420 ;
        RECT 0.560 129.100 2324.000 131.300 ;
        RECT 1.420 127.980 2324.000 129.100 ;
        RECT 1.420 127.940 2323.140 127.980 ;
        RECT 0.560 126.820 2323.140 127.940 ;
        RECT 0.560 124.620 2324.000 126.820 ;
        RECT 1.420 123.500 2324.000 124.620 ;
        RECT 1.420 123.460 2323.140 123.500 ;
        RECT 0.560 122.340 2323.140 123.460 ;
        RECT 0.560 120.140 2324.000 122.340 ;
        RECT 1.420 119.020 2324.000 120.140 ;
        RECT 1.420 118.980 2323.140 119.020 ;
        RECT 0.560 117.860 2323.140 118.980 ;
        RECT 0.560 115.660 2324.000 117.860 ;
        RECT 1.420 114.540 2324.000 115.660 ;
        RECT 1.420 114.500 2323.140 114.540 ;
        RECT 0.560 113.380 2323.140 114.500 ;
        RECT 0.560 111.180 2324.000 113.380 ;
        RECT 1.420 110.060 2324.000 111.180 ;
        RECT 1.420 110.020 2323.140 110.060 ;
        RECT 0.560 108.900 2323.140 110.020 ;
        RECT 0.560 106.700 2324.000 108.900 ;
        RECT 1.420 105.580 2324.000 106.700 ;
        RECT 1.420 105.540 2323.140 105.580 ;
        RECT 0.560 104.420 2323.140 105.540 ;
        RECT 0.560 102.220 2324.000 104.420 ;
        RECT 1.420 101.100 2324.000 102.220 ;
        RECT 1.420 101.060 2323.140 101.100 ;
        RECT 0.560 99.940 2323.140 101.060 ;
        RECT 0.560 97.740 2324.000 99.940 ;
        RECT 1.420 96.620 2324.000 97.740 ;
        RECT 1.420 96.580 2323.140 96.620 ;
        RECT 0.560 95.460 2323.140 96.580 ;
        RECT 0.560 93.260 2324.000 95.460 ;
        RECT 1.420 92.140 2324.000 93.260 ;
        RECT 1.420 92.100 2323.140 92.140 ;
        RECT 0.560 90.980 2323.140 92.100 ;
        RECT 0.560 88.780 2324.000 90.980 ;
        RECT 1.420 87.620 2324.000 88.780 ;
        RECT 0.560 75.900 2324.000 87.620 ;
        RECT 0.860 74.740 2324.000 75.900 ;
        RECT 0.560 73.660 2324.000 74.740 ;
        RECT 0.860 72.500 2324.000 73.660 ;
        RECT 0.560 71.420 2324.000 72.500 ;
        RECT 0.860 70.260 2324.000 71.420 ;
        RECT 0.560 69.180 2324.000 70.260 ;
        RECT 0.860 68.020 2324.000 69.180 ;
        RECT 0.560 66.940 2324.000 68.020 ;
        RECT 0.860 65.780 2324.000 66.940 ;
        RECT 0.560 64.700 2324.000 65.780 ;
        RECT 0.860 63.540 2324.000 64.700 ;
        RECT 0.560 62.460 2324.000 63.540 ;
        RECT 0.860 61.300 2324.000 62.460 ;
        RECT 0.560 60.220 2324.000 61.300 ;
        RECT 0.860 59.060 2324.000 60.220 ;
        RECT 0.560 57.980 2324.000 59.060 ;
        RECT 0.860 56.820 2324.000 57.980 ;
        RECT 0.560 55.740 2324.000 56.820 ;
        RECT 0.860 54.580 2324.000 55.740 ;
        RECT 0.560 53.500 2324.000 54.580 ;
        RECT 0.860 52.340 2324.000 53.500 ;
        RECT 0.560 51.260 2324.000 52.340 ;
        RECT 0.860 50.100 2324.000 51.260 ;
        RECT 0.560 49.020 2324.000 50.100 ;
        RECT 0.860 47.860 2324.000 49.020 ;
        RECT 0.560 46.780 2324.000 47.860 ;
        RECT 0.860 45.620 2324.000 46.780 ;
        RECT 0.560 44.540 2324.000 45.620 ;
        RECT 0.860 43.380 2324.000 44.540 ;
        RECT 0.560 42.300 2324.000 43.380 ;
        RECT 0.860 41.140 2324.000 42.300 ;
        RECT 0.560 40.060 2324.000 41.140 ;
        RECT 0.860 38.900 2324.000 40.060 ;
        RECT 0.560 37.820 2324.000 38.900 ;
        RECT 0.860 36.660 2324.000 37.820 ;
        RECT 0.560 35.580 2324.000 36.660 ;
        RECT 0.860 34.420 2324.000 35.580 ;
        RECT 0.560 33.340 2324.000 34.420 ;
        RECT 0.860 32.180 2324.000 33.340 ;
        RECT 0.560 31.100 2324.000 32.180 ;
        RECT 0.860 29.940 2324.000 31.100 ;
        RECT 0.560 28.860 2324.000 29.940 ;
        RECT 0.860 27.700 2324.000 28.860 ;
        RECT 0.560 26.620 2324.000 27.700 ;
        RECT 0.860 25.460 2324.000 26.620 ;
        RECT 0.560 24.380 2324.000 25.460 ;
        RECT 0.860 23.220 2324.000 24.380 ;
        RECT 0.560 22.140 2324.000 23.220 ;
        RECT 0.860 20.980 2324.000 22.140 ;
        RECT 0.560 19.900 2324.000 20.980 ;
        RECT 0.860 18.740 2324.000 19.900 ;
        RECT 0.560 17.660 2324.000 18.740 ;
        RECT 0.860 16.500 2324.000 17.660 ;
        RECT 0.560 15.420 2324.000 16.500 ;
        RECT 0.860 14.260 2324.000 15.420 ;
        RECT 0.560 13.180 2324.000 14.260 ;
        RECT 0.860 12.020 2324.000 13.180 ;
        RECT 0.560 10.940 2324.000 12.020 ;
        RECT 0.860 9.780 2324.000 10.940 ;
        RECT 0.560 8.700 2324.000 9.780 ;
        RECT 0.860 7.540 2324.000 8.700 ;
        RECT 0.560 6.460 2324.000 7.540 ;
        RECT 0.860 5.300 2324.000 6.460 ;
        RECT 0.560 0.140 2324.000 5.300 ;
      LAYER Metal4 ;
        RECT 9.660 3595.500 2308.740 3595.670 ;
        RECT 9.660 3524.380 161.940 3595.500 ;
        RECT 9.660 76.420 19.140 3524.380 ;
        RECT 21.340 76.420 22.440 3524.380 ;
        RECT 24.640 76.420 119.140 3524.380 ;
        RECT 121.340 76.420 122.440 3524.380 ;
        RECT 124.640 76.420 161.940 3524.380 ;
        RECT 9.660 5.690 161.940 76.420 ;
        RECT 164.140 5.690 165.240 3595.500 ;
        RECT 167.440 5.690 261.940 3595.500 ;
        RECT 264.140 5.690 265.240 3595.500 ;
        RECT 267.440 5.690 361.940 3595.500 ;
        RECT 364.140 5.690 365.240 3595.500 ;
        RECT 367.440 5.690 449.220 3595.500 ;
        RECT 451.420 5.690 452.520 3595.500 ;
        RECT 454.720 5.690 549.220 3595.500 ;
        RECT 551.420 5.690 552.520 3595.500 ;
        RECT 554.720 5.690 649.220 3595.500 ;
        RECT 651.420 5.690 652.520 3595.500 ;
        RECT 654.720 5.690 736.500 3595.500 ;
        RECT 738.700 5.690 739.800 3595.500 ;
        RECT 742.000 5.690 836.500 3595.500 ;
        RECT 838.700 5.690 839.800 3595.500 ;
        RECT 842.000 5.690 936.500 3595.500 ;
        RECT 938.700 5.690 939.800 3595.500 ;
        RECT 942.000 5.690 1023.780 3595.500 ;
        RECT 1025.980 5.690 1027.080 3595.500 ;
        RECT 1029.280 5.690 1123.780 3595.500 ;
        RECT 1125.980 5.690 1127.080 3595.500 ;
        RECT 1129.280 5.690 1223.780 3595.500 ;
        RECT 1225.980 5.690 1227.080 3595.500 ;
        RECT 1229.280 5.690 1345.780 3595.500 ;
        RECT 1347.980 5.690 1349.080 3595.500 ;
        RECT 1351.280 5.690 1445.780 3595.500 ;
        RECT 1447.980 5.690 1449.080 3595.500 ;
        RECT 1451.280 5.690 1545.780 3595.500 ;
        RECT 1547.980 5.690 1549.080 3595.500 ;
        RECT 1551.280 5.690 1633.060 3595.500 ;
        RECT 1635.260 5.690 1636.360 3595.500 ;
        RECT 1638.560 5.690 1733.060 3595.500 ;
        RECT 1735.260 5.690 1736.360 3595.500 ;
        RECT 1738.560 5.690 1833.060 3595.500 ;
        RECT 1835.260 5.690 1836.360 3595.500 ;
        RECT 1838.560 5.690 1896.820 3595.500 ;
        RECT 1899.020 5.690 1900.120 3595.500 ;
        RECT 1902.320 5.690 1996.820 3595.500 ;
        RECT 1999.020 5.690 2000.120 3595.500 ;
        RECT 2002.320 5.690 2096.820 3595.500 ;
        RECT 2099.020 5.690 2100.120 3595.500 ;
        RECT 2102.320 5.690 2184.100 3595.500 ;
        RECT 2186.300 5.690 2187.400 3595.500 ;
        RECT 2189.600 5.690 2284.100 3595.500 ;
        RECT 2286.300 5.690 2287.400 3595.500 ;
        RECT 2289.600 5.690 2308.740 3595.500 ;
  END
END eFPGA
END LIBRARY

