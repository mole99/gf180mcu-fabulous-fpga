* NGSPICE file created from S_term_single2.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

.subckt S_term_single2 FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0]
+ N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10]
+ N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4]
+ N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12]
+ NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5]
+ NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3] S2END[0]
+ S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1]
+ S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VDD VSS
XFILLER_10_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_9_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_505 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_527 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_11_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_062_ S2MID[1] net63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_438 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_045_ FrameStrobe[13] net37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_444 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_028_ FrameData[28] net21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput53 net53 N1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput42 net42 FrameStrobe_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput97 net97 NN4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput75 net75 N4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput86 net86 N4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput64 net64 N2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput20 net20 FrameData_O[27] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput7 net7 FrameData_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_2_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput31 net31 FrameData_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_9_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_12_Right_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_061_ S2MID[2] net62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_9_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_044_ FrameStrobe[12] net36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_15_560 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_478 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_027_ FrameData[27] net20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_6_Right_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput87 net87 N4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput65 net65 N2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput54 net54 N1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput43 net43 FrameStrobe_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput98 net98 NN4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput76 net76 N4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput21 net21 FrameData_O[28] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput10 net10 FrameData_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput8 net8 FrameData_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_2_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput32 net32 FrameData_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_10_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_060_ S2MID[3] net61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_043_ FrameStrobe[11] net35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_487 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_531 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_026_ FrameData[26] net19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_6_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput33 net33 FrameStrobe_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput99 net99 NN4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput44 net44 FrameStrobe_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput88 net88 N4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput77 net77 N4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput55 net55 N1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput22 net22 FrameData_O[29] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput66 net66 N2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput11 net11 FrameData_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput9 net9 FrameData_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_2_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_009_ FrameData[9] net32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_9_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_408 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_540 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_12_Left_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_042_ FrameStrobe[10] net34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_025_ FrameData[25] net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput34 net34 FrameStrobe_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput78 net78 N4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput56 net56 N1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput67 net67 N2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput45 net45 FrameStrobe_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput89 net89 NN4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput12 net12 FrameData_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput23 net23 FrameData_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_5_517 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_008_ FrameData[8] net31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_15_Left_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_9_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_0_Left_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_041_ FrameStrobe[9] net52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_024_ FrameData[24] net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_6_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput46 net46 FrameStrobe_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput57 net57 N2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput13 net13 FrameData_O[20] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput35 net35 FrameStrobe_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_5_507 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput24 net24 FrameData_O[30] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput79 net79 N4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput68 net68 N2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_8_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_007_ FrameData[7] net30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_14_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_494 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_461 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_472 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_450 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_443 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_040_ FrameStrobe[8] net51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_479 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_023_ FrameData[23] net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_8_527 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_505 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput47 net47 FrameStrobe_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput36 net36 FrameStrobe_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput69 net69 N2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput14 net14 FrameData_O[21] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput25 net25 FrameData_O[31] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput58 net58 N2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_006_ FrameData[6] net29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_8_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_500 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_522 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_385 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_447 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_099_ SS4END[4] net91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_022_ FrameData[22] net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_6_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput37 net37 FrameStrobe_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput59 net59 N2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput48 net48 FrameStrobe_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput15 net15 FrameData_O[22] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_12_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Right_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput26 net26 FrameData_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_7_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_005_ FrameData[5] net28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_4_531 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_460 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_486 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_098_ SS4END[5] net90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_021_ FrameData[21] net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_7_Left_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_6_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput49 net49 FrameStrobe_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput16 net16 FrameData_O[23] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput38 net38 FrameStrobe_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput27 net27 FrameData_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_12_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_004_ FrameData[4] net27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_4_521 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_15_Right_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_442 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_438 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_097_ SS4END[6] net104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_020_ FrameData[20] net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_15_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput39 net39 FrameStrobe_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput17 net17 FrameData_O[24] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput28 net28 FrameData_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_8_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_003_ FrameData[3] net26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_15_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_096_ SS4END[7] net103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_527 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput18 net18 FrameData_O[25] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput29 net29 FrameData_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_079_ S4END[8] net86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_8_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_002_ FrameData[2] net23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_5_Right_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_3_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_488 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_095_ SS4END[8] net102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_078_ S4END[9] net85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput19 net19 FrameData_O[26] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_001_ FrameData[1] net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_4_513 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_11_Right_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_13_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_427 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_482 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_094_ SS4END[9] net101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_11_Left_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_077_ S4END[10] net84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_6_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_000_ FrameData[0] net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_8_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Left_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_336 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_450 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_093_ SS4END[10] net100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_497 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_512 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_076_ S4END[11] net83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_6_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_059_ S2MID[4] net60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_12_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_518 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Right_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_400 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_506 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_092_ SS4END[11] net99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_2_465 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_075_ S4END[12] net82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_12_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_527 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_058_ S2MID[5] net59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_8_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_3_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_316 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_415 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_426 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_091_ SS4END[12] net98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_514 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_074_ S4END[13] net81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_2_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_057_ S2MID[6] net58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_8_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_0_Right_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Left_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_090_ SS4END[13] net97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_500 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_073_ S4END[14] net80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_056_ S2MID[7] net57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_6_Left_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_039_ FrameStrobe[7] net50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_13_458 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_072_ S4END[15] net73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_055_ S1END[0] net56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_038_ FrameStrobe[6] net49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_13_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_481 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Right_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_502 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_071_ S2END[0] net72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_14_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_054_ S1END[1] net55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_520 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_13_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_037_ FrameStrobe[5] net48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_7_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_512 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_4_Right_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_10_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_4_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_555 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_070_ S2END[1] net71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_15_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_053_ S1END[2] net54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_546 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_036_ FrameStrobe[4] net47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_019_ FrameData[19] net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_4_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_482 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_508 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_316 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_522 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_052_ S1END[3] net53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_10_Left_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_7_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_035_ FrameStrobe[3] net46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_13_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_104_ UserCLK net105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_473 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_018_ FrameData[18] net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_4_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_513 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_524 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_450 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_531 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_10_Right_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_051_ FrameStrobe[19] net43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_7_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_103_ SS4END[0] net95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_034_ FrameStrobe[2] net45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_13_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_397 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Right_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_4_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_017_ FrameData[17] net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_1_440 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput100 net100 NN4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_050_ FrameStrobe[18] net42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_14_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_033_ FrameStrobe[1] net44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_102_ SS4END[1] net94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_016_ FrameData[16] net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_8_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_4_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_438 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_559 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_515 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput101 net101 NN4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_7_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_032_ FrameStrobe[0] net33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_101_ SS4END[2] net93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_388 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_015_ FrameData[15] net7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_4_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_450 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_2_Left_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput102 net102 NN4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_7_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_031_ FrameData[31] net25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_100_ SS4END[3] net92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_12_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_5_Left_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_014_ FrameData[14] net6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_4_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_531 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_513 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput103 net103 NN4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_11_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_516 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_475 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_030_ FrameData[30] net24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_8_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_013_ FrameData[13] net5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_4_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_500 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput104 net104 NN4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_9_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_089_ SS4END[14] net96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_12_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_483 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_012_ FrameData[12] net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_3_Right_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_497 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput105 net105 UserCLKo VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_15_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_444 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_088_ SS4END[15] net89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_9_Left_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_011_ FrameData[11] net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_13_Right_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_527 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_353 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_508 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_467 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_087_ S4END[0] net79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_8_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_010_ FrameData[10] net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_388 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_2_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_531 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_446 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_086_ S4END[1] net78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_069_ S2END[2] net70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_442 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_423 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_434 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_7_Right_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput90 net90 NN4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_13_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_2_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_12_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_085_ S4END[2] net77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_487 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_068_ S2END[3] net69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_12_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_5_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_556 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput1 net1 FrameData_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput91 net91 NN4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput80 net80 N4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_10_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_15_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_084_ S4END[3] net76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_400 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_13_Left_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_067_ S2END[4] net68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_2_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_425 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_527 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput70 net70 N2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput92 net92 NN4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput81 net81 N4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_2_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput2 net2 FrameData_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_14_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_1_Left_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_15_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_361 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_083_ S4END[4] net75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_5_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Left_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_066_ S2END[5] net67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_049_ FrameStrobe[17] net41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_5_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput93 net93 NN4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput60 net60 N2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput82 net82 N4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput71 net71 N2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput3 net3 FrameData_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_5_521 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_082_ S4END[5] net74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_12_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_486 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_065_ S2END[6] net66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_048_ FrameStrobe[16] net40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_1_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput50 net50 FrameStrobe_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput94 net94 NN4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput83 net83 N4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput72 net72 N2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput61 net61 N2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput4 net4 FrameData_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_13_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_374 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_081_ S4END[6] net88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_14_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_064_ S2END[7] net65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_047_ FrameStrobe[15] net39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_5_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_2_Right_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_531 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput95 net95 NN4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput73 net73 N4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput51 net51 FrameStrobe_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput40 net40 FrameStrobe_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_13_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput62 net62 N2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput84 net84 N4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput5 net5 FrameData_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_10_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_080_ S4END[7] net87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_11_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_063_ S2MID[0] net64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_9_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_8_Left_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_046_ FrameStrobe[14] net38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_029_ FrameData[29] net22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput41 net41 FrameStrobe_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput52 net52 FrameStrobe_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_2_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput30 net30 FrameData_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput6 net6 FrameData_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput96 net96 NN4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput63 net63 N2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput85 net85 N4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput74 net74 N4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_8_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
.ends

