* NGSPICE file created from DSP.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latq_1 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

.subckt DSP Tile_X0Y0_E1BEG[0] Tile_X0Y0_E1BEG[1] Tile_X0Y0_E1BEG[2] Tile_X0Y0_E1BEG[3]
+ Tile_X0Y0_E1END[0] Tile_X0Y0_E1END[1] Tile_X0Y0_E1END[2] Tile_X0Y0_E1END[3] Tile_X0Y0_E2BEG[0]
+ Tile_X0Y0_E2BEG[1] Tile_X0Y0_E2BEG[2] Tile_X0Y0_E2BEG[3] Tile_X0Y0_E2BEG[4] Tile_X0Y0_E2BEG[5]
+ Tile_X0Y0_E2BEG[6] Tile_X0Y0_E2BEG[7] Tile_X0Y0_E2BEGb[0] Tile_X0Y0_E2BEGb[1] Tile_X0Y0_E2BEGb[2]
+ Tile_X0Y0_E2BEGb[3] Tile_X0Y0_E2BEGb[4] Tile_X0Y0_E2BEGb[5] Tile_X0Y0_E2BEGb[6]
+ Tile_X0Y0_E2BEGb[7] Tile_X0Y0_E2END[0] Tile_X0Y0_E2END[1] Tile_X0Y0_E2END[2] Tile_X0Y0_E2END[3]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_E2END[5] Tile_X0Y0_E2END[6] Tile_X0Y0_E2END[7] Tile_X0Y0_E2MID[0]
+ Tile_X0Y0_E2MID[1] Tile_X0Y0_E2MID[2] Tile_X0Y0_E2MID[3] Tile_X0Y0_E2MID[4] Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_E2MID[6] Tile_X0Y0_E2MID[7] Tile_X0Y0_E6BEG[0] Tile_X0Y0_E6BEG[10] Tile_X0Y0_E6BEG[11]
+ Tile_X0Y0_E6BEG[1] Tile_X0Y0_E6BEG[2] Tile_X0Y0_E6BEG[3] Tile_X0Y0_E6BEG[4] Tile_X0Y0_E6BEG[5]
+ Tile_X0Y0_E6BEG[6] Tile_X0Y0_E6BEG[7] Tile_X0Y0_E6BEG[8] Tile_X0Y0_E6BEG[9] Tile_X0Y0_E6END[0]
+ Tile_X0Y0_E6END[10] Tile_X0Y0_E6END[11] Tile_X0Y0_E6END[1] Tile_X0Y0_E6END[2] Tile_X0Y0_E6END[3]
+ Tile_X0Y0_E6END[4] Tile_X0Y0_E6END[5] Tile_X0Y0_E6END[6] Tile_X0Y0_E6END[7] Tile_X0Y0_E6END[8]
+ Tile_X0Y0_E6END[9] Tile_X0Y0_EE4BEG[0] Tile_X0Y0_EE4BEG[10] Tile_X0Y0_EE4BEG[11]
+ Tile_X0Y0_EE4BEG[12] Tile_X0Y0_EE4BEG[13] Tile_X0Y0_EE4BEG[14] Tile_X0Y0_EE4BEG[15]
+ Tile_X0Y0_EE4BEG[1] Tile_X0Y0_EE4BEG[2] Tile_X0Y0_EE4BEG[3] Tile_X0Y0_EE4BEG[4]
+ Tile_X0Y0_EE4BEG[5] Tile_X0Y0_EE4BEG[6] Tile_X0Y0_EE4BEG[7] Tile_X0Y0_EE4BEG[8]
+ Tile_X0Y0_EE4BEG[9] Tile_X0Y0_EE4END[0] Tile_X0Y0_EE4END[10] Tile_X0Y0_EE4END[11]
+ Tile_X0Y0_EE4END[12] Tile_X0Y0_EE4END[13] Tile_X0Y0_EE4END[14] Tile_X0Y0_EE4END[15]
+ Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[2] Tile_X0Y0_EE4END[3] Tile_X0Y0_EE4END[4]
+ Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[6] Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[8]
+ Tile_X0Y0_EE4END[9] Tile_X0Y0_FrameData[0] Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData[11]
+ Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData[13] Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData[15]
+ Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData[17] Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData[19]
+ Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData[20] Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData[22]
+ Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData[24] Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData[26]
+ Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData[28] Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData[2]
+ Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData[31] Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData[4]
+ Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData[6] Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData[8]
+ Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[0] Tile_X0Y0_FrameData_O[10] Tile_X0Y0_FrameData_O[11]
+ Tile_X0Y0_FrameData_O[12] Tile_X0Y0_FrameData_O[13] Tile_X0Y0_FrameData_O[14] Tile_X0Y0_FrameData_O[15]
+ Tile_X0Y0_FrameData_O[16] Tile_X0Y0_FrameData_O[17] Tile_X0Y0_FrameData_O[18] Tile_X0Y0_FrameData_O[19]
+ Tile_X0Y0_FrameData_O[1] Tile_X0Y0_FrameData_O[20] Tile_X0Y0_FrameData_O[21] Tile_X0Y0_FrameData_O[22]
+ Tile_X0Y0_FrameData_O[23] Tile_X0Y0_FrameData_O[24] Tile_X0Y0_FrameData_O[25] Tile_X0Y0_FrameData_O[26]
+ Tile_X0Y0_FrameData_O[27] Tile_X0Y0_FrameData_O[28] Tile_X0Y0_FrameData_O[29] Tile_X0Y0_FrameData_O[2]
+ Tile_X0Y0_FrameData_O[30] Tile_X0Y0_FrameData_O[31] Tile_X0Y0_FrameData_O[3] Tile_X0Y0_FrameData_O[4]
+ Tile_X0Y0_FrameData_O[5] Tile_X0Y0_FrameData_O[6] Tile_X0Y0_FrameData_O[7] Tile_X0Y0_FrameData_O[8]
+ Tile_X0Y0_FrameData_O[9] Tile_X0Y0_FrameStrobe_O[0] Tile_X0Y0_FrameStrobe_O[10]
+ Tile_X0Y0_FrameStrobe_O[11] Tile_X0Y0_FrameStrobe_O[12] Tile_X0Y0_FrameStrobe_O[13]
+ Tile_X0Y0_FrameStrobe_O[14] Tile_X0Y0_FrameStrobe_O[15] Tile_X0Y0_FrameStrobe_O[16]
+ Tile_X0Y0_FrameStrobe_O[17] Tile_X0Y0_FrameStrobe_O[18] Tile_X0Y0_FrameStrobe_O[19]
+ Tile_X0Y0_FrameStrobe_O[1] Tile_X0Y0_FrameStrobe_O[2] Tile_X0Y0_FrameStrobe_O[3]
+ Tile_X0Y0_FrameStrobe_O[4] Tile_X0Y0_FrameStrobe_O[5] Tile_X0Y0_FrameStrobe_O[6]
+ Tile_X0Y0_FrameStrobe_O[7] Tile_X0Y0_FrameStrobe_O[8] Tile_X0Y0_FrameStrobe_O[9]
+ Tile_X0Y0_N1BEG[0] Tile_X0Y0_N1BEG[1] Tile_X0Y0_N1BEG[2] Tile_X0Y0_N1BEG[3] Tile_X0Y0_N2BEG[0]
+ Tile_X0Y0_N2BEG[1] Tile_X0Y0_N2BEG[2] Tile_X0Y0_N2BEG[3] Tile_X0Y0_N2BEG[4] Tile_X0Y0_N2BEG[5]
+ Tile_X0Y0_N2BEG[6] Tile_X0Y0_N2BEG[7] Tile_X0Y0_N2BEGb[0] Tile_X0Y0_N2BEGb[1] Tile_X0Y0_N2BEGb[2]
+ Tile_X0Y0_N2BEGb[3] Tile_X0Y0_N2BEGb[4] Tile_X0Y0_N2BEGb[5] Tile_X0Y0_N2BEGb[6]
+ Tile_X0Y0_N2BEGb[7] Tile_X0Y0_N4BEG[0] Tile_X0Y0_N4BEG[10] Tile_X0Y0_N4BEG[11] Tile_X0Y0_N4BEG[12]
+ Tile_X0Y0_N4BEG[13] Tile_X0Y0_N4BEG[14] Tile_X0Y0_N4BEG[15] Tile_X0Y0_N4BEG[1] Tile_X0Y0_N4BEG[2]
+ Tile_X0Y0_N4BEG[3] Tile_X0Y0_N4BEG[4] Tile_X0Y0_N4BEG[5] Tile_X0Y0_N4BEG[6] Tile_X0Y0_N4BEG[7]
+ Tile_X0Y0_N4BEG[8] Tile_X0Y0_N4BEG[9] Tile_X0Y0_NN4BEG[0] Tile_X0Y0_NN4BEG[10] Tile_X0Y0_NN4BEG[11]
+ Tile_X0Y0_NN4BEG[12] Tile_X0Y0_NN4BEG[13] Tile_X0Y0_NN4BEG[14] Tile_X0Y0_NN4BEG[15]
+ Tile_X0Y0_NN4BEG[1] Tile_X0Y0_NN4BEG[2] Tile_X0Y0_NN4BEG[3] Tile_X0Y0_NN4BEG[4]
+ Tile_X0Y0_NN4BEG[5] Tile_X0Y0_NN4BEG[6] Tile_X0Y0_NN4BEG[7] Tile_X0Y0_NN4BEG[8]
+ Tile_X0Y0_NN4BEG[9] Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[1] Tile_X0Y0_S1END[2] Tile_X0Y0_S1END[3]
+ Tile_X0Y0_S2END[0] Tile_X0Y0_S2END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_S2END[3] Tile_X0Y0_S2END[4]
+ Tile_X0Y0_S2END[5] Tile_X0Y0_S2END[6] Tile_X0Y0_S2END[7] Tile_X0Y0_S2MID[0] Tile_X0Y0_S2MID[1]
+ Tile_X0Y0_S2MID[2] Tile_X0Y0_S2MID[3] Tile_X0Y0_S2MID[4] Tile_X0Y0_S2MID[5] Tile_X0Y0_S2MID[6]
+ Tile_X0Y0_S2MID[7] Tile_X0Y0_S4END[0] Tile_X0Y0_S4END[10] Tile_X0Y0_S4END[11] Tile_X0Y0_S4END[12]
+ Tile_X0Y0_S4END[13] Tile_X0Y0_S4END[14] Tile_X0Y0_S4END[15] Tile_X0Y0_S4END[1] Tile_X0Y0_S4END[2]
+ Tile_X0Y0_S4END[3] Tile_X0Y0_S4END[4] Tile_X0Y0_S4END[5] Tile_X0Y0_S4END[6] Tile_X0Y0_S4END[7]
+ Tile_X0Y0_S4END[8] Tile_X0Y0_S4END[9] Tile_X0Y0_SS4END[0] Tile_X0Y0_SS4END[10] Tile_X0Y0_SS4END[11]
+ Tile_X0Y0_SS4END[12] Tile_X0Y0_SS4END[13] Tile_X0Y0_SS4END[14] Tile_X0Y0_SS4END[15]
+ Tile_X0Y0_SS4END[1] Tile_X0Y0_SS4END[2] Tile_X0Y0_SS4END[3] Tile_X0Y0_SS4END[4]
+ Tile_X0Y0_SS4END[5] Tile_X0Y0_SS4END[6] Tile_X0Y0_SS4END[7] Tile_X0Y0_SS4END[8]
+ Tile_X0Y0_SS4END[9] Tile_X0Y0_UserCLKo Tile_X0Y0_W1BEG[0] Tile_X0Y0_W1BEG[1] Tile_X0Y0_W1BEG[2]
+ Tile_X0Y0_W1BEG[3] Tile_X0Y0_W1END[0] Tile_X0Y0_W1END[1] Tile_X0Y0_W1END[2] Tile_X0Y0_W1END[3]
+ Tile_X0Y0_W2BEG[0] Tile_X0Y0_W2BEG[1] Tile_X0Y0_W2BEG[2] Tile_X0Y0_W2BEG[3] Tile_X0Y0_W2BEG[4]
+ Tile_X0Y0_W2BEG[5] Tile_X0Y0_W2BEG[6] Tile_X0Y0_W2BEG[7] Tile_X0Y0_W2BEGb[0] Tile_X0Y0_W2BEGb[1]
+ Tile_X0Y0_W2BEGb[2] Tile_X0Y0_W2BEGb[3] Tile_X0Y0_W2BEGb[4] Tile_X0Y0_W2BEGb[5]
+ Tile_X0Y0_W2BEGb[6] Tile_X0Y0_W2BEGb[7] Tile_X0Y0_W2END[0] Tile_X0Y0_W2END[1] Tile_X0Y0_W2END[2]
+ Tile_X0Y0_W2END[3] Tile_X0Y0_W2END[4] Tile_X0Y0_W2END[5] Tile_X0Y0_W2END[6] Tile_X0Y0_W2END[7]
+ Tile_X0Y0_W2MID[0] Tile_X0Y0_W2MID[1] Tile_X0Y0_W2MID[2] Tile_X0Y0_W2MID[3] Tile_X0Y0_W2MID[4]
+ Tile_X0Y0_W2MID[5] Tile_X0Y0_W2MID[6] Tile_X0Y0_W2MID[7] Tile_X0Y0_W6BEG[0] Tile_X0Y0_W6BEG[10]
+ Tile_X0Y0_W6BEG[11] Tile_X0Y0_W6BEG[1] Tile_X0Y0_W6BEG[2] Tile_X0Y0_W6BEG[3] Tile_X0Y0_W6BEG[4]
+ Tile_X0Y0_W6BEG[5] Tile_X0Y0_W6BEG[6] Tile_X0Y0_W6BEG[7] Tile_X0Y0_W6BEG[8] Tile_X0Y0_W6BEG[9]
+ Tile_X0Y0_W6END[0] Tile_X0Y0_W6END[10] Tile_X0Y0_W6END[11] Tile_X0Y0_W6END[1] Tile_X0Y0_W6END[2]
+ Tile_X0Y0_W6END[3] Tile_X0Y0_W6END[4] Tile_X0Y0_W6END[5] Tile_X0Y0_W6END[6] Tile_X0Y0_W6END[7]
+ Tile_X0Y0_W6END[8] Tile_X0Y0_W6END[9] Tile_X0Y0_WW4BEG[0] Tile_X0Y0_WW4BEG[10] Tile_X0Y0_WW4BEG[11]
+ Tile_X0Y0_WW4BEG[12] Tile_X0Y0_WW4BEG[13] Tile_X0Y0_WW4BEG[14] Tile_X0Y0_WW4BEG[15]
+ Tile_X0Y0_WW4BEG[1] Tile_X0Y0_WW4BEG[2] Tile_X0Y0_WW4BEG[3] Tile_X0Y0_WW4BEG[4]
+ Tile_X0Y0_WW4BEG[5] Tile_X0Y0_WW4BEG[6] Tile_X0Y0_WW4BEG[7] Tile_X0Y0_WW4BEG[8]
+ Tile_X0Y0_WW4BEG[9] Tile_X0Y0_WW4END[0] Tile_X0Y0_WW4END[10] Tile_X0Y0_WW4END[11]
+ Tile_X0Y0_WW4END[12] Tile_X0Y0_WW4END[13] Tile_X0Y0_WW4END[14] Tile_X0Y0_WW4END[15]
+ Tile_X0Y0_WW4END[1] Tile_X0Y0_WW4END[2] Tile_X0Y0_WW4END[3] Tile_X0Y0_WW4END[4]
+ Tile_X0Y0_WW4END[5] Tile_X0Y0_WW4END[6] Tile_X0Y0_WW4END[7] Tile_X0Y0_WW4END[8]
+ Tile_X0Y0_WW4END[9] Tile_X0Y1_E1BEG[0] Tile_X0Y1_E1BEG[1] Tile_X0Y1_E1BEG[2] Tile_X0Y1_E1BEG[3]
+ Tile_X0Y1_E1END[0] Tile_X0Y1_E1END[1] Tile_X0Y1_E1END[2] Tile_X0Y1_E1END[3] Tile_X0Y1_E2BEG[0]
+ Tile_X0Y1_E2BEG[1] Tile_X0Y1_E2BEG[2] Tile_X0Y1_E2BEG[3] Tile_X0Y1_E2BEG[4] Tile_X0Y1_E2BEG[5]
+ Tile_X0Y1_E2BEG[6] Tile_X0Y1_E2BEG[7] Tile_X0Y1_E2BEGb[0] Tile_X0Y1_E2BEGb[1] Tile_X0Y1_E2BEGb[2]
+ Tile_X0Y1_E2BEGb[3] Tile_X0Y1_E2BEGb[4] Tile_X0Y1_E2BEGb[5] Tile_X0Y1_E2BEGb[6]
+ Tile_X0Y1_E2BEGb[7] Tile_X0Y1_E2END[0] Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_E2END[3]
+ Tile_X0Y1_E2END[4] Tile_X0Y1_E2END[5] Tile_X0Y1_E2END[6] Tile_X0Y1_E2END[7] Tile_X0Y1_E2MID[0]
+ Tile_X0Y1_E2MID[1] Tile_X0Y1_E2MID[2] Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[4] Tile_X0Y1_E2MID[5]
+ Tile_X0Y1_E2MID[6] Tile_X0Y1_E2MID[7] Tile_X0Y1_E6BEG[0] Tile_X0Y1_E6BEG[10] Tile_X0Y1_E6BEG[11]
+ Tile_X0Y1_E6BEG[1] Tile_X0Y1_E6BEG[2] Tile_X0Y1_E6BEG[3] Tile_X0Y1_E6BEG[4] Tile_X0Y1_E6BEG[5]
+ Tile_X0Y1_E6BEG[6] Tile_X0Y1_E6BEG[7] Tile_X0Y1_E6BEG[8] Tile_X0Y1_E6BEG[9] Tile_X0Y1_E6END[0]
+ Tile_X0Y1_E6END[10] Tile_X0Y1_E6END[11] Tile_X0Y1_E6END[1] Tile_X0Y1_E6END[2] Tile_X0Y1_E6END[3]
+ Tile_X0Y1_E6END[4] Tile_X0Y1_E6END[5] Tile_X0Y1_E6END[6] Tile_X0Y1_E6END[7] Tile_X0Y1_E6END[8]
+ Tile_X0Y1_E6END[9] Tile_X0Y1_EE4BEG[0] Tile_X0Y1_EE4BEG[10] Tile_X0Y1_EE4BEG[11]
+ Tile_X0Y1_EE4BEG[12] Tile_X0Y1_EE4BEG[13] Tile_X0Y1_EE4BEG[14] Tile_X0Y1_EE4BEG[15]
+ Tile_X0Y1_EE4BEG[1] Tile_X0Y1_EE4BEG[2] Tile_X0Y1_EE4BEG[3] Tile_X0Y1_EE4BEG[4]
+ Tile_X0Y1_EE4BEG[5] Tile_X0Y1_EE4BEG[6] Tile_X0Y1_EE4BEG[7] Tile_X0Y1_EE4BEG[8]
+ Tile_X0Y1_EE4BEG[9] Tile_X0Y1_EE4END[0] Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[11]
+ Tile_X0Y1_EE4END[12] Tile_X0Y1_EE4END[13] Tile_X0Y1_EE4END[14] Tile_X0Y1_EE4END[15]
+ Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[2] Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[4]
+ Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[6] Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[8]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData[11]
+ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData[15]
+ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData[19]
+ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData[22]
+ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData[26]
+ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData[2]
+ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData[4]
+ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData[8]
+ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[0] Tile_X0Y1_FrameData_O[10] Tile_X0Y1_FrameData_O[11]
+ Tile_X0Y1_FrameData_O[12] Tile_X0Y1_FrameData_O[13] Tile_X0Y1_FrameData_O[14] Tile_X0Y1_FrameData_O[15]
+ Tile_X0Y1_FrameData_O[16] Tile_X0Y1_FrameData_O[17] Tile_X0Y1_FrameData_O[18] Tile_X0Y1_FrameData_O[19]
+ Tile_X0Y1_FrameData_O[1] Tile_X0Y1_FrameData_O[20] Tile_X0Y1_FrameData_O[21] Tile_X0Y1_FrameData_O[22]
+ Tile_X0Y1_FrameData_O[23] Tile_X0Y1_FrameData_O[24] Tile_X0Y1_FrameData_O[25] Tile_X0Y1_FrameData_O[26]
+ Tile_X0Y1_FrameData_O[27] Tile_X0Y1_FrameData_O[28] Tile_X0Y1_FrameData_O[29] Tile_X0Y1_FrameData_O[2]
+ Tile_X0Y1_FrameData_O[30] Tile_X0Y1_FrameData_O[31] Tile_X0Y1_FrameData_O[3] Tile_X0Y1_FrameData_O[4]
+ Tile_X0Y1_FrameData_O[5] Tile_X0Y1_FrameData_O[6] Tile_X0Y1_FrameData_O[7] Tile_X0Y1_FrameData_O[8]
+ Tile_X0Y1_FrameData_O[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_FrameStrobe[11]
+ Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_FrameStrobe[13] Tile_X0Y1_FrameStrobe[14] Tile_X0Y1_FrameStrobe[15]
+ Tile_X0Y1_FrameStrobe[16] Tile_X0Y1_FrameStrobe[17] Tile_X0Y1_FrameStrobe[18] Tile_X0Y1_FrameStrobe[19]
+ Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_FrameStrobe[4]
+ Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_FrameStrobe[8]
+ Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_N1END[0] Tile_X0Y1_N1END[1] Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[0] Tile_X0Y1_N2END[1] Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3]
+ Tile_X0Y1_N2END[4] Tile_X0Y1_N2END[5] Tile_X0Y1_N2END[6] Tile_X0Y1_N2END[7] Tile_X0Y1_N2MID[0]
+ Tile_X0Y1_N2MID[1] Tile_X0Y1_N2MID[2] Tile_X0Y1_N2MID[3] Tile_X0Y1_N2MID[4] Tile_X0Y1_N2MID[5]
+ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2MID[7] Tile_X0Y1_N4END[0] Tile_X0Y1_N4END[10] Tile_X0Y1_N4END[11]
+ Tile_X0Y1_N4END[12] Tile_X0Y1_N4END[13] Tile_X0Y1_N4END[14] Tile_X0Y1_N4END[15]
+ Tile_X0Y1_N4END[1] Tile_X0Y1_N4END[2] Tile_X0Y1_N4END[3] Tile_X0Y1_N4END[4] Tile_X0Y1_N4END[5]
+ Tile_X0Y1_N4END[6] Tile_X0Y1_N4END[7] Tile_X0Y1_N4END[8] Tile_X0Y1_N4END[9] Tile_X0Y1_NN4END[0]
+ Tile_X0Y1_NN4END[10] Tile_X0Y1_NN4END[11] Tile_X0Y1_NN4END[12] Tile_X0Y1_NN4END[13]
+ Tile_X0Y1_NN4END[14] Tile_X0Y1_NN4END[15] Tile_X0Y1_NN4END[1] Tile_X0Y1_NN4END[2]
+ Tile_X0Y1_NN4END[3] Tile_X0Y1_NN4END[4] Tile_X0Y1_NN4END[5] Tile_X0Y1_NN4END[6]
+ Tile_X0Y1_NN4END[7] Tile_X0Y1_NN4END[8] Tile_X0Y1_NN4END[9] Tile_X0Y1_S1BEG[0] Tile_X0Y1_S1BEG[1]
+ Tile_X0Y1_S1BEG[2] Tile_X0Y1_S1BEG[3] Tile_X0Y1_S2BEG[0] Tile_X0Y1_S2BEG[1] Tile_X0Y1_S2BEG[2]
+ Tile_X0Y1_S2BEG[3] Tile_X0Y1_S2BEG[4] Tile_X0Y1_S2BEG[5] Tile_X0Y1_S2BEG[6] Tile_X0Y1_S2BEG[7]
+ Tile_X0Y1_S2BEGb[0] Tile_X0Y1_S2BEGb[1] Tile_X0Y1_S2BEGb[2] Tile_X0Y1_S2BEGb[3]
+ Tile_X0Y1_S2BEGb[4] Tile_X0Y1_S2BEGb[5] Tile_X0Y1_S2BEGb[6] Tile_X0Y1_S2BEGb[7]
+ Tile_X0Y1_S4BEG[0] Tile_X0Y1_S4BEG[10] Tile_X0Y1_S4BEG[11] Tile_X0Y1_S4BEG[12] Tile_X0Y1_S4BEG[13]
+ Tile_X0Y1_S4BEG[14] Tile_X0Y1_S4BEG[15] Tile_X0Y1_S4BEG[1] Tile_X0Y1_S4BEG[2] Tile_X0Y1_S4BEG[3]
+ Tile_X0Y1_S4BEG[4] Tile_X0Y1_S4BEG[5] Tile_X0Y1_S4BEG[6] Tile_X0Y1_S4BEG[7] Tile_X0Y1_S4BEG[8]
+ Tile_X0Y1_S4BEG[9] Tile_X0Y1_SS4BEG[0] Tile_X0Y1_SS4BEG[10] Tile_X0Y1_SS4BEG[11]
+ Tile_X0Y1_SS4BEG[12] Tile_X0Y1_SS4BEG[13] Tile_X0Y1_SS4BEG[14] Tile_X0Y1_SS4BEG[15]
+ Tile_X0Y1_SS4BEG[1] Tile_X0Y1_SS4BEG[2] Tile_X0Y1_SS4BEG[3] Tile_X0Y1_SS4BEG[4]
+ Tile_X0Y1_SS4BEG[5] Tile_X0Y1_SS4BEG[6] Tile_X0Y1_SS4BEG[7] Tile_X0Y1_SS4BEG[8]
+ Tile_X0Y1_SS4BEG[9] Tile_X0Y1_UserCLK Tile_X0Y1_W1BEG[0] Tile_X0Y1_W1BEG[1] Tile_X0Y1_W1BEG[2]
+ Tile_X0Y1_W1BEG[3] Tile_X0Y1_W1END[0] Tile_X0Y1_W1END[1] Tile_X0Y1_W1END[2] Tile_X0Y1_W1END[3]
+ Tile_X0Y1_W2BEG[0] Tile_X0Y1_W2BEG[1] Tile_X0Y1_W2BEG[2] Tile_X0Y1_W2BEG[3] Tile_X0Y1_W2BEG[4]
+ Tile_X0Y1_W2BEG[5] Tile_X0Y1_W2BEG[6] Tile_X0Y1_W2BEG[7] Tile_X0Y1_W2BEGb[0] Tile_X0Y1_W2BEGb[1]
+ Tile_X0Y1_W2BEGb[2] Tile_X0Y1_W2BEGb[3] Tile_X0Y1_W2BEGb[4] Tile_X0Y1_W2BEGb[5]
+ Tile_X0Y1_W2BEGb[6] Tile_X0Y1_W2BEGb[7] Tile_X0Y1_W2END[0] Tile_X0Y1_W2END[1] Tile_X0Y1_W2END[2]
+ Tile_X0Y1_W2END[3] Tile_X0Y1_W2END[4] Tile_X0Y1_W2END[5] Tile_X0Y1_W2END[6] Tile_X0Y1_W2END[7]
+ Tile_X0Y1_W2MID[0] Tile_X0Y1_W2MID[1] Tile_X0Y1_W2MID[2] Tile_X0Y1_W2MID[3] Tile_X0Y1_W2MID[4]
+ Tile_X0Y1_W2MID[5] Tile_X0Y1_W2MID[6] Tile_X0Y1_W2MID[7] Tile_X0Y1_W6BEG[0] Tile_X0Y1_W6BEG[10]
+ Tile_X0Y1_W6BEG[11] Tile_X0Y1_W6BEG[1] Tile_X0Y1_W6BEG[2] Tile_X0Y1_W6BEG[3] Tile_X0Y1_W6BEG[4]
+ Tile_X0Y1_W6BEG[5] Tile_X0Y1_W6BEG[6] Tile_X0Y1_W6BEG[7] Tile_X0Y1_W6BEG[8] Tile_X0Y1_W6BEG[9]
+ Tile_X0Y1_W6END[0] Tile_X0Y1_W6END[10] Tile_X0Y1_W6END[11] Tile_X0Y1_W6END[1] Tile_X0Y1_W6END[2]
+ Tile_X0Y1_W6END[3] Tile_X0Y1_W6END[4] Tile_X0Y1_W6END[5] Tile_X0Y1_W6END[6] Tile_X0Y1_W6END[7]
+ Tile_X0Y1_W6END[8] Tile_X0Y1_W6END[9] Tile_X0Y1_WW4BEG[0] Tile_X0Y1_WW4BEG[10] Tile_X0Y1_WW4BEG[11]
+ Tile_X0Y1_WW4BEG[12] Tile_X0Y1_WW4BEG[13] Tile_X0Y1_WW4BEG[14] Tile_X0Y1_WW4BEG[15]
+ Tile_X0Y1_WW4BEG[1] Tile_X0Y1_WW4BEG[2] Tile_X0Y1_WW4BEG[3] Tile_X0Y1_WW4BEG[4]
+ Tile_X0Y1_WW4BEG[5] Tile_X0Y1_WW4BEG[6] Tile_X0Y1_WW4BEG[7] Tile_X0Y1_WW4BEG[8]
+ Tile_X0Y1_WW4BEG[9] Tile_X0Y1_WW4END[0] Tile_X0Y1_WW4END[10] Tile_X0Y1_WW4END[11]
+ Tile_X0Y1_WW4END[12] Tile_X0Y1_WW4END[13] Tile_X0Y1_WW4END[14] Tile_X0Y1_WW4END[15]
+ Tile_X0Y1_WW4END[1] Tile_X0Y1_WW4END[2] Tile_X0Y1_WW4END[3] Tile_X0Y1_WW4END[4]
+ Tile_X0Y1_WW4END[5] Tile_X0Y1_WW4END[6] Tile_X0Y1_WW4END[7] Tile_X0Y1_WW4END[8]
+ Tile_X0Y1_WW4END[9] VDD VSS
Xclkbuf_2_2__f_Tile_X0Y1_UserCLK_regs clknet_0_Tile_X0Y1_UserCLK_regs clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3155_ _1459_ _1460_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3086_ _1390_ _1394_ _1396_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_54_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3988_ _0199_ _2171_ _2172_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5727_ Tile_X0Y1_N4END[9] net128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2939_ _1218_ _1248_ _1249_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_99_Left_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5658_ Tile_X0Y0_FrameData[4] net75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5589_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4609_ _0491_ _0493_ _0497_ _0498_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_112_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_400 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_428 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_398 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_79_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_320 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4960_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4891_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3911_ Tile_X0Y0_S2MID[0] Tile_X0Y0_S4END[7] Tile_X0Y1_W6END[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3842_ _2062_ _2061_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3773_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y0_S1END[2] Tile_X0Y0_E1END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q _2004_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5512_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2724_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q _1040_ _1041_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5443_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2655_ _0142_ _0974_ _0975_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5374_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4325_ Tile_X0Y1_N1END[1] Tile_X0Y1_N2END[3] Tile_X0Y1_N4END[3] Tile_X0Y1_E2END[3]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q
+ _0229_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2586_ _0883_ _0907_ _0908_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4256_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q _0160_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4187_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q _0091_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_2_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3207_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q _1507_ _1508_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3138_ _1443_ _1429_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q
+ _1444_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_85_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3069_ _1089_ _1378_ _1088_ _1379_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_25_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_283 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_285 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_366 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2440_ _0751_ _0772_ _0773_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_142_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2371_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q _0707_ _0708_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5090_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_78_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4110_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1781_ _0014_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4041_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ _2218_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_394 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4943_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_90_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4874_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3825_ _2045_ _2047_ _2048_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3756_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ _1988_ _1989_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_30_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2707_ Tile_X0Y1_E2MID[4] _0147_ _1023_ _1024_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5426_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3687_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1942_ _1943_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput242 net242 Tile_X0Y1_EE4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2638_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q
+ _0959_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput231 net231 Tile_X0Y1_E6BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput220 net220 Tile_X0Y1_E2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput253 net253 Tile_X0Y1_FrameData_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2569_ Tile_X0Y1_N2MID[4] Tile_X0Y1_N4END[4] Tile_X0Y0_E1END[2] Tile_X0Y0_E2END[4]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q
+ _0893_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput286 net286 Tile_X0Y1_S2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput275 net275 Tile_X0Y1_FrameData_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5357_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput264 net264 Tile_X0Y1_FrameData_O[22] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput297 net297 Tile_X0Y1_S2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5288_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4308_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 _0212_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_445 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4239_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q _0143_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_445 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_137_Right_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_128_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_438 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_45_Left_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_334 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3610_ _0033_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q _1875_
+ _1876_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_104_Right_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4590_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3
+ _0479_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3541_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q
+ _1813_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_54_Left_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_115_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3472_ _1755_ _1756_ _1757_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5211_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2423_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q _0754_ _0756_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q _0757_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5142_ _0008_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[8\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2354_ _0691_ _0690_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q
+ _0692_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2285_ Tile_X0Y0_E2MID[7] _0062_ _0065_ _0626_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_437 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4024_ Tile_X0Y1_N1END[0] Tile_X0Y1_E1END[0] Tile_X0Y1_W1END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q
+ _2204_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_84_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5975_ Tile_X0Y1_WW4END[8] net376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4926_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4857_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3808_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q _2033_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q
+ _2034_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4788_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3739_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ _1973_ _1974_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5409_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_79_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_109_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2972_ _0719_ _0720_ _1122_ _1282_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5760_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 net155 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5691_ Tile_X0Y1_FrameStrobe[5] net96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4711_ Tile_X0Y1_N2MID[0] Tile_X0Y0_E2END[0] Tile_X0Y0_S2END[0] Tile_X0Y0_WW4END[3]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q
+ _0593_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_62_Left_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4642_ _0163_ _0526_ _0527_ _0528_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4573_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q _0460_ _0461_
+ _0463_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_3524_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1799_ _1800_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3455_ Tile_X0Y1_N2END[7] Tile_X0Y1_EE4END[2] Tile_X0Y0_S2MID[7] Tile_X0Y1_W2END[7]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q
+ _1741_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_130_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2406_ Tile_X0Y1_N4END[0] Tile_X0Y0_S4END[4] Tile_X0Y1_E6END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q
+ _0741_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3386_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q _1673_ _1675_
+ _1676_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_71_Left_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5125_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2337_ _0105_ _0673_ _0675_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q
+ _0676_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_84_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2268_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q
+ _0610_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_57_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5056_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4007_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q _1608_ _2189_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5958_ Tile_X0Y1_W2MID[7] net353 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_80_Left_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4909_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5889_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 net284 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_444 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_289 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_119_Left_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_128_Left_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_5 Tile_X0Y0_EE4END[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3240_ Tile_X0Y1_N1END[0] Tile_X0Y1_E1END[0] Tile_X0Y1_N2END[0] Tile_X0Y1_E2END[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q
+ _1539_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3171_ _0121_ _1464_ _1474_ _1475_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_137_Left_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_77_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5812_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 net207 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5743_ Tile_X0Y1_NN4END[9] net144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2955_ _1263_ _1264_ _1265_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5674_ Tile_X0Y0_FrameData[20] net61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_60_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2886_ _1163_ _1195_ _1197_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4625_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q _0208_ _0512_
+ _0513_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4556_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q
+ _0448_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3507_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[4\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ _1789_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4487_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q _0378_ _0380_
+ _0383_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q _0384_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_131_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3438_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q _1724_ _1723_
+ _1725_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3369_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6
+ _1658_ _1659_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5108_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_68_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5039_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_122_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_1081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_392 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput31 net31 Tile_X0Y0_E6BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput42 net42 Tile_X0Y0_EE4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput20 net20 Tile_X0Y0_E2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput7 net7 Tile_X0Y0_E2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput64 net64 Tile_X0Y0_FrameData_O[23] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput53 net53 Tile_X0Y0_FrameData_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput75 net75 Tile_X0Y0_FrameData_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_8_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput86 net86 Tile_X0Y0_FrameStrobe_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput97 net97 Tile_X0Y0_FrameStrobe_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2740_ _0598_ _1053_ _1055_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2671_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q Tile_X0Y1_DSP_bot.A1
+ _0987_ _0989_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4410_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q _0309_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q
+ _0310_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5390_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4341_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q _0243_ _0244_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_445 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4272_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q _0176_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3223_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q
+ _1523_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_98_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3154_ Tile_X0Y1_N2MID[7] Tile_X0Y0_EE4END[2] Tile_X0Y0_S2END[7] Tile_X0Y0_W2END[7]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q
+ _1459_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_65_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3085_ _1390_ _1394_ _1395_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3987_ _0955_ _1188_ _1730_ _1651_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q _2171_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5726_ Tile_X0Y1_N4END[8] net121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2938_ _1219_ _1247_ _1248_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5657_ Tile_X0Y0_FrameData[3] net74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2869_ _1178_ _1181_ _1182_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5588_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4608_ _0495_ _0496_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q
+ _0497_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4539_ _0024_ _0430_ _0432_ _0433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_112_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_318 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4890_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3910_ Tile_X0Y1_E6END[0] Tile_X0Y0_S2MID[3] Tile_X0Y0_S4END[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3841_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y0_S1END[2] Tile_X0Y0_W1END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q _2062_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_32_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3772_ _2000_ _2002_ _2003_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5511_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2723_ Tile_X0Y1_NN4END[3] Tile_X0Y1_E1END[1] Tile_X0Y1_E2END[3] Tile_X0Y1_E6END[1]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q
+ _1040_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5442_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2654_ Tile_X0Y1_N1END[2] Tile_X0Y1_N2END[4] Tile_X0Y1_N4END[0] Tile_X0Y1_E2END[4]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q
+ _0974_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5373_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2585_ _0906_ _0132_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q
+ _0907_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4324_ _0045_ _0227_ _0228_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4255_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q _0159_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4186_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q _0090_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3206_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ _1507_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3137_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 Tile_X0Y0_E2MID[2] Tile_X0Y0_S2MID[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q _1443_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_118_Right_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3068_ _1146_ _1377_ _1147_ _1378_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_443 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5709_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 net104 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2370_ _0139_ _0254_ _0707_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4040_ _1026_ _1701_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q
+ _2217_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4942_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4873_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3824_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q _0346_ _2046_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q _2047_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3755_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q _1430_ _1988_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3686_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[1\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ _1943_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2706_ _0027_ _0147_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q
+ _1023_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5425_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput210 net210 Tile_X0Y1_E2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_12_Right_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2637_ _0145_ _0957_ _0958_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput243 net243 Tile_X0Y1_EE4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput221 net221 Tile_X0Y1_E2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput232 net232 Tile_X0Y1_E6BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2568_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q _0891_ _0090_
+ _0892_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput276 net276 Tile_X0Y1_FrameData_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5356_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput254 net254 Tile_X0Y1_FrameData_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput265 net265 Tile_X0Y1_FrameData_O[23] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4307_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 _0211_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput287 net287 Tile_X0Y1_S2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput298 net298 Tile_X0Y1_S2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2499_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q
+ _0828_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5287_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_98_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4238_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q _0142_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4169_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q _0073_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_21_Right_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_30_Right_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_118_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_100_Left_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_46_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3540_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q
+ _1812_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5210_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3471_ _1684_ _1698_ _1756_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2422_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ _0755_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q _0756_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5141_ _0007_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[7\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2353_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q
+ _0691_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_69_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5072_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4023_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q _2200_ _2202_
+ _2203_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2284_ _0061_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q
+ _0625_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_95_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5974_ Tile_X0Y1_WW4END[7] net375 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4925_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4856_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3807_ _2032_ _2033_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4787_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_20_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3738_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q _0916_ _1973_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3669_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q _0188_ _1927_
+ _1928_ _1929_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5408_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5339_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_109_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_90_408 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_370 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2971_ _1148_ _1262_ _1281_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5690_ Tile_X0Y1_FrameStrobe[4] net95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4710_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q _0589_ _0591_
+ _0592_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4641_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[14\]
+ _0527_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4572_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q _0460_ _0461_
+ _0462_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_143_432 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3523_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[9\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ _1800_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3454_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q _1739_ _1738_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q _1740_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2405_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q _0738_ _0740_
+ _0734_ _0736_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3385_ _0063_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q
+ _1674_ _1675_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5124_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_29_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2336_ _0105_ _0374_ _0675_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2267_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q
+ _0609_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5055_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4006_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ _2187_ _2188_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ Tile_X0Y1_W2MID[6] net352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4908_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5888_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 net283 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4839_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_106_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_6 Tile_X0Y0_EE4END[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3170_ _0097_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q
+ _1473_ _1474_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_77_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5811_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 net206 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5742_ Tile_X0Y1_NN4END[8] net137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2954_ _1209_ _1215_ _1264_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5673_ Tile_X0Y0_FrameData[19] net59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2885_ _1163_ _1195_ _1196_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4624_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q _0512_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_6_Right_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4555_ _0446_ _0447_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3506_ _1758_ _1759_ _1788_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4486_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q _0382_ _0383_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3437_ Tile_X0Y0_S2MID[3] Tile_X0Y1_WW4END[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q
+ _1724_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3368_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q _0421_ _1658_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5107_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2319_ _0631_ _0634_ _0655_ _0098_ _0659_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3299_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q _1582_ _1592_
+ _1554_ _1580_ Tile_X0Y1_DSP_bot.C8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_68_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5038_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_0_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_1082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput21 net21 Tile_X0Y0_E6BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput32 net32 Tile_X0Y0_E6BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput43 net43 Tile_X0Y0_EE4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput8 net8 Tile_X0Y0_E2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput10 net10 Tile_X0Y0_E2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput65 net65 Tile_X0Y0_FrameData_O[24] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput54 net54 Tile_X0Y0_FrameData_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput76 net76 Tile_X0Y0_FrameData_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput98 net98 Tile_X0Y0_FrameStrobe_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput87 net87 Tile_X0Y0_FrameStrobe_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Right_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2670_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q _0146_ _0986_
+ _0988_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4340_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q
+ _0243_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4271_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q _0175_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3222_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q
+ _1522_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3153_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q _1457_ _1455_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q _1458_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_68_Right_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3084_ _1392_ _1393_ _1394_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3986_ _0199_ _2169_ _2170_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_77_Right_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5725_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 net120 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2937_ _1220_ _1246_ _1247_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5656_ Tile_X0Y0_FrameData[2] net71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2868_ _0156_ _1180_ _1181_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4607_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q Tile_X0Y1_W1END[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q _0496_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5587_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2799_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 _1113_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4538_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q Tile_X0Y1_W6END[0]
+ _0431_ _0432_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_112_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4469_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q _0366_ _0367_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_86_Right_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_85_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_441 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_95_Right_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_1211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3840_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q _2058_ _2060_
+ _2061_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3771_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q _0875_ _2001_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q _2002_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5510_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2722_ _0151_ _1038_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q
+ _1039_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5441_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2653_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q _0972_ _0143_
+ _0973_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5372_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2584_ _0906_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4323_ Tile_X0Y1_E6END[1] Tile_X0Y0_S2MID[3] Tile_X0Y1_W2END[3] Tile_X0Y1_W6END[1]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q
+ _0227_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_99_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4254_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q _0158_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4185_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q _0089_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3205_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ _1505_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q _1506_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3136_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q _1441_ _1440_
+ _1442_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3067_ _1207_ _1257_ _1374_ _1206_ _1377_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_42_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5708_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 net103 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3969_ Tile_X0Y1_N1END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q
+ _2155_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5639_ Tile_X0Y0_EE4END[5] net40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_385 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_396 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4941_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4872_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3823_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q _0771_ _2046_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_447 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3754_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q _0346_ _1986_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q _1987_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3685_ _1750_ _1751_ _1942_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2705_ _1021_ _1022_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5424_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2636_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q
+ _0957_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput200 net200 Tile_X0Y0_WW4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput222 net222 Tile_X0Y1_E6BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput233 net233 Tile_X0Y1_E6BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput211 net211 Tile_X0Y1_E2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput244 net244 Tile_X0Y1_EE4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2567_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q
+ _0891_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5355_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput255 net255 Tile_X0Y1_FrameData_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput266 net266 Tile_X0Y1_FrameData_O[24] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput277 net277 Tile_X0Y1_FrameData_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2498_ _0826_ _0827_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput299 net299 Tile_X0Y1_S2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput288 net288 Tile_X0Y1_S2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5286_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4306_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 _0210_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_98_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4237_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q _0141_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4168_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q _0072_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4099_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1790_ _0003_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_38_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3119_ _1089_ _1378_ _1426_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_81_821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_439 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_336 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3470_ _1718_ _1754_ _1755_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2421_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q _0213_ _0755_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5140_ _0006_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[6\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2352_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q
+ _0690_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2283_ _0498_ _0503_ _0508_ _0062_ _0624_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5071_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4022_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q _1651_ _2201_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q _2202_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_95_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_439 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5973_ Tile_X0Y1_WW4END[6] net374 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4924_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_35_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4855_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3806_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q
+ _2032_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4786_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_20_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3737_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 _0374_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2
+ _0407_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3668_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[18\]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q _1928_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5407_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2619_ _0775_ _0927_ _0940_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3599_ _0130_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 _1864_ _1865_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5338_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5269_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_87_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_439 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2970_ _1278_ _1279_ _1280_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4640_ _0162_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X
+ _0526_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_441 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4571_ Tile_X0Y1_N4END[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q
+ _0461_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3522_ _1549_ _1550_ _1769_ _1799_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3453_ Tile_X0Y1_N4END[3] Tile_X0Y1_E2END[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q
+ _1739_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2404_ _0135_ _0739_ _0740_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5123_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3384_ Tile_X0Y1_WW4END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q
+ _1674_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2335_ _0673_ _0674_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5054_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4005_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q _0956_ _2187_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5956_ Tile_X0Y1_W2MID[5] net351 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4907_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5887_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 net282 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4838_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4769_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_134_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_7 Tile_X0Y0_EE4END[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5810_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 net205 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5741_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 net127 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2953_ _0882_ _1121_ _1262_ _1263_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5672_ Tile_X0Y0_FrameData[18] net58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_60_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2884_ _0599_ _1194_ _1195_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4623_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q
+ _0511_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4554_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q
+ _0446_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_400 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3505_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1786_ _1787_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4485_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ _0381_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q _0382_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3436_ _0043_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q
+ _1722_ _1723_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3367_ _1362_ _1364_ _1657_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5106_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2318_ _0632_ _0633_ _0654_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ _0658_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5037_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_57_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3298_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6
+ _1591_ _1592_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_1083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5939_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 net334 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput22 net22 Tile_X0Y0_E6BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput33 net33 Tile_X0Y0_EE4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput11 net11 Tile_X0Y0_E2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput9 net9 Tile_X0Y0_E2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput55 net55 Tile_X0Y0_FrameData_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput66 net66 Tile_X0Y0_FrameData_O[25] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput44 net44 Tile_X0Y0_EE4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput99 net99 Tile_X0Y0_FrameStrobe_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput77 net77 Tile_X0Y0_FrameData_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput88 net88 Tile_X0Y0_FrameStrobe_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4270_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q _0174_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3221_ _1518_ _1519_ _1517_ _1520_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q _1521_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3152_ _0057_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q _1456_
+ _1457_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3083_ _1381_ _1383_ _1385_ _1393_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_59_Left_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3985_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q
+ _2169_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5724_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 net119 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2936_ _1221_ _1243_ _1246_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5655_ Tile_X0Y0_FrameData[1] net60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2867_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q _1179_ _1180_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4606_ _0020_ Tile_X0Y1_W1END[2] _0495_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2798_ _1110_ _1112_ _1108_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5586_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_68_Left_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_117_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4537_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q _0023_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q
+ _0431_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_112_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4468_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q
+ _0366_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3419_ _0185_ _1706_ _1705_ _1707_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4399_ Tile_X0Y1_E6END[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q
+ _0299_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_77_Left_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_399 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_86_Left_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_95_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_87_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_141_1212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3770_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q _0525_ _2001_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2721_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q
+ _1038_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_132_Right_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5440_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2652_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q
+ _0972_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_8_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5371_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2583_ _0899_ _0905_ _0886_ _0906_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4322_ _0045_ _0225_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q
+ _0226_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4253_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q _0157_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3204_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q _0207_ _1505_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4184_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q _0088_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3135_ Tile_X0Y0_S2END[3] Tile_X0Y0_WW4END[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q
+ _1441_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3066_ _1207_ _1257_ _1374_ _1376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_50_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3968_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q _0489_ _2153_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q _2154_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5707_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 net102 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2919_ Tile_X0Y1_E2MID[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q
+ _1230_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3899_ Tile_X0Y1_N1END[3] Tile_X0Y1_N4END[1] Tile_X0Y1_N2END[1] Tile_X0Y1_EE4END[1]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q
+ _2104_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5638_ Tile_X0Y0_EE4END[4] net33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5569_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_2_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_445 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4940_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4871_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3822_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ _2044_ _2045_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3753_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q _0880_ _1986_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2704_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q _1021_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3684_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1940_ _1941_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5423_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2635_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q _0954_ _0953_
+ _0956_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput201 net201 Tile_X0Y0_WW4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput234 net234 Tile_X0Y1_EE4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput212 net212 Tile_X0Y1_E2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5354_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput223 net223 Tile_X0Y1_E6BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2566_ _0089_ _0889_ _0890_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput245 net245 Tile_X0Y1_EE4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput267 net267 Tile_X0Y1_FrameData_O[25] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput256 net256 Tile_X0Y1_FrameData_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4305_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 _0209_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5285_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2497_ Tile_X0Y1_N2MID[4] Tile_X0Y1_E2MID[4] Tile_X0Y1_W2MID[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q
+ _0826_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput289 net289 Tile_X0Y1_S2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput278 net278 Tile_X0Y1_FrameData_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_98_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4236_ Tile_X0Y0_SS4END[4] _0140_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4167_ Tile_X0Y0_E2MID[3] _0071_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3118_ _0161_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q _1423_
+ _1424_ _1425_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4098_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1783_ _0002_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_38_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3049_ _1347_ _1348_ _1359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_81_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_426 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_408 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_280 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_14_Left_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_441 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2420_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ _0753_ _0754_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2351_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q _0688_ _0689_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2282_ _0499_ _0502_ _0509_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q
+ _0623_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5070_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4021_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q _0716_ _2201_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_95_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5972_ Tile_X0Y1_WW4END[5] net373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_32_Left_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_35_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4923_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4854_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3805_ Tile_X0Y0_E1END[2] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_W1END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q _2031_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4785_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_20_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3736_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1
+ _0346_ _0321_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Left_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3667_ _0162_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X
+ _1927_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5406_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2618_ _0680_ _0883_ _0939_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3598_ Tile_X0Y0_W2MID[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q
+ _1864_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2549_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 Tile_X0Y0_W2MID[2] Tile_X0Y0_E2MID[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q _0874_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5337_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_87_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5268_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4219_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q _0123_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5199_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_50_Left_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_440 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4570_ Tile_X0Y0_E2END[2] _0031_ _0460_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3521_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1797_ _1798_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3452_ _0044_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q
+ _1737_ _1738_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2403_ Tile_X0Y0_S2MID[2] Tile_X0Y1_W2END[2] Tile_X0Y0_S4END[6] Tile_X0Y1_W6END[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q
+ _0739_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3383_ Tile_X0Y1_N2END[7] Tile_X0Y1_E2END[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q
+ _1673_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5122_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2334_ _0672_ _0104_ _0103_ _0617_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q _0673_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5053_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4004_ _2181_ _2186_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5955_ Tile_X0Y1_W2MID[4] net350 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4906_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5886_ Tile_X0Y1_FrameData[31] net274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4837_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4768_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_134_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3719_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q _1965_ _1966_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4699_ _0255_ Tile_X0Y1_N2MID[2] Tile_X0Y0_E2END[2] Tile_X0Y0_E6END[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q _0582_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_106_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_8 Tile_X0Y0_EE4END[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5740_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 net126 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_106_Left_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2952_ _1213_ _1258_ _1259_ _1262_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5671_ Tile_X0Y0_FrameData[17] net57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2883_ _1192_ _1193_ _1194_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_60_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4622_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 Tile_X0Y0_S2MID[7] Tile_X0Y0_E2MID[7]
+ Tile_X0Y0_W2MID[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q _0510_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4553_ _0445_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3504_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[0\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ _1787_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4484_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q _0213_ _0381_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3435_ Tile_X0Y1_N2END[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q
+ _1722_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_318 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3366_ _0163_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[5\] _1655_ _1656_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5105_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3297_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q _0421_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q
+ _1591_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2317_ _0656_ _0657_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5036_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_0_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5938_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 net324 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_0_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_1084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5869_ Tile_X0Y1_FrameData[14] net255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput23 net23 Tile_X0Y0_E6BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput34 net34 Tile_X0Y0_EE4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput12 net12 Tile_X0Y0_E2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput67 net67 Tile_X0Y0_FrameData_O[26] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput56 net56 Tile_X0Y0_FrameData_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput45 net45 Tile_X0Y0_EE4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput89 net89 Tile_X0Y0_FrameStrobe_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput78 net78 Tile_X0Y0_FrameData_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_113_Right_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3220_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q
+ _1520_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3151_ Tile_X0Y1_N4END[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q
+ _1456_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3082_ _0679_ _0824_ _1391_ _1392_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3984_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q _2167_ _2168_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5723_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 net118 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2935_ _1244_ _1245_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5654_ Tile_X0Y0_FrameData[0] net49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2866_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q
+ _1179_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4605_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q _0492_ _0494_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2797_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q _1111_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q
+ _1112_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5585_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4536_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q Tile_X0Y0_S2MID[2]
+ _0429_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q _0430_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_112_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4467_ _0361_ _0362_ _0363_ _0364_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q
+ _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3418_ Tile_X0Y1_W2MID[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q
+ _1706_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4398_ Tile_X0Y1_N2END[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q _0298_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3349_ _1366_ _1368_ _1640_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5019_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_42_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_1139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_324 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_1213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2720_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q _1036_ _1037_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2651_ _0142_ _0970_ _0971_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_10_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5370_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2582_ _0901_ _0904_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q
+ _0905_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4321_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q
+ _0225_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4252_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q _0156_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3203_ _0170_ _1503_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q
+ _1504_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4183_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q _0087_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3134_ _0057_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q
+ _1439_ _1440_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3065_ _1257_ _1374_ _1375_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3967_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q _0207_ _2153_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5706_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 net101 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2918_ _1228_ _1229_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3898_ _0197_ _2102_ _2103_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5637_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 net23 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2849_ _1151_ _1159_ _1161_ _1162_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5568_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_2_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4519_ Tile_X0Y0_S2MID[7] _0094_ _0095_ _0414_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5499_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_58_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4870_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_32_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3821_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q _1430_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q
+ _2044_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_102_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_287 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3752_ _1985_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2703_ _1007_ _1012_ _1017_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q
+ _1020_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3683_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[18\]
+ _1941_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5422_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2634_ _0952_ _0954_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q
+ _0955_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2565_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q
+ _0889_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput224 net224 Tile_X0Y1_E6BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5353_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput202 net202 Tile_X0Y1_E1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput235 net235 Tile_X0Y1_EE4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput213 net213 Tile_X0Y1_E2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput246 net246 Tile_X0Y1_EE4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput257 net257 Tile_X0Y1_FrameData_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput268 net268 Tile_X0Y1_FrameData_O[26] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4304_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 _0208_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5284_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput279 net279 Tile_X0Y1_FrameData_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2496_ _0824_ _0825_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4235_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q _0139_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_98_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4166_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q _0070_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3117_ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[12\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q _1424_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4097_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1942_ _0001_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_38_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3048_ _1357_ _1358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_81_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4999_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_21_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_1178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2350_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q _0687_ _0688_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2281_ _0621_ _0622_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4020_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ _2199_ _2200_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_95_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ Tile_X0Y1_WW4END[4] net366 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4922_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4853_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_60_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3804_ _2025_ _2028_ _2029_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q _2030_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4784_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3735_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 _0630_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0
+ _0653_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3666_ _1926_ _1925_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5405_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3597_ _1862_ _1863_ _1860_ _1861_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2617_ _0928_ _0932_ _0930_ _0938_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5336_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2548_ _0867_ _0869_ _0871_ _0873_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5267_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4218_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q _0122_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2479_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 _0809_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5198_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_141_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4149_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q _0053_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkload0 clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs clkload0/ZN VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_137_443 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3520_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[7\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ _1798_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3451_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3
+ _1737_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2402_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q _0737_ _0738_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3382_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q _1669_ _1671_
+ _0182_ _1672_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2333_ _0672_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5121_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_127_Right_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5052_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4003_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q _2182_ _2185_
+ _2186_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5954_ Tile_X0Y1_W2MID[3] net349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5885_ Tile_X0Y1_FrameData[30] net273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4905_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4836_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4767_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_119_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3718_ _1964_ _1965_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4698_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q _0575_ _0580_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q _0581_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3649_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ _1912_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_136_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5319_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_102_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_9 Tile_X0Y0_EE4END[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_1159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2951_ _1213_ _1259_ _1261_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5670_ Tile_X0Y0_FrameData[16] net56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2882_ _0131_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[1\] _1193_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_60_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4621_ _0498_ _0503_ _0508_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_402 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4552_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q _0444_ _0441_
+ _0445_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3503_ _1750_ _1785_ _1786_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4483_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q _0210_ _0379_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q _0380_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3434_ Tile_X0Y1_NN4END[2] Tile_X0Y0_S4END[6] Tile_X0Y1_E2END[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q
+ _1721_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3365_ _0163_ _1653_ _1654_ _1655_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3296_ _1585_ _1586_ _1588_ _1590_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2316_ _0632_ _0633_ _0654_ _0656_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5104_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_57_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5035_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_122_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5937_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 net323 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_1085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5868_ Tile_X0Y1_FrameData[13] net254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4819_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5799_ Tile_X0Y0_WW4END[12] net200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput24 net24 Tile_X0Y0_E6BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput13 net13 Tile_X0Y0_E2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput57 net57 Tile_X0Y0_FrameData_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput35 net35 Tile_X0Y0_EE4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput46 net46 Tile_X0Y0_EE4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput68 net68 Tile_X0Y0_FrameData_O[27] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput79 net79 Tile_X0Y0_FrameData_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_19_Right_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_28_Right_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3150_ _0059_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q
+ _1454_ _1455_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3081_ _0598_ _0775_ _1391_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_37_Right_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5722_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 net117 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3983_ Tile_X0Y1_E1END[3] Tile_X0Y1_W1END[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q _2167_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2934_ _0598_ _1221_ _1242_ _1244_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5653_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 net39 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2865_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q _1177_ _1178_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_13_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5584_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_46_Right_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4604_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q _0492_ _0493_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2796_ Tile_X0Y0_S1END[3] Tile_X0Y0_W1END[1] Tile_X0Y0_S2END[7] Tile_X0Y0_W1END[3]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q
+ _1111_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4535_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q _0022_ _0429_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4466_ _0078_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q
+ _0364_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3417_ _0027_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q _0185_
+ _1704_ _1705_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4397_ Tile_X0Y1_N1END[3] _0051_ _0297_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3348_ _0163_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[6\] _1636_ _1638_ _1639_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_97_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3279_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q
+ _1575_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_55_Right_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5018_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_38_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_108_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_447 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_64_Right_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_125_Left_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_5_315 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_73_Right_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_134_Left_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_87_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_336 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_141_1214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_82_Right_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_143_Left_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2650_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q
+ _0970_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_139_1198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2581_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q _0903_ _0904_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4320_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q _0223_ _0224_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4251_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q _0155_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3202_ Tile_X0Y1_N1END[2] Tile_X0Y1_E1END[2] Tile_X0Y1_N2END[6] Tile_X0Y1_E2END[6]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q
+ _1503_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_91_Right_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4182_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q _0086_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3133_ Tile_X0Y1_N2MID[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q
+ _1439_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_2_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3064_ _1255_ _1256_ _1371_ _1372_ _1280_ _1374_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_105_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3966_ _2152_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5705_ Tile_X0Y1_FrameStrobe[19] net91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2917_ Tile_X0Y1_W2MID[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q _1228_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5636_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 net22 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3897_ Tile_X0Y1_E6END[1] Tile_X0Y1_W2END[1] Tile_X0Y0_S2MID[1] Tile_X0Y1_W6END[1]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q
+ _2102_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_128_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2848_ _1129_ _1135_ _1161_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5567_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2779_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q _1091_ _1093_
+ _1094_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5498_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4518_ _0375_ _0377_ _0410_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q
+ _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4449_ _0346_ _0347_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3820_ _2043_ _2042_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_102_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3751_ _1980_ _1983_ _1984_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q
+ _1985_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2702_ _1008_ _1011_ _1018_ _0147_ _1019_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_30_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3682_ _1836_ _1930_ _1932_ _1940_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2633_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 Tile_X0Y1_W2MID[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q
+ _0954_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5421_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput203 net203 Tile_X0Y1_E1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput214 net214 Tile_X0Y1_E2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5352_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput225 net225 Tile_X0Y1_E6BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2564_ _0083_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q _0888_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xoutput236 net236 Tile_X0Y1_EE4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput247 net247 Tile_X0Y1_EE4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput258 net258 Tile_X0Y1_FrameData_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4303_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 _0207_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5283_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2495_ _0822_ _0823_ _0824_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput269 net269 Tile_X0Y1_FrameData_O[27] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_385 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4234_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q _0138_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_98_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4165_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q _0069_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3116_ _0162_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X
+ _1423_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4096_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1786_ _0000_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_38_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3047_ _1351_ _1356_ _1357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_82_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4998_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_21_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3949_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 _1629_ _1708_ _0978_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q _2138_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_136_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5619_ Tile_X0Y0_E2MID[1] net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_1179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_108_Right_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_108_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2280_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q _0620_ _0621_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_96_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_95_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5970_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 net356 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4921_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4852_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3803_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q
+ _2029_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4783_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3734_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 _0482_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3
+ _0468_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3665_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4
+ _0189_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q _1926_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_9_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5404_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2616_ _0935_ _0936_ _0934_ _0937_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3596_ Tile_X0Y0_S1END[1] Tile_X0Y0_S2END[7] Tile_X0Y0_S1END[3] Tile_X0Y0_W1END[3]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q
+ _1863_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5335_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2547_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q _0872_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q
+ _0873_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2478_ _0806_ _0808_ _0804_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5266_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4217_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q _0121_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5197_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4148_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q _0052_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4079_ _0203_ _0827_ _2251_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q
+ _2252_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_43_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_49_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_444 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3450_ _0163_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[0\] _1736_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2401_ Tile_X0Y1_N1END[0] Tile_X0Y1_N2END[2] Tile_X0Y1_E2END[2] Tile_X0Y1_E6END[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q
+ _0737_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3381_ Tile_X0Y1_EE4END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q _1670_ _1671_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5120_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2332_ _0667_ _0670_ _0621_ _0672_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5051_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4002_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q _2184_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q
+ _2185_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_108_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5953_ Tile_X0Y1_W2MID[2] net348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5884_ Tile_X0Y1_FrameData[29] net271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4904_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4835_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_60_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4766_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3717_ Tile_X0Y0_E6END[1] Tile_X0Y0_W2END[1] Tile_X0Y0_SS4END[1] Tile_X0Y0_W6END[1]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q
+ _1964_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4697_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q _0577_ _0579_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q _0580_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3648_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q
+ _1911_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_134_447 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3579_ Tile_X0Y0_E2MID[4] Tile_X0Y0_W2MID[4] Tile_X0Y0_S2MID[4] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q
+ _1848_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_114_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5318_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5249_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_16_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2950_ _1213_ _1259_ _1260_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2881_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q _1165_ _1187_
+ _1190_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q _1192_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4620_ _0508_ _0509_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4551_ _0442_ _0443_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q
+ _0444_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3502_ _1352_ _1749_ _1785_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4482_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ _0379_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3433_ _0163_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[1\] _1720_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5103_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3364_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[5\]
+ _1654_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_29_Left_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_57_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3295_ _0173_ _1589_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q
+ _1590_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2315_ _0654_ _0655_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5034_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_76_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5936_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 net322 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_121_1086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_38_Left_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5867_ Tile_X0Y1_FrameData[12] net253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4818_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5798_ Tile_X0Y0_WW4END[11] net199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4749_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_134_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput25 net25 Tile_X0Y0_E6BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput14 net14 Tile_X0Y0_E2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput58 net58 Tile_X0Y0_FrameData_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput36 net36 Tile_X0Y0_EE4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput47 net47 Tile_X0Y0_EE4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput69 net69 Tile_X0Y0_FrameData_O[28] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_8_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_47_Left_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_88_375 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_283 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_357 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3080_ _1079_ _1080_ _1082_ _1384_ _1390_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_35_445 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3982_ _2166_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_73_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5721_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 net116 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2933_ _0598_ _1242_ _1243_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5652_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 net38 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2864_ _1176_ _1177_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2795_ _0127_ _1109_ _1110_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_13_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5583_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4603_ _0020_ Tile_X0Y0_S2MID[0] _0492_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4534_ _0024_ _0424_ _0427_ _0428_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4465_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3416_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4
+ _1704_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4396_ Tile_X0Y0_S2MID[1] Tile_X0Y0_S4END[5] Tile_X0Y1_W2END[1] Tile_X0Y1_W6END[1]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q
+ _0296_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_5_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3347_ _0163_ _1637_ _1638_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3278_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q
+ _1574_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5017_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_108_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_423 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5919_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 net305 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_1215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_1199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2580_ Tile_X0Y0_S2MID[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q _0902_ _0903_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_4_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4250_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q _0154_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3201_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q _1499_ _1501_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q _1502_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4181_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q _0085_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3132_ _1432_ _1434_ _1436_ _1438_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_2_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3063_ _1371_ _1372_ _1280_ _1373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_326 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3965_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q _2146_ _2151_
+ _2152_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5704_ Tile_X0Y1_FrameStrobe[18] net90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3896_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q _2100_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q
+ _2101_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2916_ _0666_ _0671_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q
+ _0622_ _1227_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5635_ Tile_X0Y0_E6END[11] net32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2847_ _1151_ _1159_ _1160_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5566_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2778_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q _0153_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q
+ _1092_ _1093_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5497_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_2_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4517_ _0411_ _0412_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4448_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 Tile_X0Y0_E2MID[3] Tile_X0Y0_S2MID[3]
+ Tile_X0Y0_W2MID[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q _0346_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4379_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q
+ _0280_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_415 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3750_ _0456_ Tile_X0Y0_W1END[3] Tile_X0Y0_E1END[3] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q
+ _1984_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_102_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2701_ _1007_ _1012_ _1017_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3681_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1938_ _1939_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2632_ _0144_ _0952_ _0953_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5420_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput204 net204 Tile_X0Y1_E1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput226 net226 Tile_X0Y1_E6BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput215 net215 Tile_X0Y1_E2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5351_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2563_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q _0218_ _0417_
+ _0420_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q _0887_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4302_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q _0206_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput237 net237 Tile_X0Y1_EE4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput248 net248 Tile_X0Y1_EE4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5282_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput259 net259 Tile_X0Y1_FrameData_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_364 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4233_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q _0137_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2494_ _0131_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[6\] _0823_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_98_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4164_ Tile_X0Y0_SS4END[1] _0068_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4095_ _0206_ _2262_ _2264_ _2266_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3115_ _1421_ _1422_ _1419_ _0653_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_38_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3046_ _1122_ _1194_ _1338_ _1355_ _1356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_TAPCELL_ROW_81_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4997_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_23_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3948_ _2137_ _2136_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q
+ Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3879_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q _2092_ _2094_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q _2095_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5618_ Tile_X0Y0_E2MID[0] net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5549_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_46_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_364 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4920_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4851_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3802_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q _2027_ _2028_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4782_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3733_ Tile_X0Y0_S2END[1] Tile_X0Y0_S4END[0] Tile_X0Y0_W6END[0] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3664_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q _1922_ _1923_
+ _1924_ _1925_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5403_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2615_ _0910_ _0933_ _0936_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3595_ _0456_ Tile_X0Y0_E1END[3] Tile_X0Y1_N2MID[7] Tile_X0Y0_E2END[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q _1862_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5334_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2546_ Tile_X0Y1_E6END[1] Tile_X0Y0_S2MID[3] Tile_X0Y1_W2END[3] Tile_X0Y1_WW4END[1]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q
+ _0872_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_125_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2477_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q _0807_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q
+ _0808_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_10_Left_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5265_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4216_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q _0120_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5196_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4147_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q _0051_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4078_ _0203_ _1026_ _2251_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3029_ _0989_ _1192_ _1193_ _1339_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_70_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_320 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_141_Right_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_32_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2400_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q _0735_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q
+ _0736_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3380_ _0042_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q _1670_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2331_ _0670_ _0671_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5050_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4001_ _2183_ _2184_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_108_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5952_ Tile_X0Y1_W2MID[1] net347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4903_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5883_ Tile_X0Y1_FrameData[28] net270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4834_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4765_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3716_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q _1957_ _1962_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q _1963_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4696_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ _0578_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q _0579_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_134_437 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3647_ _0190_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 _1909_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q
+ _1910_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3578_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q _1846_ _1847_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2529_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ _0855_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q _0856_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_114_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5317_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_406 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5248_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5179_ Tile_X0Y1_DSP_bot.C9 clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[9\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_389 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_126_1113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2880_ _1191_ Tile_X0Y1_DSP_bot.B1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4550_ Tile_X0Y0_S2MID[3] Tile_X0Y1_W2END[3] Tile_X0Y0_S4END[7] Tile_X0Y1_W6END[1]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q
+ _0443_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3501_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1783_ _1784_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4481_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q
+ _0378_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3432_ _1338_ _1353_ _1719_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3363_ _0162_ Tile_X0Y1_DSP_bot.C5 _1653_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5102_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_111_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3294_ Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[7] Tile_X0Y1_E1END[3] Tile_X0Y1_E2END[7]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q
+ _1589_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2314_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q _0652_ _0647_
+ _0102_ _0654_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_68_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_76_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5935_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 net321 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5866_ Tile_X0Y1_FrameData[11] net252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4817_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_119_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5797_ Tile_X0Y0_WW4END[10] net198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4748_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_107_426 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4679_ _0106_ _0562_ _0563_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput15 net15 Tile_X0Y0_E2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_1_Right_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput26 net26 Tile_X0Y0_E6BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput37 net37 Tile_X0Y0_EE4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput48 net48 Tile_X0Y0_EE4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput59 net59 Tile_X0Y0_FrameData_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_8_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3981_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q _2165_ _2164_
+ _2166_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_73_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5720_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 net115 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2932_ _1238_ _1241_ _1242_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5651_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 net37 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2863_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q
+ _1176_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_87_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2794_ _0456_ Tile_X0Y0_E1END[3] Tile_X0Y1_N2MID[7] Tile_X0Y0_E2END[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q _1109_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_13_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5582_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4602_ _0469_ _0481_ _0487_ _0020_ _0491_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_7_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4533_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q _0426_ _0427_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4464_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ _0079_ _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3415_ _0186_ _0287_ _1702_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q
+ _1703_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4395_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q _0289_ _0294_
+ _0053_ _0295_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_5_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3346_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[6\]
+ _1637_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3277_ _0175_ _1572_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q
+ _1573_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5016_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_108_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5918_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 net304 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5849_ Tile_X0Y1_EE4END[14] net235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Left_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_79_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_1216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3200_ _0083_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q
+ _1500_ _1501_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4180_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q _0084_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3131_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q _1437_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q
+ _1438_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_2_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3062_ _1278_ _1279_ _1372_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3964_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q _2150_ _2148_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q _2151_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5703_ Tile_X0Y1_FrameStrobe[17] net89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3895_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q
+ _2100_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2915_ _0667_ _0670_ _0158_ _0621_ _1226_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5634_ Tile_X0Y0_E6END[10] net31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2846_ _1151_ _1157_ _1158_ _1159_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_128_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5565_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2777_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q Tile_X0Y1_W2END[6]
+ _1092_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5496_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4516_ _0375_ _0377_ _0410_ _0411_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4447_ _0340_ _0341_ _0343_ _0345_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4378_ _0054_ _0278_ _0279_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3329_ _1369_ _1370_ _1621_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_421 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2700_ _1017_ _1018_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_65_Left_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3680_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[13\]
+ _1939_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2631_ Tile_X0Y1_N2MID[3] Tile_X0Y1_E2MID[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q
+ _0952_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_351 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput216 net216 Tile_X0Y1_E2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput205 net205 Tile_X0Y1_E1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5350_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2562_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q _0408_ _0885_
+ _0886_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput227 net227 Tile_X0Y1_E6BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput249 net249 Tile_X0Y1_EE4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4301_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q _0205_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5281_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput238 net238 Tile_X0Y1_EE4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4232_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q _0136_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2493_ _0817_ _0820_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q
+ _0796_ _0822_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_87_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4163_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q _0067_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_74_Left_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_95_441 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4094_ _0205_ _2265_ _0206_ _2266_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3114_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 Tile_X0Y0_S2MID[5] Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_W2MID[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q _1422_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3045_ _1306_ _1325_ _1339_ _1355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_38_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4996_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_23_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_408 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3947_ Tile_X0Y1_N1END[0] Tile_X0Y1_E1END[0] Tile_X0Y1_W1END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q
+ _2137_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_23_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_83_Left_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_136_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3878_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q _1421_ _2093_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q _2094_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5617_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 net12 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2829_ _1138_ _1141_ _1142_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5548_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5479_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_92_Left_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_129_1133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_122_Right_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_445 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4850_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3801_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q _1421_ _2026_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q _2027_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4781_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3732_ Tile_X0Y0_S2END[0] Tile_X0Y0_W6END[1] Tile_X0Y0_S4END[3] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3663_ _0189_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q
+ _1924_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5402_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2614_ _0723_ _0724_ _0935_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3594_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q
+ _1861_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5333_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2545_ _0111_ _0870_ _0871_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2476_ Tile_X0Y0_S1END[1] Tile_X0Y0_W1END[1] Tile_X0Y0_S2END[5] Tile_X0Y0_W1END[3]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q
+ _0807_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5264_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_141_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4215_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q _0119_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5195_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4146_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q _0050_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4077_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q _2246_ _2249_
+ _2250_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3028_ _0988_ _1239_ _1240_ _1338_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_51_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4979_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_137_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2330_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q _0669_ _0670_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4000_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q
+ _2183_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_77_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5951_ Tile_X0Y1_W2MID[0] net346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4902_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5882_ Tile_X0Y1_FrameData[27] net269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4833_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4764_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3715_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q _1959_ _1961_
+ _1962_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4695_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q _0214_ _0578_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3646_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7
+ _1909_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3577_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 Tile_X0Y0_S2MID[5] Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_W2MID[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q _1846_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2528_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q _0208_ _0855_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5316_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5247_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_102_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2459_ Tile_X0Y0_S4END[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q _0789_ _0790_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_28_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5178_ Tile_X0Y1_DSP_bot.C8 clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[8\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_126_1114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4129_ Tile_X0Y1_N2MID[1] _0033_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_54_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3500_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[2\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ _1784_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4480_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q _0376_ _0377_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3431_ _1700_ _1717_ _1718_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_114_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3362_ _1645_ _1648_ _1650_ _1652_ Tile_X0Y1_DSP_bot.C5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2313_ _0652_ _0653_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5101_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3293_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q _1587_ _1588_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_366 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5032_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_111_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_400 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5934_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 net320 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5865_ Tile_X0Y1_FrameData[10] net251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_51_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4816_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5796_ Tile_X0Y0_WW4END[9] net197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4747_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4678_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q
+ _0562_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3629_ _1889_ _1890_ _1891_ _1892_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q
+ _1893_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_103_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput49 net49 Tile_X0Y0_FrameData_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput27 net27 Tile_X0Y0_E6BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput38 net38 Tile_X0Y0_EE4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput16 net16 Tile_X0Y0_E2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_8_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_359 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3980_ Tile_X0Y1_N1END[1] Tile_X0Y1_E1END[1] _0657_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q
+ _2165_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2931_ _1240_ _1241_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_73_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5650_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 net36 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2862_ _1171_ _1174_ _1175_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4601_ _0470_ _0480_ _0486_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q
+ _0490_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2793_ _0127_ _1102_ _1107_ _1108_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_13_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5581_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4532_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q _0425_ _0426_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_392 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4463_ _0078_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 _0361_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3414_ _0186_ _1701_ _1702_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_15_Right_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4394_ _0290_ _0291_ _0292_ _0293_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q
+ _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3345_ _1628_ _1635_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q
+ _1636_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3276_ Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[7] Tile_X0Y1_E1END[3] Tile_X0Y1_E2END[7]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q
+ _1572_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5015_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_38_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_425 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_436 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_447 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_391 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_24_Right_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5917_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 net303 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5848_ Tile_X0Y1_EE4END[13] net249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5779_ Tile_X0Y0_W6END[2] net174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_33_Right_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_88_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Right_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_103_Left_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_51_Right_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_10_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_136_Right_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_112_Left_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_99_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3130_ Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[2] Tile_X0Y0_S2END[6] Tile_X0Y0_W1END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q
+ _1437_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3061_ _1369_ _1370_ _1304_ _1371_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_60_Right_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_121_Left_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_391 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3963_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ _2149_ _2150_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5702_ Tile_X0Y1_FrameStrobe[16] net88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3894_ _0197_ _2098_ _2099_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2914_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q _1224_ _1225_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5633_ Tile_X0Y0_E6END[9] net30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2845_ _1149_ _1150_ _1158_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5564_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_130_Left_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2776_ Tile_X0Y1_N2END[6] Tile_X0Y1_E2END[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q
+ _1091_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4515_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q _0408_ _0409_
+ _0410_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_103_Right_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5495_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_104_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4446_ _0072_ _0344_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q
+ _0345_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4377_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q
+ _0278_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3328_ _1619_ _1620_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3259_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q _1556_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_84_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_443 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2630_ _0725_ _0950_ _0951_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xoutput217 net217 Tile_X0Y1_E2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput206 net206 Tile_X0Y1_E2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2561_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q _0884_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q
+ _0885_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4300_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q _0204_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5280_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput239 net239 Tile_X0Y1_EE4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput228 net228 Tile_X0Y1_E6BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2492_ _0821_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4231_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q _0135_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4162_ Tile_X0Y0_S2END[1] _0066_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3113_ _1420_ _1421_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4093_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q _0204_ _2265_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3044_ _1122_ _1194_ _1338_ _1354_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4995_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_23_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3946_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 _1651_ _1730_ _1164_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q _2136_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3877_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q _1849_ _2093_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5616_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 net11 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2828_ _1139_ _1140_ _1141_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5547_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2759_ _0940_ _1072_ _1074_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_2_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5478_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4429_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q _0328_ _0329_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_129_1134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3800_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q _1849_ _2026_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4780_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3731_ Tile_X0Y0_E6END[0] Tile_X0Y0_S4END[2] Tile_X0Y0_S2END[3] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3662_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6
+ _1923_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3593_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q
+ _1860_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5401_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_62_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2613_ _0910_ _0933_ _0934_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_117_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2544_ Tile_X0Y1_N2END[3] Tile_X0Y1_N4END[3] Tile_X0Y1_E1END[1] Tile_X0Y1_E2END[3]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q
+ _0870_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5332_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_114_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2475_ _0115_ _0805_ _0806_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5263_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5194_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_87_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4214_ Tile_X0Y0_SS4END[0] _0118_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4145_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q _0049_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4076_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q _2248_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q
+ _2249_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3027_ _1324_ _1329_ _1337_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_70_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4978_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3929_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q _2122_ _2123_
+ _2120_ _2121_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_50_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_375 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_406 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_439 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_428 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5950_ Tile_X0Y1_W2END[7] net345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4901_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5881_ Tile_X0Y1_FrameData[26] net268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4832_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_60_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4763_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3714_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ _1960_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q _1961_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4694_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ _0576_ _0577_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3645_ _1907_ _1908_ _1905_ _1906_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3576_ _0128_ _1843_ _0129_ _1845_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2527_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q
+ _0854_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5315_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_114_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5246_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2458_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q _0788_ _0789_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_89_Right_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_102_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5177_ Tile_X0Y1_DSP_bot.C7 clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[7\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2389_ _0723_ _0724_ _0725_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_126_1115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4128_ Tile_X0Y1_E2MID[7] _0032_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4059_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q _1707_ _2234_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_98_Right_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_124_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3430_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[2\] _1716_ _0163_ _1717_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_114_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3361_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q _1651_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q
+ _1652_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5100_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2312_ _0649_ _0651_ _0652_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5031_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3292_ _0412_ Tile_X0Y1_W1END[1] Tile_X0Y0_S2MID[7] Tile_X0Y1_W1END[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q _1587_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_57_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5933_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 net319 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5864_ Tile_X0Y1_FrameData[9] net281 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_51_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_334 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4815_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5795_ Tile_X0Y0_WW4END[8] net196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4746_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4677_ _0554_ _0556_ _0558_ _0560_ _0561_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3628_ Tile_X0Y0_E2END[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q
+ _0193_ _1892_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput28 net28 Tile_X0Y0_E6BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput39 net39 Tile_X0Y0_EE4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_132_1152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput17 net17 Tile_X0Y0_E2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_8_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3559_ _0163_ _1827_ _1828_ _1829_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5229_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_102_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_16_Left_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Right_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_90 net366 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2930_ _0131_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[0\] _1240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_73_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2861_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q _1173_ _1174_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4600_ _0469_ _0481_ _0487_ _0489_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2792_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q _1106_ _1107_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_13_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5580_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4531_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q
+ _0425_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4462_ _0356_ _0359_ _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3413_ Tile_X0Y1_N2END[5] Tile_X0Y1_E2END[5] Tile_X0Y0_SS4END[5] Tile_X0Y1_W2END[5]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q
+ _1701_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4393_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ _0052_ _0293_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3344_ _1628_ _1635_ Tile_X0Y1_DSP_bot.C6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3275_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q _1570_ _1571_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_359 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_26_415 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5916_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 net317 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5847_ Tile_X0Y1_EE4END[12] net248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5778_ Tile_X0Y0_W2MID[7] net173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4729_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_88_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_70_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3060_ _1275_ _1276_ _1302_ _1370_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_67_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5701_ Tile_X0Y1_FrameStrobe[15] net87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3962_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q _0827_ _2149_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3893_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q
+ _2098_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_31_440 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2913_ _1222_ _1223_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q
+ _1224_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5632_ Tile_X0Y0_E6END[8] net29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2844_ _1132_ _1152_ _1154_ _1157_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5563_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2775_ _0951_ _1069_ _1090_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4514_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q _0409_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5494_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4445_ Tile_X0Y1_N2END[4] Tile_X0Y1_E1END[2] Tile_X0Y1_N4END[0] Tile_X0Y1_E2END[4]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q
+ _0344_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4376_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q _0275_ _0277_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3327_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q _1618_ _1598_
+ _1619_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3258_ _0172_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 _1555_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3189_ Tile_X0Y1_N1END[0] Tile_X0Y1_E1END[0] Tile_X0Y1_N2END[0] Tile_X0Y1_E2END[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q
+ _1492_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_104_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_1191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_440 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2560_ Tile_X0Y1_N2MID[6] Tile_X0Y0_E2END[6] Tile_X0Y0_SS4END[3] Tile_X0Y0_W2END[6]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q
+ _0884_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput207 net207 Tile_X0Y1_E2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput218 net218 Tile_X0Y1_E2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput229 net229 Tile_X0Y1_E6BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2491_ _0817_ _0820_ _0796_ _0821_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4230_ Tile_X0Y0_S4END[6] _0134_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_389 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4161_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q _0065_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3112_ _0672_ _0104_ _0039_ _0454_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q _1420_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4092_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 _2258_ _2263_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q _2264_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_67_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3043_ _1122_ _1192_ _1193_ _1353_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4994_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_46_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3945_ _2135_ _2134_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q
+ Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3876_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q _0674_ _2091_
+ _2092_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5615_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 net10 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2827_ _0998_ _1061_ _1136_ _1140_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5546_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2758_ _0679_ _0775_ _1073_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5477_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2689_ _1000_ _1002_ _1006_ _1007_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4428_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q _0325_ _0327_
+ _0328_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_48_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4359_ _0047_ _0260_ _0261_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_129_1135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_425 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_8_Left_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_446 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3730_ Tile_X0Y0_E6END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3661_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6
+ _1921_ _1922_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5400_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2612_ _0928_ _0932_ _0933_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3592_ _0163_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[17\] _1859_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_114_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2543_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q _0868_ _0112_
+ _0869_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5331_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_141_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2474_ _0306_ Tile_X0Y0_E1END[1] Tile_X0Y1_N2MID[5] Tile_X0Y0_E2END[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q _0805_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5262_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_141_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5193_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4213_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q _0117_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4144_ Tile_X0Y1_W2MID[7] _0048_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4075_ _2247_ _2248_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3026_ _1333_ _1334_ _1336_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4977_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3928_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ _2123_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3859_ _2072_ _2075_ _2076_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q
+ _2077_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_109_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5529_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_135_1172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_443 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_437 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4900_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5880_ Tile_X0Y1_FrameData[25] net267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4831_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_31_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4762_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_60_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3713_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q _0214_ _1960_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4693_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q _0210_ _0576_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3644_ Tile_X0Y0_S1END[0] Tile_X0Y0_S2END[0] Tile_X0Y0_W1END[0] Tile_X0Y0_W1END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q
+ _1908_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3575_ _1843_ _1844_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5314_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2526_ _0849_ _0850_ _0853_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5245_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2457_ _0788_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5176_ Tile_X0Y1_DSP_bot.C6 clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[6\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2388_ _0598_ _0721_ _0724_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_126_1116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4127_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q _0031_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4058_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q _1629_ _2232_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q _2233_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3009_ _1315_ _1316_ _1319_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_24_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_89_Left_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_435 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_98_Left_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3360_ Tile_X0Y1_N2MID[3] Tile_X0Y1_E2MID[3] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3
+ Tile_X0Y1_W2MID[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q _1651_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2311_ _0068_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q
+ _0650_ _0651_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5030_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3291_ _0173_ _1583_ _0174_ _1586_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_402 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_68_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5932_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 net333 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_76_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5863_ Tile_X0Y1_FrameData[8] net280 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5794_ Tile_X0Y0_WW4END[7] net195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4814_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_119_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4745_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4676_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q _0559_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q
+ _0560_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3627_ Tile_X0Y0_E1END[0] _0192_ _1891_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput29 net29 Tile_X0Y0_E6BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput18 net18 Tile_X0Y0_E2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3558_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[15\]
+ _1828_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_132_1153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2509_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q _0836_ _0837_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3489_ _1772_ _1773_ _1453_ _1774_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5228_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5159_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X
+ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[5\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_80 Tile_X0Y0_E6END[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_91 net375 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2860_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q _1172_ _1173_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2791_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q _1103_ _1105_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q _1106_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4530_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q
+ _0424_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4461_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q _0358_ _0359_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3412_ _1354_ _1355_ _1700_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4392_ _0051_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 _0292_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3343_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q _1629_ _1634_
+ _1635_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3274_ _0657_ _0412_ Tile_X0Y0_S2MID[7] Tile_X0Y1_W1END[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q _1570_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5013_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_26_438 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Right_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5915_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 net316 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5846_ Tile_X0Y1_EE4END[11] net247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2989_ _1297_ _1298_ _1299_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5777_ Tile_X0Y0_W2MID[6] net172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4728_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4659_ Tile_X0Y0_S2MID[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q _0543_ _0544_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_107_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_351 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3961_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q _1026_ _2147_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q _2148_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5700_ Tile_X0Y1_FrameStrobe[14] net86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2912_ Tile_X0Y1_E2END[3] Tile_X0Y1_WW4END[2] Tile_X0Y0_SS4END[7] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q
+ _1223_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_35_Left_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3892_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 _0254_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3
+ _0231_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5631_ Tile_X0Y0_E6END[7] net28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2843_ _0551_ _0747_ _1132_ _1156_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5562_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2774_ _1070_ _1087_ _1089_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4513_ _0407_ _0408_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5493_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4444_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q _0342_ _0343_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_44_Left_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4375_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q _0275_ _0276_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3326_ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[7\] Tile_X0Y1_DSP_bot.C7 _0162_ _1618_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3257_ _0177_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 _1553_ _1554_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_1_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3188_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q _1488_ _1490_
+ _1491_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_26_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_53_Left_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_441 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5829_ Tile_X0Y1_E6END[4] net226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_1192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput208 net208 Tile_X0Y1_E2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput219 net219 Tile_X0Y1_E2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2490_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q _0819_ _0820_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4160_ Tile_X0Y0_W2MID[7] _0064_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3111_ Tile_X0Y1_N2MID[5] Tile_X0Y0_SS4END[1] Tile_X0Y0_E2END[5] Tile_X0Y0_W2END[5]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q
+ _1419_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4091_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q _0241_ _2263_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3042_ _1121_ _1242_ _1352_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4993_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3944_ Tile_X0Y1_N1END[3] Tile_X0Y1_E1END[3] Tile_X0Y1_W1END[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q
+ _2135_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3875_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q _0816_ _2091_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_101_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5614_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2826_ _1057_ _1132_ _1134_ _1139_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5545_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2757_ _0679_ _0824_ _1072_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5476_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2688_ _1004_ _1005_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q
+ _1006_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4427_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q _0211_ _0326_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q _0327_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4358_ Tile_X0Y0_S1END[0] Tile_X0Y0_S2END[0] Tile_X0Y0_W1END[0] Tile_X0Y0_W1END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ _0260_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4289_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q _0193_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_129_1136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3309_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q _0693_ _1601_
+ _1602_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_61_Left_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_70_Left_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_109_Left_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_43_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3660_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q _0315_ _1921_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2611_ _0930_ _0931_ _0932_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3591_ _1854_ _1855_ _1853_ _1858_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2542_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q
+ _0868_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5330_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_141_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5261_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2473_ _0115_ _0797_ _0803_ _0804_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4212_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q _0116_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_118_Left_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5192_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4143_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q _0047_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4074_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q
+ _2247_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_94_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3025_ _1333_ _1334_ _1335_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_127_Left_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_34_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4976_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3927_ _0198_ _0272_ _2122_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3858_ _0306_ Tile_X0Y0_W1END[1] Tile_X0Y0_S1END[1] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q
+ _2076_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3789_ Tile_X0Y0_E1END[3] Tile_X0Y0_W1END[3] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q _2016_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2809_ _1121_ _1122_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5528_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_3_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_1173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_136_Left_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_105_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5459_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_132_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_2_1__f_Tile_X0Y1_UserCLK_regs clknet_0_Tile_X0Y1_UserCLK_regs clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_128_427 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4830_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_33_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4761_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3712_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ _1958_ _1959_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4692_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q
+ _0575_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3643_ _0255_ Tile_X0Y1_N2MID[0] Tile_X0Y0_E1END[0] Tile_X0Y0_EE4END[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q _1907_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5313_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3574_ Tile_X0Y1_NN4END[5] Tile_X0Y0_S2END[5] Tile_X0Y0_E2END[5] Tile_X0Y0_W2END[5]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q
+ _1843_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2525_ _0849_ _0850_ _0852_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5244_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2456_ _0783_ _0787_ _0788_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5175_ Tile_X0Y1_DSP_bot.C5 clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[5\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4126_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q _0030_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2387_ _0551_ _0679_ _0723_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_126_1117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4057_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q _0839_ _2232_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3008_ _1305_ _1311_ _1310_ _1318_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_355 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4959_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_126_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput380 net380 Tile_X0Y1_WW4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2310_ Tile_X0Y1_N4END[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q
+ _0650_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3290_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q _1584_ _1585_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5931_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 net332 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5862_ Tile_X0Y1_FrameData[7] net279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_51_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5793_ Tile_X0Y0_WW4END[6] net194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4813_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4744_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_119_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4675_ Tile_X0Y0_S2END[4] Tile_X0Y0_W2END[4] Tile_X0Y0_S4END[0] Tile_X0Y0_W6END[0]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q
+ _0559_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3626_ Tile_X0Y1_N2MID[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q _1890_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_131_Right_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput19 net19 Tile_X0Y0_E2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3557_ _0162_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X
+ _1827_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_132_1154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2508_ Tile_X0Y1_N4END[1] Tile_X0Y1_W6END[1] Tile_X0Y1_E6END[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q
+ _0836_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5227_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3488_ _1451_ _1452_ _1773_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2439_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q _0770_ _0769_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q _0772_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5158_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X
+ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[4\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5089_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_56_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1938_ _0013_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_70 Tile_X0Y1_NN4END[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_81 Tile_X0Y0_E6END[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_92 net376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2790_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q _0211_ _1104_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q _1105_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_120_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4460_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q _0357_ _0358_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3411_ _1684_ _1698_ _1699_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4391_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q _0291_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3342_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q _1633_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q
+ _1634_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3273_ _0177_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 _1569_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5012_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_38_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5914_ Tile_X0Y0_S4END[15] net315 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5845_ Tile_X0Y1_EE4END[10] net246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2988_ _1266_ _1272_ _1298_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5776_ Tile_X0Y0_W2MID[5] net171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4727_ _0602_ _0605_ _0607_ _0105_ _0608_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4658_ _0064_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q _0543_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3609_ Tile_X0Y0_EE4END[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q _1875_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4589_ _0472_ _0474_ _0476_ _0478_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_450 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_11_Right_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_431 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_20_Right_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_78_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3960_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q _1742_ _2147_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2911_ Tile_X0Y1_NN4END[3] Tile_X0Y1_E2END[6] Tile_X0Y0_S2MID[6] Tile_X0Y1_W2END[6]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q
+ _1222_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3891_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 _0455_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2
+ _0436_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5630_ Tile_X0Y0_E6END[6] net27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2842_ _0551_ _0747_ _1132_ _1155_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_129_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5561_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2773_ _1070_ _1087_ _1088_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5492_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4512_ Tile_X0Y1_NN4END[7] Tile_X0Y0_WW4END[0] Tile_X0Y0_S4END[3] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q
+ _0407_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_104_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4443_ Tile_X0Y1_E6END[0] Tile_X0Y0_S2MID[4] Tile_X0Y1_W2END[4] Tile_X0Y1_W6END[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q
+ _0342_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4374_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ _0275_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3325_ _1610_ _1617_ Tile_X0Y1_DSP_bot.C7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3256_ _0177_ _0693_ _0171_ _1553_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_1_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3187_ _0140_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q
+ _1489_ _1490_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5828_ Tile_X0Y1_E6END[3] net225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5759_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 net154 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_138_1193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_442 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput209 net209 Tile_X0Y1_E2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3110_ _1416_ _1417_ _1418_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4090_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q _2259_ _2261_
+ _2262_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3041_ _1340_ _1345_ _1351_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4992_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_16_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3943_ _2131_ _2133_ _2134_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_46_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3874_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q _2086_ _2089_
+ _2090_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_101_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5613_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2825_ _1062_ _1136_ _1137_ _1138_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_129_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5544_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2756_ _0942_ _0944_ _1071_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5475_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2687_ Tile_X0Y1_W1END[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q _1005_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4426_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ _0326_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4357_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q _0258_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q
+ _0259_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_412 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4288_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q _0192_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_129_1137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3308_ Tile_X0Y1_W2END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q _1601_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_97_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3239_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q _1535_ _1537_
+ _1538_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_37_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_399 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2610_ _0748_ _0776_ _0825_ _0907_ _0931_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3590_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1856_ _1857_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2541_ _0111_ _0866_ _0867_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2472_ _0799_ _0802_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q
+ _0803_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5260_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_141_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4211_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q _0115_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5191_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4142_ Tile_X0Y1_N2MID[0] _0046_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073_ Tile_X0Y1_E1END[2] Tile_X0Y1_W1END[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q _2246_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_94_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3024_ _1315_ _1316_ _1318_ _1334_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4975_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_34_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_397 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3926_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q _2121_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3857_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q _2074_ _2075_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3788_ _2014_ _2015_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2808_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q _1119_ _1120_
+ _1121_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5527_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2739_ _1050_ _1051_ _1054_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_135_1174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5458_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5389_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4409_ Tile_X0Y0_E1END[1] Tile_X0Y0_E2END[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ _0309_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_445 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4760_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_60_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_112_Right_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3711_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q _0210_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q
+ _1958_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4691_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q _0570_ _0573_
+ _0574_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3642_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q
+ _1906_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5312_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_49_Right_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3573_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q _1839_ _1841_
+ _1842_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2524_ _0850_ _0851_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5243_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2455_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q _0786_ _0787_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5174_ Tile_X0Y1_DSP_bot.C4 clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[4\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2386_ _0679_ _0721_ _0722_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4125_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q _0029_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_1118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4056_ Tile_X0Y1_N1END[1] Tile_X0Y1_W1END[1] _0657_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q
+ _2231_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_58_Right_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3007_ _1315_ _1316_ _1317_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_54_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4958_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4889_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3909_ Tile_X0Y1_E6END[1] Tile_X0Y0_S4END[5] Tile_X0Y0_S2MID[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_67_Right_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput370 net370 Tile_X0Y1_WW4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput381 net381 Tile_X0Y1_WW4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_437 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_76_Right_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_289 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_334 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_85_Right_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_128_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Right_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5930_ Tile_X0Y0_SS4END[15] net331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5861_ Tile_X0Y1_FrameData[6] net278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5792_ Tile_X0Y0_WW4END[5] net193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4812_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4743_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4674_ _0108_ _0557_ _0558_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3625_ _0192_ _0255_ _1889_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3556_ _1817_ _1818_ _1826_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_442 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_1155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2507_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q _0833_ _0835_
+ _0829_ _0831_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5226_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3487_ _1482_ _1551_ _1770_ _1481_ _1772_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2438_ _0770_ _0771_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2369_ _0694_ _0695_ _0705_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q
+ _0139_ _0706_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5157_ Tile_X0Y1_DSP_bot.A3 clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[3\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5088_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_67_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4108_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1806_ _0012_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4039_ _2216_ _2215_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_60 Tile_X0Y1_NN4END[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_71 Tile_X0Y1_NN4END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_82 Tile_X0Y0_EE4END[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_93 Tile_X0Y0_EE4END[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3410_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q _0183_ _1696_
+ _1697_ _1698_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4390_ _0051_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 _0290_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3341_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q _1630_ _1632_
+ _1633_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3272_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q _1561_ _1568_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5011_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_97_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_64_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5913_ Tile_X0Y0_S4END[14] net314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5844_ Tile_X0Y1_EE4END[9] net245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2987_ _1281_ _1294_ _1296_ _1297_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5775_ Tile_X0Y0_W2MID[4] net170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4726_ _0606_ _0607_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4657_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7
+ _0541_ _0542_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3608_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q _1868_ _1873_
+ _1874_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4588_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q _0477_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q
+ _0478_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3539_ _1389_ _1395_ _1396_ _1810_ _1811_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_107_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5209_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_4_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_107_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2910_ _1210_ _1212_ _1214_ _1221_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3890_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1
+ _1651_ _1604_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2841_ _0551_ _0747_ _1154_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5560_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2772_ _1084_ _1085_ _1087_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4511_ _0400_ _0402_ _0404_ _0406_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5491_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4442_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q _0338_ _0073_
+ _0341_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4373_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q _0269_ _0271_
+ _0274_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3324_ _1614_ _1615_ _1616_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q _1617_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3255_ _0163_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[8\] _1552_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_1_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3186_ Tile_X0Y1_WW4END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q
+ _1489_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_140_1210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5827_ Tile_X0Y1_E6END[2] net222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5758_ clknet_1_0__leaf_Tile_X0Y1_UserCLK net153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4709_ Tile_X0Y1_N4END[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q
+ _0590_ _0591_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5689_ Tile_X0Y1_FrameStrobe[3] net94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_138_1194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_Tile_X0Y1_UserCLK_regs Tile_X0Y1_UserCLK_regs clknet_0_Tile_X0Y1_UserCLK_regs
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3040_ _1347_ _1348_ _1350_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4991_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3942_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ _2132_ _2133_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_46_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3873_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q _2088_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q
+ _2089_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_101_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5612_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 net7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2824_ _0998_ _1061_ _1137_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5543_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2755_ _1065_ _1068_ _0951_ _1070_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5474_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2686_ Tile_X0Y1_W1END[3] _0148_ _1004_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4425_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q _0208_ _0324_
+ _0325_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4356_ Tile_X0Y0_E1END[0] Tile_X0Y0_E2END[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q
+ _0258_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3307_ _0022_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q
+ _1599_ _1600_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_140_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4287_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q _0191_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_129_1138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3238_ _0060_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q
+ _1536_ _1537_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3169_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5
+ _1473_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_126_Right_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_80_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2540_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q
+ _0866_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_141_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2471_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q _0801_ _0802_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4210_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q _0114_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5190_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4141_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q _0045_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4072_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q _2239_ _2241_
+ _2243_ _2245_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3023_ _1328_ _1330_ _1331_ _1333_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4974_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3925_ _0198_ _0286_ _2120_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3856_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q _1848_ _2073_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q _2074_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3787_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 _1421_ _1848_ _0884_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q
+ _2015_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2807_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[0\]
+ _1120_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5526_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2738_ _1049_ _1052_ _1053_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_135_1175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5457_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2669_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q _0146_ _0987_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4408_ Tile_X0Y1_N2MID[5] _0076_ _0308_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5388_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4339_ _0234_ _0235_ _0240_ _0242_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_438 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_431 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_392 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_332 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3710_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q
+ _1957_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4690_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q _0572_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q
+ _0573_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3641_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q
+ _1905_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3572_ _0058_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q _1840_
+ _1841_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5311_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2523_ _0776_ _0847_ _0850_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_432 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5242_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2454_ _0784_ _0785_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q
+ _0786_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5173_ Tile_X0Y1_DSP_bot.C3 clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[3\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2385_ _0719_ _0720_ _0721_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4124_ Tile_X0Y0_E6END[0] _0028_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_438 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_126_1119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4055_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q _2230_ _2226_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3006_ _1281_ _1292_ _1293_ _1316_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_83_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4957_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4888_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3908_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2
+ _0455_ _0436_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3839_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q _0875_ _2059_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q _2060_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5509_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput360 net360 Tile_X0Y1_W6BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput371 net371 Tile_X0Y1_WW4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_58_Left_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_67_Left_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_76_Left_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_97_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5860_ Tile_X0Y1_FrameData[5] net277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4811_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5791_ Tile_X0Y0_WW4END[4] net186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4742_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_21_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4673_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y0_E2END[4] Tile_X0Y1_N2MID[4]
+ Tile_X0Y0_E6END[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q _0557_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3624_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q _0454_ _1887_
+ _0191_ _1888_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3555_ _1820_ _1823_ _1824_ _0126_ _1826_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_1156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2506_ _0136_ _0834_ _0835_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3486_ _1551_ _1770_ _1771_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5225_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2437_ Tile_X0Y1_N2MID[0] Tile_X0Y0_S2END[0] Tile_X0Y0_EE4END[1] Tile_X0Y0_W2END[0]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q
+ _0770_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_130_446 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2368_ _0137_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 _0704_ _0705_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5156_ Tile_X0Y1_DSP_bot.A2 clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[2\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5087_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2299_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q _0639_ _0640_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4107_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1803_ _0011_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_143_1230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4038_ Tile_X0Y1_N1END[2] Tile_X0Y1_W1END[2] _0351_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q
+ _2216_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_56_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_50 Tile_X0Y1_N4END[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_61 Tile_X0Y1_NN4END[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_72 Tile_X0Y1_NN4END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_83 Tile_X0Y0_EE4END[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_94 Tile_X0Y0_W2END[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput190 net190 Tile_X0Y0_WW4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_7_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3340_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q _0454_ _1631_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q _1632_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5010_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3271_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q _1562_ _1567_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q _1568_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_38_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5912_ Tile_X0Y0_S4END[13] net313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5843_ Tile_X0Y1_EE4END[8] net244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2986_ _1290_ _1291_ _1293_ _1296_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5774_ Tile_X0Y0_W2MID[3] net169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4725_ Tile_X0Y1_N2MID[4] Tile_X0Y0_S2END[4] Tile_X0Y0_EE4END[0] Tile_X0Y0_W2END[4]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q
+ _0606_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4656_ _0061_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q
+ _0541_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4587_ Tile_X0Y0_E6END[0] Tile_X0Y0_S2END[4] Tile_X0Y0_W2END[4] Tile_X0Y0_W6END[0]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q
+ _0477_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3607_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q _1870_ _1872_
+ _1873_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3538_ _1395_ _1809_ _1810_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3469_ _1752_ _1753_ _1754_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5208_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_4_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5139_ _0005_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[5\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_90_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_366 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_444 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2840_ _0721_ _0747_ _1153_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2771_ _1084_ _1085_ _1086_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4510_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q _0405_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q
+ _0406_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5490_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4441_ _0072_ _0339_ _0340_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_9_Right_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4372_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q _0269_ _0271_
+ _0273_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3323_ Tile_X0Y1_N2MID[1] Tile_X0Y1_E2MID[1] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1
+ Tile_X0Y1_W2MID[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q _1616_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_107_Right_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_13_Left_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3254_ _1549_ _1550_ _1551_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_1_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3185_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q _0488_ _1487_
+ _1488_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_92_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_22_Left_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5826_ Tile_X0Y1_E2MID[7] net221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5757_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 net143 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2969_ _1253_ _1254_ _1279_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4708_ _0028_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q
+ _0590_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5688_ Tile_X0Y1_FrameStrobe[2] net93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_138_1195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4639_ _0459_ _0510_ _0524_ _0523_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_89_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Left_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_91_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Left_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_426 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4990_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3941_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q _0827_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q
+ _2132_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_46_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3872_ _2087_ _2088_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5611_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 net6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2823_ _1129_ _1135_ _1128_ _1136_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_101_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5542_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2754_ _1065_ _1068_ _1069_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5473_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2685_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q _1001_ _1003_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4424_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q _0324_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4355_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q _0255_ _0256_
+ _0257_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3306_ Tile_X0Y1_NN4END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q
+ _1599_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4286_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q _0190_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3237_ Tile_X0Y1_W1END[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q
+ _1536_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3168_ _1466_ _1468_ _1470_ _1472_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3099_ _0124_ _1408_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q
+ _1409_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5809_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 net204 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_399 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2470_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q _0211_ _0800_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q _0801_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_55_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4140_ Tile_X0Y1_W2END[3] _0044_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4071_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q _2244_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q
+ _2245_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3022_ _1312_ _1314_ _1330_ _1332_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_48_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4973_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3924_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q _2119_ _2114_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3855_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q _0607_ _2073_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3786_ _0306_ Tile_X0Y0_S1END[1] Tile_X0Y0_E1END[1] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q
+ _2014_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2806_ _1119_ Tile_X0Y1_DSP_bot.A0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5525_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2737_ _1051_ _1052_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_135_1176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2668_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q Tile_X0Y1_DSP_bot.A1
+ _0986_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5456_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4407_ _0274_ _0276_ _0304_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ _0307_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5387_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2599_ Tile_X0Y1_NN4END[4] Tile_X0Y0_S2END[2] Tile_X0Y0_E2END[2] Tile_X0Y0_W2END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q
+ _0921_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4338_ _0041_ _0239_ _0236_ _0241_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4269_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q _0173_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3640_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q _1888_ _1903_
+ _1904_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3571_ Tile_X0Y0_S4END[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q _1840_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5310_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2522_ _0748_ _0822_ _0823_ _0849_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_114_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5241_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2453_ Tile_X0Y0_S2END[3] Tile_X0Y0_W2END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_W6END[1]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q
+ _0785_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5172_ Tile_X0Y1_DSP_bot.C2 clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[2\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2384_ _0131_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[3\] _0720_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4123_ Tile_X0Y1_N2MID[4] _0027_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4054_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q _2229_ _2228_
+ _2230_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3005_ _1312_ _1314_ _1315_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4956_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4887_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3907_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1
+ _1651_ _1604_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3838_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q _1844_ _2059_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3769_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ _1999_ _2000_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5508_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_133_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5439_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput361 net361 Tile_X0Y1_W6BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput350 net350 Tile_X0Y1_W2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_5_Left_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput372 net372 Tile_X0Y1_WW4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4810_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5790_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 net176 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4741_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_14_391 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4672_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q _0555_ _0109_
+ _0556_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3623_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7
+ _1887_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3554_ _1824_ _1825_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_132_1157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2505_ Tile_X0Y0_S4END[6] Tile_X0Y0_SS4END[6] Tile_X0Y1_W2END[2] Tile_X0Y1_W6END[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q
+ _0834_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3485_ _1549_ _1550_ _1597_ _1768_ _1770_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5224_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2436_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q _0766_ _0768_
+ _0769_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5155_ Tile_X0Y1_DSP_bot.A1 clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2367_ _0046_ _0137_ _0704_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5086_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_110_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2298_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q _0211_ _0638_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q _0639_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_67_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4106_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1801_ _0010_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4037_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q _2214_ _2212_
+ _2215_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_143_1231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_431 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4939_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_40 Tile_X0Y1_FrameStrobe[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_51 Tile_X0Y1_N4END[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_73 Tile_X0Y1_NN4END[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_62 Tile_X0Y1_NN4END[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_84 Tile_X0Y0_EE4END[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_361 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_95 net354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput180 net180 Tile_X0Y0_W6BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput191 net191 Tile_X0Y0_WW4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3270_ _1563_ _1564_ _1566_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q _1567_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_97_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5911_ Tile_X0Y0_S4END[12] net312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_64_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_280 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5842_ Tile_X0Y1_EE4END[7] net243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5773_ Tile_X0Y0_W2MID[2] net168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2985_ _1292_ _1293_ _1295_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4724_ _0105_ _0604_ _0605_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4655_ _0538_ _0539_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q
+ _0540_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4586_ _0029_ _0475_ _0476_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3606_ _0025_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q
+ _1871_ _1872_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3537_ _1072_ _1393_ _1391_ _1809_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3468_ _1354_ _1355_ _1717_ _1753_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_130_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5207_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3399_ _0025_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q
+ _1687_ _1688_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_76_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2419_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q _0210_ _0753_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5138_ _0004_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[4\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_95_Left_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5069_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_107_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2770_ _0937_ _0949_ _0950_ _0725_ _1085_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_129_366 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4440_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q
+ _0339_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4371_ _0269_ _0271_ _0272_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3322_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q _1612_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q
+ _1615_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3253_ _1255_ _1256_ _1373_ _1550_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_3184_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q _0351_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q
+ _1487_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_1_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5825_ Tile_X0Y1_E2MID[6] net220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_92_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5756_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 net142 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2968_ _1273_ _1274_ _1277_ _1278_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5687_ Tile_X0Y1_FrameStrobe[1] net92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4707_ Tile_X0Y0_S4END[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q _0588_ _0589_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_138_1196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4638_ _0524_ _0525_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2899_ _0907_ _1054_ _1210_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4569_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 Tile_X0Y0_E2MID[6] Tile_X0Y0_S2MID[6]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q _0459_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_1_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3940_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q _1026_ _2130_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q _2131_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_46_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3871_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q
+ _2087_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5610_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 net5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2822_ _1130_ _1133_ _1135_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_101_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_140_Right_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5541_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2753_ _1066_ _1067_ _1068_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5472_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2684_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q _1001_ _1002_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4423_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q
+ _0323_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4354_ _0046_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ _0256_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3305_ _0163_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[7\] _1598_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4285_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q _0189_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3236_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q _0488_ _1534_
+ _1535_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3167_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q _1471_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q
+ _1472_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3098_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y0_E1END[2] Tile_X0Y1_N2MID[6]
+ Tile_X0Y0_E2END[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q _1408_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5808_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 net203 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5739_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 net125 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4070_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q
+ _2244_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3021_ _1312_ _1314_ _1331_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4972_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3923_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q _2118_ _2117_
+ _2119_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3854_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q _1420_ _2071_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q _2072_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2805_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q _1096_ _1101_
+ _1118_ _1119_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3785_ _2013_ _2012_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5524_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2736_ _0131_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[2\] _1051_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_135_1177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2667_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q _0979_ _0983_
+ _0985_ Tile_X0Y1_DSP_bot.A1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5455_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4406_ _0273_ _0277_ _0305_ _0306_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2598_ Tile_X0Y0_EE4END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_W2END[7] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q
+ _0920_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5386_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4337_ _0041_ _0239_ _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4268_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q _0172_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3219_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q
+ _1519_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4199_ Tile_X0Y0_E2MID[4] _0103_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3570_ _0080_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q
+ _1838_ _1839_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2521_ _0822_ _0823_ _0847_ _0848_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5240_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_5_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2452_ Tile_X0Y1_NN4END[7] Tile_X0Y0_E1END[1] Tile_X0Y0_E2END[3] Tile_X0Y0_E6END[1]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q
+ _0784_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_18_Right_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5171_ Tile_X0Y1_DSP_bot.C1 clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2383_ _0706_ _0708_ _0714_ _0717_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q
+ _0719_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4122_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q _0026_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4053_ _1651_ _1045_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q
+ _2229_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3004_ _1288_ _1313_ _1314_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_27_Right_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4955_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3906_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q _2108_ _2109_
+ _2106_ _2107_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4886_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3837_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ _2057_ _2058_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3768_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q _0916_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q
+ _1999_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2719_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q
+ _1036_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5507_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3699_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q
+ _1954_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_105_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5438_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput362 net362 Tile_X0Y1_W6BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput351 net351 Tile_X0Y1_W2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput340 net340 Tile_X0Y1_W2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_36_Right_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5369_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput373 net373 Tile_X0Y1_WW4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_45_Right_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_53_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_54_Right_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_115_Left_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_97_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_1110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_63_Right_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_124_Left_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_76_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4740_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_16_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4671_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q
+ _0555_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3622_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1885_ _1886_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_72_Right_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_133_Left_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_127_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3553_ Tile_X0Y1_N2MID[3] Tile_X0Y0_E2END[3] Tile_X0Y0_SS4END[0] Tile_X0Y0_W2END[3]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q
+ _1824_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_132_1158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2504_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q _0832_ _0833_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3484_ _1597_ _1768_ _1769_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5223_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2435_ Tile_X0Y1_N4END[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q
+ _0767_ _0768_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5154_ Tile_X0Y1_DSP_bot.A0 clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[0\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4105_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1799_ _0009_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2366_ _0697_ _0699_ _0701_ _0703_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5085_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2297_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ _0638_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_81_Right_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_96_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_142_Left_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4036_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ _2213_ _2214_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_143_1232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4938_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_41 Tile_X0Y1_FrameStrobe[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_30 Tile_X0Y1_FrameStrobe[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4869_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_74 Tile_X0Y1_NN4END[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_63 Tile_X0Y1_NN4END[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_52 Tile_X0Y1_N4END[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_90_Right_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_85 Tile_X0Y0_SS4END[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_96 net368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_307 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput170 net170 Tile_X0Y0_W2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput181 net181 Tile_X0Y0_W6BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_7_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput192 net192 Tile_X0Y0_WW4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5910_ Tile_X0Y0_S4END[11] net311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_64_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5841_ Tile_X0Y1_EE4END[6] net242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2984_ _1290_ _1291_ _1293_ _1294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5772_ Tile_X0Y0_W2MID[1] net167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4723_ _0058_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q
+ _0603_ _0604_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4654_ Tile_X0Y0_E2END[3] Tile_X0Y0_WW4END[2] Tile_X0Y0_SS4END[3] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q
+ _0539_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4585_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y1_N4END[4] Tile_X0Y1_N2MID[4]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q _0475_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3605_ Tile_X0Y0_W2MID[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q
+ _1871_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3536_ _1399_ _1779_ _1808_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5206_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3467_ _1719_ _1720_ _1734_ _1750_ _1751_ _1752_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_88_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3398_ Tile_X0Y1_W2END[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q
+ _1687_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2418_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q
+ _0752_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_4_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5137_ _0003_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[3\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2349_ Tile_X0Y1_N1END[1] Tile_X0Y1_N2END[5] Tile_X0Y1_E1END[1] Tile_X0Y1_E2END[5]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q
+ _0687_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_84_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5068_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4019_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q _1731_ _2199_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_0_Right_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_446 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_121_Right_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4370_ Tile_X0Y1_N2MID[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q
+ _0049_ _0270_ _0271_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3321_ _0046_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q _1613_
+ _1614_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3252_ _1548_ _1549_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3183_ _0165_ _1484_ _1485_ _1486_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_1_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5824_ Tile_X0Y1_E2MID[5] net219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_92_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5755_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 net141 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2967_ _1275_ _1276_ _1277_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5686_ Tile_X0Y1_FrameStrobe[0] net81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2898_ _1149_ _1208_ _1209_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4706_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q _0587_ _0588_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4637_ Tile_X0Y1_N2MID[7] Tile_X0Y0_S2END[7] Tile_X0Y0_E2END[7] Tile_X0Y0_WW4END[0]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q
+ _0524_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_138_1197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4568_ _0457_ _0458_ _0422_ _0423_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_103_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3519_ _1766_ _1796_ _1797_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4499_ _0395_ _0396_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3870_ Tile_X0Y0_E1END[2] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_W1END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q _2086_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2821_ _1130_ _1133_ _1134_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5540_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2752_ _1063_ _1064_ _1067_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5471_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2683_ Tile_X0Y0_S2MID[5] _0148_ _1001_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4422_ _0317_ _0318_ _0319_ _0320_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q
+ _0322_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4353_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 _0242_ _0254_ _0231_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q _0255_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_140_351 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4284_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[18\] _0188_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3304_ _1595_ _1596_ _1597_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3235_ Tile_X0Y0_S2MID[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q _1534_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3166_ Tile_X0Y0_S1END[2] Tile_X0Y0_S2END[6] Tile_X0Y0_W1END[0] Tile_X0Y0_W1END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q
+ _1471_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_104_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3097_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q _1406_ _1407_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3999_ Tile_X0Y1_E1END[2] Tile_X0Y1_W1END[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q _2182_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5807_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 net202 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5738_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 net124 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5669_ Tile_X0Y0_FrameData[15] net55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_1130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3020_ _1308_ _1323_ _1329_ _1330_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_36_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4971_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3922_ Tile_X0Y1_NN4END[1] Tile_X0Y1_E1END[3] Tile_X0Y1_E2END[1] Tile_X0Y1_E6END[1]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q
+ _2118_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3853_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ _2071_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2804_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q _1117_ _1118_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3784_ _0255_ Tile_X0Y0_S1END[0] Tile_X0Y0_E1END[0] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q
+ _2013_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5523_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2735_ _1027_ _1035_ _1047_ _0131_ _1050_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2666_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q _0978_ _0984_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q _0985_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5454_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_132_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5385_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4405_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q _0288_ _0303_
+ _0305_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_132_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2597_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q _0916_ _0918_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q _0919_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4336_ _0237_ _0238_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q
+ _0239_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4267_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q _0171_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3218_ Tile_X0Y1_N1END[0] Tile_X0Y1_E1END[0] Tile_X0Y1_N2END[0] Tile_X0Y1_E2END[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q
+ _1518_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4198_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q _0102_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3149_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3
+ _1454_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_19_Left_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_131_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Left_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_104_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_37_Left_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_92_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_46_Left_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2520_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[2\]
+ _0844_ _0847_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2451_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q _0777_ _0782_
+ _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5170_ Tile_X0Y1_DSP_bot.C0 clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[0\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2382_ _0709_ _0718_ Tile_X0Y1_DSP_bot.B3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4121_ Tile_X0Y0_S2MID[1] _0025_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4052_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q _1731_ _2227_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q _2228_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3003_ _1285_ _1286_ _1287_ _1313_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_83_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4954_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3905_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ _2109_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4885_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_32_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3836_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q _0916_ _2057_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3767_ _1998_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5506_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2718_ _0152_ _1033_ _1035_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3698_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q _1952_ _1953_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2649_ Tile_X0Y1_EE4END[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q
+ _0968_ _0969_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput330 net330 Tile_X0Y1_SS4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput341 net341 Tile_X0Y1_W2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput352 net352 Tile_X0Y1_W2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5437_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_120_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5368_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput363 net363 Tile_X0Y1_W6BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput374 net374 Tile_X0Y1_WW4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4319_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q
+ _0223_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5299_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_15_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_1111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_400 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4670_ _0108_ _0553_ _0554_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3621_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[17\]
+ _1886_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3552_ _1822_ _1823_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2503_ Tile_X0Y1_NN4END[2] Tile_X0Y1_EE4END[2] Tile_X0Y1_E1END[0] Tile_X0Y1_E6END[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q
+ _0832_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3483_ _1622_ _1766_ _1767_ _1768_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5222_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2434_ _0118_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q
+ _0767_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_135_Right_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2365_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q _0702_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q
+ _0703_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5153_ _0019_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[19\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4104_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1946_ _0008_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_363 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5084_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2296_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ _0636_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q _0637_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_67_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4035_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q _0956_ _2213_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_143_1233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5986_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 net372 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_50_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4937_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_31 Tile_X0Y1_FrameStrobe[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4868_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_20 Tile_X0Y1_E6END[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_64 Tile_X0Y1_NN4END[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_53 Tile_X0Y1_N4END[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_42 Tile_X0Y1_FrameStrobe[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_363 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_75 Tile_X0Y1_W2MID[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_3819_ _0456_ Tile_X0Y0_W1END[3] Tile_X0Y0_E1END[3] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q
+ _2043_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4799_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_97 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_86 Tile_X0Y0_SS4END[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput160 net160 Tile_X0Y0_W2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput182 net182 Tile_X0Y0_W6BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_7_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput171 net171 Tile_X0Y0_W2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput193 net193 Tile_X0Y0_WW4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_102_Right_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_87_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_120_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_427 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5840_ Tile_X0Y1_EE4END[5] net241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2983_ _0907_ _1194_ _1293_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5771_ Tile_X0Y0_W2MID[0] net166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4722_ Tile_X0Y1_N4END[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q
+ _0603_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4653_ Tile_X0Y1_NN4END[7] Tile_X0Y0_S2END[6] Tile_X0Y0_E2END[6] Tile_X0Y0_W2END[6]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q
+ _0538_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4584_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q _0473_ _0030_
+ _0474_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3604_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q _0428_ _0435_
+ _1869_ _1870_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3535_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1806_ _1807_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3466_ _1338_ _1353_ _1735_ _1751_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5205_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2417_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q _0749_ _0750_
+ _0751_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3397_ Tile_X0Y1_NN4END[2] Tile_X0Y1_E2END[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q
+ _1686_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_4_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5136_ _0002_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[2\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2348_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q _0681_ _0682_
+ _0685_ _0686_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2279_ _0618_ _0619_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q
+ _0620_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5067_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_96_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4018_ _2198_ _2197_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5969_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 net355 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_111_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3320_ Tile_X0Y1_E2MID[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q _1613_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3251_ _0163_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[9\] _1547_ _1548_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3182_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q _1483_ _1485_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_100_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5823_ Tile_X0Y1_E2MID[4] net218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_92_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5754_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 net140 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2966_ _1273_ _1274_ _1276_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5685_ Tile_X0Y0_FrameData[31] net73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2897_ _0882_ _0988_ _1121_ _0824_ _1208_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4705_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 _0587_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4636_ Tile_X0Y1_N4END[7] Tile_X0Y0_S4END[3] Tile_X0Y0_EE4END[0] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q
+ _0523_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4567_ Tile_X0Y0_S1END[3] Tile_X0Y0_W1END[1] Tile_X0Y0_S2END[7] Tile_X0Y0_W1END[3]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q
+ _0458_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3518_ _1641_ _1764_ _1765_ _1796_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4498_ Tile_X0Y0_E6END[1] Tile_X0Y0_S2END[3] Tile_X0Y0_W2END[3] Tile_X0Y0_W6END[1]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q
+ _0395_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3449_ _1720_ _1734_ _1735_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5119_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_72_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_429 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2820_ _1059_ _1131_ _1133_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2751_ _1056_ _1058_ _1060_ _1066_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5470_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2682_ _0631_ _0634_ _0655_ _0148_ _1000_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4421_ _0317_ _0318_ _0319_ _0320_ _0321_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4352_ Tile_X0Y1_N2MID[1] Tile_X0Y1_E2MID[1] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1
+ Tile_X0Y1_W2MID[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q _0254_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4283_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q _0187_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3303_ _1371_ _1372_ _1596_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3234_ _0168_ _1531_ _1532_ _1533_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_322 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3165_ _0119_ _1469_ _1470_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3096_ Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[2] Tile_X0Y0_S2END[6] Tile_X0Y0_W1END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q
+ _1406_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3998_ _2176_ _2179_ _2180_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q _2181_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_22_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5806_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 net192 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5737_ Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A net123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2949_ _0552_ _0989_ _1259_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5668_ Tile_X0Y0_FrameData[14] net54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5599_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4619_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q _0504_ _0507_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q _0508_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_336 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_1131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4970_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3921_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q _2116_ _2117_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3852_ _2070_ _2069_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_42_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2803_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q _1116_ _1115_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q _1117_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3783_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 _0346_ _1429_ _0538_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q
+ _2012_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5522_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2734_ _1028_ _1034_ _1048_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q
+ _1049_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2665_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q _0967_ _0969_
+ _0984_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5453_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_132_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2596_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q _0917_ _0918_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5384_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4404_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q _0288_ _0303_
+ _0304_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4335_ Tile_X0Y0_S2MID[4] Tile_X0Y0_S4END[4] Tile_X0Y1_W2END[4] Tile_X0Y1_W6END[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q
+ _0238_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_113_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4266_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q _0170_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4197_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q _0101_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3217_ _0489_ _0351_ Tile_X0Y0_S2MID[0] Tile_X0Y1_W1END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q _1517_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_67_450 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_420 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3148_ _1451_ _1452_ _1453_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_42_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3079_ _1379_ _1387_ _1388_ _1389_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_110 net381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_391 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_116_Right_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2450_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q _0779_ _0781_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q _0782_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2381_ _0714_ _0717_ _0718_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4120_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q _0024_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4051_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ _2227_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3002_ _1305_ _1308_ _1309_ _1312_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_83_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4953_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3904_ _0196_ _0272_ _2108_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4884_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_62_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3835_ _2056_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3766_ _1993_ _1996_ _1997_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q
+ _1998_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5505_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2717_ _0152_ _1033_ _1034_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3697_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q
+ _1952_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5436_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_126_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2648_ _0134_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q
+ _0968_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput353 net353 Tile_X0Y1_W2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput320 net320 Tile_X0Y1_SS4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput331 net331 Tile_X0Y1_SS4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput342 net342 Tile_X0Y1_W2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput364 net364 Tile_X0Y1_W6BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5367_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput375 net375 Tile_X0Y1_WW4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2579_ _0064_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q _0902_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5298_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4318_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q _0221_ _0220_
+ _0222_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4249_ Tile_X0Y0_SS4END[7] _0153_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_53_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_1112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_361 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_1_Left_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3620_ _1836_ _1858_ _1883_ _1885_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_3551_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q _1821_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q
+ _1822_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2502_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q _0830_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q
+ _0831_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3482_ _1371_ _1372_ _1595_ _1767_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_142_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5221_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2433_ Tile_X0Y0_W6END[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q _0765_ _0766_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2364_ Tile_X0Y0_S2END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_W2END[1] Tile_X0Y0_W6END[1]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q
+ _0702_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5152_ _0018_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[18\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4103_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1797_ _0007_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5083_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2295_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q _0208_ _0636_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4034_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q _1188_ _2211_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q _2212_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_67_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_1234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5985_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 net371 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_50_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4936_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_32 Tile_X0Y1_FrameStrobe[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4867_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_10 Tile_X0Y0_EE4END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_21 Tile_X0Y1_E6END[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_54 Tile_X0Y1_N4END[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_43 Tile_X0Y1_N4END[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_65 Tile_X0Y1_NN4END[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_353 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3818_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 _0674_ _0815_ _1410_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q
+ _2042_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4798_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_98 net181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_87 Tile_X0Y0_SS4END[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_76 net357 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_3749_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q _1982_ _1983_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput150 net150 Tile_X0Y0_NN4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5419_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_79_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput161 net161 Tile_X0Y0_W2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput183 net183 Tile_X0Y0_W6BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput172 net172 Tile_X0Y0_W2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput194 net194 Tile_X0Y0_WW4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2982_ _1290_ _1291_ _1292_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5770_ Tile_X0Y0_W2END[7] net165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4721_ Tile_X0Y0_W6END[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q _0601_ _0602_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4652_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q _0535_ _0537_
+ _0531_ _0533_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3603_ Tile_X0Y0_E2MID[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q _1869_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4583_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q
+ _0473_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3534_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[12\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ _1807_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3465_ _1121_ _1242_ _1736_ _1748_ _1750_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5204_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2416_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q _0483_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q
+ _0750_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3396_ Tile_X0Y1_EE4END[3] Tile_X0Y1_WW4END[1] Tile_X0Y0_S4END[4] _0242_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q _1685_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5135_ _0001_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2347_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q _0684_ _0685_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2278_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q
+ _0619_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5066_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4017_ Tile_X0Y1_N1END[3] Tile_X0Y1_E1END[3] Tile_X0Y1_W1END[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q
+ _2198_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_25_434 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_64_Left_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5968_ Tile_X0Y1_W6END[11] net365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4919_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_40_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5899_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 net294 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_73_Left_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_334 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_82_Left_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_113_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_423 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_91_Left_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3250_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q _1545_ _1546_
+ _0163_ _1547_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3181_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q
+ _1484_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_120_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_140_1204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5822_ Tile_X0Y1_E2MID[3] net217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5753_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A net139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4704_ _0581_ _0586_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2965_ _1267_ _1271_ _1270_ _1275_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5684_ Tile_X0Y0_FrameData[30] net72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2896_ _1204_ _1205_ _1207_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4635_ _0518_ _0522_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4566_ _0456_ Tile_X0Y0_E1END[3] Tile_X0Y1_N2MID[7] Tile_X0Y0_E2END[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q _0457_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3517_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1794_ _1795_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_361 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4497_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q _0386_ _0388_
+ _0392_ _0394_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XPHY_EDGE_ROW_139_Left_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3448_ _0162_ Tile_X0Y1_DSP_bot.C1 _1733_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q
+ _1734_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3379_ Tile_X0Y0_S4END[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q
+ _1668_ _1669_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5118_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_84_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5049_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_138_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2750_ _0997_ _1062_ _1064_ _1065_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2681_ _0632_ _0633_ _0654_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ _0999_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4420_ Tile_X0Y0_E6END[0] _0075_ _0077_ _0320_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4351_ _0253_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4282_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q _0186_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3302_ _1552_ _1594_ _1595_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3233_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q _1530_ _1532_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_58_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3164_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y0_E1END[2] Tile_X0Y1_N2MID[6]
+ Tile_X0Y0_E2END[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q _1469_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3095_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q _1404_ _0125_
+ _1405_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3997_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q
+ _2180_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5805_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 net191 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5736_ Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A net122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_289 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2948_ _0747_ _1050_ _1051_ _1258_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5667_ Tile_X0Y0_FrameData[13] net53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_20_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2879_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q _1165_ _1187_
+ _1190_ _1191_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4618_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q _0506_ _0507_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5598_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4549_ Tile_X0Y1_N1END[1] Tile_X0Y1_N2END[3] Tile_X0Y1_E2END[3] Tile_X0Y1_E6END[1]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q
+ _0442_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_89_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_353 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_128_1132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3920_ _2115_ _2116_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_34_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3851_ _0255_ Tile_X0Y0_W1END[0] Tile_X0Y0_S1END[0] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q
+ _2070_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3782_ _2011_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_42_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2802_ Tile_X0Y1_W2MID[6] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q
+ _1116_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5521_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2733_ _1027_ _1035_ _1047_ Tile_X0Y1_DSP_bot.B2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2664_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q _0980_ _0982_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q _0983_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5452_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2595_ Tile_X0Y0_E2MID[2] Tile_X0Y0_W2MID[2] Tile_X0Y0_S2MID[2] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q
+ _0917_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5383_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4403_ _0295_ _0302_ _0050_ _0303_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4334_ Tile_X0Y1_N1END[2] Tile_X0Y1_N2END[4] Tile_X0Y1_E2END[4] Tile_X0Y1_E6END[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q
+ _0237_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_59_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4265_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q _0169_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3216_ _1502_ _1504_ _1516_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4196_ Tile_X0Y0_EE4END[1] _0100_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3147_ _1090_ _1145_ _1377_ _1452_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3078_ _1086_ _1386_ _1388_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5719_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 net114 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_447 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_100 net193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_1095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2380_ _0139_ _0716_ _0141_ _0717_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4050_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q _2225_ _2224_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q _2226_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3001_ _1308_ _1309_ _1311_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4952_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4883_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3903_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q _2107_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_392 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3834_ _2051_ _2054_ _2055_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q
+ _2056_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_62_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3765_ _0306_ Tile_X0Y0_W1END[1] Tile_X0Y0_E1END[1] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q
+ _1997_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3696_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q _1948_ _1950_
+ _1951_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5504_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2716_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q _1032_ _1030_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q _1033_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2647_ Tile_X0Y1_W2END[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q _0966_ _0967_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xoutput310 net310 Tile_X0Y1_S4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5435_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput332 net332 Tile_X0Y1_SS4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput321 net321 Tile_X0Y1_SS4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput343 net343 Tile_X0Y1_W2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput365 net365 Tile_X0Y1_W6BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput354 net354 Tile_X0Y1_W6BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5366_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput376 net376 Tile_X0Y1_WW4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2578_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7
+ _0900_ _0901_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5297_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4317_ _0208_ _0210_ _0211_ _0213_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q _0221_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_101_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4248_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q _0152_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4179_ Tile_X0Y0_S2MID[6] _0083_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Right_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_136_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_23_Right_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_32_Right_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3550_ Tile_X0Y1_N4END[6] Tile_X0Y0_SS4END[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q
+ _1821_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2501_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q
+ _0830_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5220_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3481_ _1641_ _1764_ _1765_ _1766_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_41_Right_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2432_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q _0764_ _0765_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2363_ _0092_ _0700_ _0701_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5151_ _0017_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[17\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_102_Left_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5082_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_110_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4102_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1794_ _0006_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2294_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q
+ _0635_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4033_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q _1627_ _2211_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_143_1235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_1224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Right_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5984_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 net370 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_111_Left_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_50_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4935_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4866_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_11 Tile_X0Y0_EE4END[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_22 Tile_X0Y1_E6END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_33 Tile_X0Y1_FrameStrobe[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_66 Tile_X0Y1_NN4END[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_55 Tile_X0Y1_N4END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_44 Tile_X0Y1_N4END[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4797_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3817_ _2041_ _2040_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3748_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q _0815_ _1981_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q _1982_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_99 net182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_77 net364 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_88 Tile_X0Y0_W2END[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_3679_ _1416_ _1417_ _1777_ _1938_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_1
Xoutput151 net151 Tile_X0Y0_NN4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput140 net140 Tile_X0Y0_NN4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_120_Left_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5418_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_133_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput184 net184 Tile_X0Y0_W6BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5349_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput162 net162 Tile_X0Y0_W2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput195 net195 Tile_X0Y0_WW4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput173 net173 Tile_X0Y0_W2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_332 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_432 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_131_1150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_324 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2981_ _1284_ _1288_ _1289_ _1291_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4720_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q _0253_ _0601_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4651_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q _0536_ _0537_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3602_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q _1865_ _1866_
+ _1867_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q _1868_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4582_ _0029_ _0471_ _0472_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3533_ _1776_ _1805_ _1806_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3464_ _1736_ _1748_ _1749_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5203_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_88_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2415_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 Tile_X0Y0_W2MID[0] Tile_X0Y0_S2MID[0]
+ _0316_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q
+ _0749_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5134_ _0000_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[0\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3395_ _1340_ _1345_ _1356_ _1684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2346_ Tile_X0Y0_S2MID[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q _0683_ _0684_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2277_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q
+ _0618_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5065_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4016_ _2194_ _2196_ _2197_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5967_ Tile_X0Y1_W6END[10] net364 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4918_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_52_287 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5898_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 net293 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4849_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_4_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_394 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3180_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q
+ _1483_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_19_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_1205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5821_ Tile_X0Y1_E2MID[2] net216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5752_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A net138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2964_ _1219_ _1247_ _1274_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4703_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q _0582_ _0585_
+ _0586_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5683_ Tile_X0Y0_FrameData[29] net70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2895_ _1204_ _1205_ _1206_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4634_ _0110_ _0519_ _0521_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q
+ _0522_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4565_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2
+ _0455_ _0436_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q
+ _0456_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3516_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[6\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ _1795_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Right_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4496_ _0387_ _0389_ _0391_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q _0393_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3447_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[1\]
+ _1733_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3378_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q _0672_ _1668_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5117_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2329_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q _0668_ _0669_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5048_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_83_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_287 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2680_ _0995_ _0996_ _0998_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4350_ _0247_ _0252_ _0253_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3301_ _0162_ Tile_X0Y1_DSP_bot.C8 _1593_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q
+ _1594_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4281_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q _0185_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3232_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q
+ _1531_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_97_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3163_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q _1467_ _0120_
+ _1468_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3094_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q
+ _1404_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_37_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5804_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 net190 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3996_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q _2178_ _2179_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_45_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5735_ Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A net136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2947_ _1255_ _1256_ _1257_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5666_ Tile_X0Y0_FrameData[12] net52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_20_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2878_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q _1189_ _1190_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4617_ _0505_ _0506_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5597_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_116_351 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4548_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q _0438_ _0440_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q _0441_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4479_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_79_Right_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_88_Right_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_117_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_97_Right_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_59_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3850_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q _2066_ _2068_
+ _2069_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3781_ _2006_ _2009_ _2010_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q
+ _2011_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_42_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2801_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q _1113_ _1114_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q _1115_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5520_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2732_ _1047_ _1048_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2663_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q _0788_ _0981_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q _0982_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5451_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2594_ _0912_ _0914_ _0916_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5382_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4402_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q _0296_ _0301_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q _0302_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4333_ _0234_ _0235_ _0236_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4264_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q _0168_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3215_ _1514_ _1515_ _1516_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4195_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q _0099_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3146_ _1428_ _1450_ _1451_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3077_ _1380_ _1386_ _1387_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5718_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 net113 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3979_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q _2163_ _2161_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q _2164_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5649_ Tile_X0Y0_EE4END[15] net35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_130_Right_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_48_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_101 net198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_1170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3000_ _1308_ _1309_ _1310_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4951_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4882_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3902_ _0196_ _0286_ _2106_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3833_ _0306_ Tile_X0Y0_W1END[1] Tile_X0Y0_E1END[1] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q
+ _2055_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_32_363 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3764_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q _1995_ _1996_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3695_ _0067_ _1949_ _1950_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5503_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2715_ Tile_X0Y1_E2MID[5] _0149_ _1031_ _1032_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2646_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q _0965_ _0966_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput300 net300 Tile_X0Y1_S2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5434_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput344 net344 Tile_X0Y1_W2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput311 net311 Tile_X0Y1_S4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput333 net333 Tile_X0Y1_SS4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput322 net322 Tile_X0Y1_SS4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput377 net377 Tile_X0Y1_WW4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput366 net366 Tile_X0Y1_WW4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput355 net355 Tile_X0Y1_W6BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5365_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2577_ _0061_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q
+ _0900_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5296_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4316_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q _0219_ _0220_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4247_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q _0151_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4178_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q _0082_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3129_ _0122_ _1435_ _1436_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2500_ _0136_ _0828_ _0829_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3480_ _1369_ _1370_ _1620_ _1765_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_115_449 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2431_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 _0764_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5150_ _0016_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[16\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2362_ Tile_X0Y1_NN4END[5] Tile_X0Y0_E1END[3] Tile_X0Y0_E2END[1] Tile_X0Y0_E6END[1]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q
+ _0700_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5081_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4101_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1792_ _0005_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2293_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ _0102_ _0634_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4032_ _2210_ _2209_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_143_1236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_1225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_regs_0_Tile_X0Y1_UserCLK Tile_X0Y1_UserCLK Tile_X0Y1_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5983_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 net369 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4934_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4865_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_32_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_23 Tile_X0Y1_EE4END[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_12 Tile_X0Y0_W1END[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_56 Tile_X0Y1_N4END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_34 Tile_X0Y1_FrameStrobe[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_45 Tile_X0Y1_N4END[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4796_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3816_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y0_E1END[2] Tile_X0Y0_W1END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q _2041_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_67 Tile_X0Y1_NN4END[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_3747_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q _1442_ _1981_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_89 net365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_78 net378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3678_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1936_ _1937_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput141 net141 Tile_X0Y0_NN4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput130 net130 Tile_X0Y0_N4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput152 net152 Tile_X0Y0_NN4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5417_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2629_ _0937_ _0949_ _0950_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_121_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput174 net174 Tile_X0Y0_W6BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput185 net185 Tile_X0Y0_W6BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5348_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput163 net163 Tile_X0Y0_W2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_322 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput196 net196 Tile_X0Y0_WW4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5279_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_46_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_131_1151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2980_ _1284_ _1288_ _1289_ _1290_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4650_ Tile_X0Y1_N2MID[3] Tile_X0Y1_N4END[7] Tile_X0Y0_E1END[1] Tile_X0Y0_E2END[3]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q
+ _0536_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_12_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3601_ Tile_X0Y0_E2MID[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q _1867_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4581_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q
+ _0471_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3532_ _1774_ _1775_ _1805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3463_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q _1746_ _1747_
+ _0163_ _1748_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5202_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2414_ _0747_ _0748_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5133_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3394_ _1681_ _1682_ _1683_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2345_ _0096_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q _0683_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5064_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_96_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2276_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 _0617_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4015_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ _2195_ _2196_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5966_ Tile_X0Y1_W6END[9] net363 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5897_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 net292 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4917_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_32_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4848_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4779_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_106_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_1206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5820_ Tile_X0Y1_E2MID[1] net215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5751_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A net152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2963_ _1266_ _1272_ _1265_ _1273_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4702_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q _0584_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q
+ _0585_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5682_ Tile_X0Y0_FrameData[28] net69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2894_ _1143_ _1144_ _1205_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4633_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q _0520_ _0521_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_7_Left_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4564_ Tile_X0Y1_N2MID[5] Tile_X0Y1_E2MID[5] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5
+ Tile_X0Y1_W2MID[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q
+ _0455_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3515_ _1762_ _1763_ _1794_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4495_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q _0391_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q
+ _0392_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_110_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3446_ _1729_ _1732_ _1727_ Tile_X0Y1_DSP_bot.C1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3377_ _1665_ _1666_ _0182_ _1664_ _1667_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5116_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_111_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2328_ Tile_X0Y1_N1END[1] Tile_X0Y1_N2END[5] Tile_X0Y1_E1END[1] Tile_X0Y1_E2END[5]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q
+ _0668_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5047_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_84_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5949_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 net344 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_91_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_363 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_1190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_363 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3300_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[8\]
+ _1593_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4280_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q _0184_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3231_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q
+ _1530_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_97_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_399 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3162_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q
+ _1467_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3093_ _0124_ _1402_ _1403_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5803_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 net189 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3995_ _0200_ _1629_ _2177_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q
+ _2178_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_45_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5734_ Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A net135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2946_ _1196_ _1203_ _1256_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5665_ Tile_X0Y0_FrameData[11] net51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_20_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2877_ _0157_ _1188_ _1189_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_100_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4616_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q
+ _0505_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_111_Right_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5596_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4547_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q _0439_ _0440_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4478_ _0370_ _0371_ _0372_ _0373_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q
+ _0375_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_89_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3429_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q _1714_ _1715_
+ _1716_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_79_Left_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_94_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_34_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_88_Left_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3780_ _0456_ Tile_X0Y0_E1END[3] Tile_X0Y0_S1END[3] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q
+ _2010_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_42_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2800_ Tile_X0Y1_N2MID[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q
+ _1114_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2731_ _0150_ _1044_ _1046_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q
+ _1047_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5450_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2662_ Tile_X0Y1_E2MID[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q
+ _0981_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4401_ _0297_ _0298_ _0300_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q _0301_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2593_ _0912_ _0914_ _0915_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5381_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_97_Left_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4332_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q _0232_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q
+ _0235_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4263_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q _0167_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3214_ _0170_ _1506_ _1509_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q
+ _1515_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4194_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q _0098_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3145_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[11\]
+ _1449_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q _1450_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3076_ _1079_ _1384_ _1386_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_94_283 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3978_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ _2162_ _2163_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5717_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 net112 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2929_ _1233_ _1236_ _0131_ _1225_ _1239_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5648_ Tile_X0Y0_EE4END[14] net34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5579_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_105_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_102 Tile_X0Y1_E6END[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_123_1097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_439 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_428 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_1171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4950_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_91_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4881_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3901_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q _2103_ _2105_
+ _2099_ _2101_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3832_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q _2053_ _2054_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3763_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q _1848_ _1994_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q _1995_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5502_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3694_ Tile_X0Y0_S2END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_W2END[1] Tile_X0Y0_W6END[1]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q
+ _1949_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2714_ Tile_X0Y1_N2MID[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q
+ _1031_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_133_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2645_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 _0965_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput301 net301 Tile_X0Y1_S2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5433_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput312 net312 Tile_X0Y1_S4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput334 net334 Tile_X0Y1_W1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput323 net323 Tile_X0Y1_SS4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5364_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput356 net356 Tile_X0Y1_W6BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput367 net367 Tile_X0Y1_WW4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput378 net378 Tile_X0Y1_WW4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput345 net345 Tile_X0Y1_W2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2576_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q _0887_ _0888_
+ _0898_ _0899_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4315_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q
+ _0219_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5295_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_99_375 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4246_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q _0150_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4177_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q _0081_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3128_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y0_E1END[2] Tile_X0Y1_N2MID[6]
+ Tile_X0Y0_E2END[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q _1435_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_35_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3059_ _1367_ _1368_ _1322_ _1369_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2430_ _0758_ _0763_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_450 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2361_ _0092_ _0698_ _0093_ _0699_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5080_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4100_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1788_ _0004_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2292_ _0099_ _0208_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q
+ _0633_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4031_ Tile_X0Y1_N1END[1] Tile_X0Y1_W1END[1] Tile_X0Y1_E1END[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q
+ _2210_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_49_250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_143_1226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5982_ Tile_X0Y1_WW4END[15] net368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_75_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4933_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_52_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4864_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_13 net177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_46 Tile_X0Y1_N4END[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_57 Tile_X0Y1_N4END[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_35 Tile_X0Y1_FrameStrobe[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_3815_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q _2037_ _2039_
+ _2040_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_25_Left_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_24 Tile_X0Y1_EE4END[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4795_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_68 Tile_X0Y1_NN4END[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_79 Tile_X0Y0_E6END[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_3746_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q _0673_ _1979_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q _1980_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5416_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3677_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[19\]
+ _1937_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput142 net142 Tile_X0Y0_NN4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput131 net131 Tile_X0Y0_N4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput120 net120 Tile_X0Y0_N2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_113_1030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2628_ _0600_ _0947_ _0949_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput153 net153 Tile_X0Y0_UserCLKo VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput175 net175 Tile_X0Y0_W6BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5347_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2559_ _0882_ _0883_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput164 net164 Tile_X0Y0_W2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput186 net186 Tile_X0Y0_WW4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5278_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_87_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput197 net197 Tile_X0Y0_WW4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4229_ Tile_X0Y1_E2MID[0] _0133_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_34_Left_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_43_Left_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_120_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_52_Left_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_445 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_72_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4580_ _0464_ _0466_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q
+ _0463_ _0470_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3600_ _0130_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 _1866_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_12_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3531_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1803_ _1804_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3462_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[0\]
+ _1747_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5201_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3393_ _1346_ _1348_ _1357_ _1682_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2413_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q _0745_ _0746_
+ _0747_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5132_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2344_ _0632_ _0633_ _0654_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ _0682_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_29_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2275_ _0611_ _0612_ _0614_ _0616_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5063_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4014_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q _0827_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q
+ _2195_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5965_ Tile_X0Y1_W6END[8] net362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5896_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 net291 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4916_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_138_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4847_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_138_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4778_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3729_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q _1972_ _1970_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_125_Right_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_26_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_60_Left_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_77_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_1207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5750_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A net151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2962_ _1267_ _1268_ _1269_ _1272_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5681_ Tile_X0Y0_FrameData[27] net68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4701_ _0583_ _0584_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4632_ Tile_X0Y0_S1END[1] Tile_X0Y0_W1END[1] Tile_X0Y0_S2END[5] Tile_X0Y0_W1END[3]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q
+ _0520_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2893_ _1196_ _1203_ _1202_ _1204_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4563_ _0454_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3514_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1792_ _1793_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4494_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q _0057_ _0390_
+ _0391_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3445_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q _1730_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q
+ _1732_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3376_ Tile_X0Y1_E2MID[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q _1666_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5115_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2327_ _0658_ _0662_ _0663_ _0664_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q
+ _0667_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XPHY_EDGE_ROW_108_Left_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5046_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_0_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_83_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_351 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 net343 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5879_ Tile_X0Y1_FrameData[24] net266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_117_Left_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_119_361 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_394 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_126_Left_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_370 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3230_ _1524_ _1525_ _1527_ _1529_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3161_ _0119_ _1465_ _1466_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_97_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3092_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q
+ _1402_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_37_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5802_ Tile_X0Y0_WW4END[15] net188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3994_ _0200_ _1707_ _2177_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5733_ Tile_X0Y1_N4END[15] net134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2945_ _1253_ _1254_ _1252_ _1255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5664_ Tile_X0Y0_FrameData[10] net50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_20_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2876_ Tile_X0Y1_N2MID[3] Tile_X0Y1_E2MID[3] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3
+ Tile_X0Y1_W2MID[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q _1188_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5595_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4615_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q
+ _0504_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4546_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q
+ _0439_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_89_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4477_ _0370_ _0371_ _0372_ _0373_ _0374_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3428_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[2\]
+ _1715_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3359_ _0178_ _1649_ _1650_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5029_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_57_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_414 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2730_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q _1045_ _1046_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2661_ Tile_X0Y1_W2MID[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q
+ _0980_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4400_ _0051_ Tile_X0Y1_E2END[1] _0299_ _0300_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2592_ _0074_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q _0913_
+ _0914_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5380_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4331_ _0040_ _0233_ _0234_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4262_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q _0166_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3213_ _1510_ _1511_ _1513_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q _1514_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_86_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4193_ Tile_X0Y0_W2MID[6] _0097_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3144_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q _1448_ _1449_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3075_ _1071_ _1078_ _1384_ _1385_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_50_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3977_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q _1707_ _2162_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5716_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 net111 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2928_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q _1224_ _1234_
+ _1237_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q _1238_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_136_437 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5647_ Tile_X0Y0_EE4END[13] net48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2859_ Tile_X0Y1_N1END[1] Tile_X0Y1_N2END[5] Tile_X0Y1_E1END[1] Tile_X0Y1_E2END[5]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q
+ _1172_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_116_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5578_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4529_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q
+ _0423_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_103 Tile_X0Y1_E6END[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_123_1098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4880_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_17_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3900_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q _2104_ _2105_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3831_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q _1848_ _2052_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q _2053_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3762_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q _0922_ _1994_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5501_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_72_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3693_ _0456_ Tile_X0Y0_E2END[1] Tile_X0Y1_N2MID[1] Tile_X0Y0_E6END[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q _1948_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2713_ Tile_X0Y1_W2MID[5] _0149_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q
+ _1029_ _1030_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2644_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q _0962_ _0964_
+ _0958_ _0960_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5432_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput313 net313 Tile_X0Y1_S4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput335 net335 Tile_X0Y1_W1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput302 net302 Tile_X0Y1_S4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput324 net324 Tile_X0Y1_SS4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5363_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2575_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q _0897_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q
+ _0898_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput357 net357 Tile_X0Y1_W6BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput368 net368 Tile_X0Y1_WW4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput346 net346 Tile_X0Y1_W2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4314_ _0216_ _0217_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q
+ _0218_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput379 net379 Tile_X0Y1_WW4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5294_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4245_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q _0149_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4176_ Tile_X0Y0_WW4END[3] _0080_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3127_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q _1433_ _0123_
+ _1434_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3058_ _1320_ _1321_ _1368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_287 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_446 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2360_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q
+ _0698_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2291_ _0623_ _0626_ _0628_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q
+ _0632_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_10_Right_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4030_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q _2208_ _2206_
+ _2209_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_143_1227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_139_Right_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ Tile_X0Y1_WW4END[14] net367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4932_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_75_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4863_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_32_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_14 net180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_36 Tile_X0Y1_FrameStrobe[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_47 Tile_X0Y1_N4END[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_3814_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q _0875_ _2038_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q _2039_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_15_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_25 Tile_X0Y1_EE4END[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4794_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_58 Tile_X0Y1_N4END[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_69 Tile_X0Y1_NN4END[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_3745_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ _1979_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput110 net110 Tile_X0Y0_N2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5415_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3676_ _1920_ _1935_ _1936_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xoutput143 net143 Tile_X0Y0_NN4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput121 net121 Tile_X0Y0_N4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput132 net132 Tile_X0Y0_N4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_113_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2627_ _0947_ _0948_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput176 net176 Tile_X0Y0_W6BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5346_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2558_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[5\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X
+ _0131_ _0882_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput154 net154 Tile_X0Y0_W1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput165 net165 Tile_X0Y0_W2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput187 net187 Tile_X0Y0_WW4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5277_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2489_ _0116_ _0818_ _0819_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput198 net198 Tile_X0Y0_WW4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4228_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[4\] _0132_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_106_Right_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4159_ Tile_X0Y0_S2MID[7] _0063_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3530_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[11\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ _1804_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3461_ _1746_ Tile_X0Y1_DSP_bot.C0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5200_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3392_ _0163_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[4\] _1680_ _1681_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2412_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[3\]
+ _0746_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5131_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2343_ _0375_ _0377_ _0410_ _0138_ _0681_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_96_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5062_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2274_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q _0615_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q
+ _0616_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4013_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q _1026_ _2193_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q _2194_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_25_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5964_ Tile_X0Y1_W6END[7] net361 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4915_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5895_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 net290 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4846_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4777_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3728_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q _0374_ _1971_
+ _1972_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3659_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[19\]
+ _1919_ _1920_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5329_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_102_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_86_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_287 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_1208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2961_ _1268_ _1269_ _1271_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5680_ Tile_X0Y0_FrameData[26] net67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4700_ Tile_X0Y0_S2END[2] Tile_X0Y0_W2END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_W6END[0]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q
+ _0583_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4631_ _0306_ Tile_X0Y0_E1END[1] Tile_X0Y1_N2MID[5] Tile_X0Y0_E2END[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q _0519_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2892_ _1199_ _1201_ _1203_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_2_0__f_Tile_X0Y1_UserCLK_regs clknet_0_Tile_X0Y1_UserCLK_regs clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4562_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q _0453_ _0450_
+ _0454_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3513_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[5\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ _1793_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4493_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q Tile_X0Y1_N4END[7]
+ _0390_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3444_ _1730_ _1731_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_110_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3375_ Tile_X0Y1_N2MID[7] _0181_ _1665_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5114_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2326_ _0659_ _0661_ _0665_ _0666_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5045_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_83_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5947_ Tile_X0Y1_W2END[4] net342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5878_ Tile_X0Y1_FrameData[23] net265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4829_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_119_1070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3160_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q
+ _1465_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_97_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3091_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 Tile_X0Y0_S2MID[1] Tile_X0Y0_E2MID[1]
+ Tile_X0Y0_W2MID[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q _1401_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_94_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Right_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_80_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5801_ Tile_X0Y0_WW4END[14] net187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5732_ Tile_X0Y1_N4END[14] net133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3993_ _0200_ _0827_ _2175_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q
+ _2176_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2944_ _1249_ _1250_ _1254_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5663_ Tile_X0Y0_FrameData[9] net80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_20_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2875_ _1183_ _1184_ _1186_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q
+ _0157_ _1187_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5594_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4614_ _0502_ _0503_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4545_ _0437_ _0438_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4476_ _0085_ Tile_X0Y0_W2MID[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q
+ _0373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3427_ _1714_ Tile_X0Y1_DSP_bot.C2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_39_Right_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3358_ Tile_X0Y1_N2MID[2] Tile_X0Y1_W2MID[2] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q _1649_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_97_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2309_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q _0617_ _0648_
+ _0649_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3289_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q
+ _1584_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5028_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_48_Right_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_139_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Right_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_79_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_66_Right_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2660_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q _0956_ _0979_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2591_ Tile_X0Y0_S2MID[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q _0913_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_75_Right_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4330_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q
+ _0233_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_125_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4261_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q _0165_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3212_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ _1512_ _1513_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4192_ Tile_X0Y1_W1END[1] _0096_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3143_ _1448_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3074_ _1381_ _1383_ _1384_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_84_Right_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_285 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3976_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q _1629_ _2160_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q _2161_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5715_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 net110 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2927_ _1233_ _1236_ _1225_ Tile_X0Y1_DSP_bot.B0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5646_ Tile_X0Y0_EE4END[12] net47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2858_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q _1166_ _1167_
+ _1170_ _1171_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XPHY_EDGE_ROW_93_Right_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2789_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ _1104_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5577_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4528_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q
+ _0422_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_116_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4459_ Tile_X0Y1_N1END[2] Tile_X0Y1_E1END[2] Tile_X0Y1_N2END[6] Tile_X0Y1_E2END[6]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_49_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_104 Tile_X0Y1_N4END[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_1099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3830_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q _0594_ _2052_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3761_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q _1420_ _1992_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q _1993_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5500_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2712_ _0149_ _0454_ _1029_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3692_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1946_ _1947_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2643_ _0145_ _0963_ _0964_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5431_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_65_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput303 net303 Tile_X0Y1_S4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput325 net325 Tile_X0Y1_SS4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput314 net314 Tile_X0Y1_S4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5362_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2574_ Tile_X0Y0_W2MID[6] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q
+ _0897_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput358 net358 Tile_X0Y1_W6BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput369 net369 Tile_X0Y1_WW4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput336 net336 Tile_X0Y1_W1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput347 net347 Tile_X0Y1_W2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4313_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ _0217_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5293_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4244_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q _0148_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_316 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4175_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q _0079_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3126_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q
+ _1433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3057_ _1361_ _1363_ _1336_ _1367_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3959_ Tile_X0Y1_N1END[3] Tile_X0Y1_E1END[3] _0412_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q
+ _2146_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5629_ Tile_X0Y0_E6END[5] net26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_377 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2290_ _0624_ _0625_ _0629_ _0099_ _0631_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_96_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_143_1228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5980_ Tile_X0Y1_WW4END[13] net381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4931_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_75_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4862_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3813_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q _1879_ _2038_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_37 Tile_X0Y1_FrameStrobe[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_48 Tile_X0Y1_N4END[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_15 net183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_26 Tile_X0Y1_EE4END[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4793_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_59 Tile_X0Y1_NN4END[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_3744_ _1978_ _1977_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3675_ _1836_ _1930_ _1933_ _1934_ _1935_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xoutput100 net100 Tile_X0Y0_FrameStrobe_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5414_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2626_ _0938_ _0945_ _0947_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput122 net122 Tile_X0Y0_N4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput133 net133 Tile_X0Y0_N4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput111 net111 Tile_X0Y0_N2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput144 net144 Tile_X0Y0_NN4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2557_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q _0877_ _0878_
+ _0881_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_113_1032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5345_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput155 net155 Tile_X0Y0_W1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput166 net166 Tile_X0Y0_W2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput177 net177 Tile_X0Y0_W6BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput199 net199 Tile_X0Y0_WW4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5276_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2488_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 Tile_X0Y0_S2MID[5] Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_W2MID[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q _0818_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput188 net188 Tile_X0Y0_WW4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4227_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q _0131_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4158_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q _0062_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4089_ _0205_ _2260_ _2261_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3109_ _1379_ _1387_ _1417_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_55_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3460_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q _1745_ _1743_
+ _1746_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3391_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q _1678_ _1679_
+ _0163_ _1680_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2411_ _0745_ Tile_X0Y1_DSP_bot.A3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5130_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_123_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2342_ _0679_ _0680_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5061_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_336 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2273_ Tile_X0Y0_S2END[4] Tile_X0Y0_W2END[4] Tile_X0Y0_S4END[0] Tile_X0Y0_WW4END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ _0615_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4012_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q _1689_ _2193_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5963_ Tile_X0Y1_W6END[6] net360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4914_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5894_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 net289 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4845_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4776_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_20_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3727_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q _0210_ _1971_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3658_ _1917_ _1918_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q
+ _1919_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3589_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[16\]
+ _1857_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2609_ _0849_ _0929_ _0930_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5328_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5259_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_86_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_140_1209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2960_ _0679_ _1242_ _1268_ _1270_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_42_280 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2891_ _1200_ _1201_ _1202_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4630_ _0110_ _0511_ _0517_ _0518_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4561_ _0451_ _0452_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q
+ _0453_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3512_ _1760_ _1761_ _1792_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4492_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q _0388_ _0389_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3443_ Tile_X0Y1_N2MID[3] Tile_X0Y1_E2MID[3] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3
+ Tile_X0Y1_W2MID[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q _1730_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5113_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_110_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3374_ _0181_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 _1663_ _1664_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2325_ _0663_ _0664_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q
+ _0665_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5044_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_83_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5946_ Tile_X0Y1_W2END[3] net341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5877_ Tile_X0Y1_FrameData[22] net264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4828_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_23_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4759_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_119_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_435 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Left_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3090_ _0529_ _1389_ _1397_ _1400_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_66_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3992_ _0200_ _1026_ _2175_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_80_819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5800_ Tile_X0Y0_WW4END[13] net201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5731_ Tile_X0Y1_N4END[13] net132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2943_ _1220_ _1246_ _1245_ _1253_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5662_ Tile_X0Y0_FrameData[8] net79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_20_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2874_ Tile_X0Y1_E2MID[2] _0154_ _1185_ _1186_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5593_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4613_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q _0501_ _0502_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4544_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q
+ _0437_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_143_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q Tile_X0Y0_S2MID[5]
+ _0372_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3426_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q _1713_ _1703_
+ _1714_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3357_ _0178_ _1646_ _0179_ _1648_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2308_ Tile_X0Y0_W2END[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q _0648_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5027_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3288_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q
+ _1583_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5929_ Tile_X0Y0_SS4END[14] net330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_1126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_1200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_57_Left_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_287 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2590_ _0071_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q
+ _0911_ _0912_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_140_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4260_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[10\] _0164_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3211_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q _0212_ _1512_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4191_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q _0095_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3142_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q _1444_ _1447_
+ _1448_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_66_Left_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3073_ _1073_ _1382_ _1383_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_93_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3975_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q _1094_ _2160_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5714_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 net109 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2926_ _1236_ _1237_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5645_ Tile_X0Y0_EE4END[11] net46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2857_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q _1169_ _1170_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2788_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q _1103_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5576_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4527_ _0421_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_116_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4458_ _0352_ _0353_ _0354_ _0355_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q
+ _0356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3409_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[3\]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q _1697_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4389_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q
+ _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_105 Tile_X0Y1_N4END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3760_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ _1992_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2711_ _1019_ _1021_ _1024_ _0150_ _1028_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3691_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[8\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ _1947_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5430_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_72_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2642_ Tile_X0Y1_E6END[0] Tile_X0Y1_W2END[2] Tile_X0Y0_S2MID[2] Tile_X0Y1_WW4END[3]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q
+ _0963_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2573_ _0890_ _0892_ _0894_ _0896_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5361_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput315 net315 Tile_X0Y1_S4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput304 net304 Tile_X0Y1_S4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput326 net326 Tile_X0Y1_SS4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput359 net359 Tile_X0Y1_W6BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput337 net337 Tile_X0Y1_W1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput348 net348 Tile_X0Y1_W2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5292_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4312_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ _0216_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_99_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4243_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q _0147_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4174_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q _0078_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3125_ _0122_ _1431_ _1432_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3056_ _1362_ _1364_ _1335_ _1366_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3958_ _2145_ _2144_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_61_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3889_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 _0272_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0
+ _0286_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2909_ _0680_ _1194_ _1220_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5628_ Tile_X0Y0_E6END[4] net25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5559_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_132_431 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_1107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_143_1229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4930_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4861_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3812_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ _2036_ _2037_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_50_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_38 Tile_X0Y1_FrameStrobe[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_120_Right_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_27 Tile_X0Y1_EE4END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4792_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_16 net196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_49 Tile_X0Y1_N4END[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_3743_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y0_E1END[2] Tile_X0Y0_W1END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q _1978_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3674_ _1836_ _1931_ _1934_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput101 net101 Tile_X0Y0_N1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5413_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2625_ _0938_ _0945_ _0946_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput123 net123 Tile_X0Y0_N4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput134 net134 Tile_X0Y0_N4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput112 net112 Tile_X0Y0_N2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5344_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput145 net145 Tile_X0Y0_NN4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2556_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q _0879_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q
+ _0881_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_113_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput156 net156 Tile_X0Y0_W1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput167 net167 Tile_X0Y0_W2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput178 net178 Tile_X0Y0_W6BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5275_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2487_ _0812_ _0814_ _0116_ _0811_ _0817_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xoutput189 net189 Tile_X0Y0_WW4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4226_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q _0130_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4157_ Tile_X0Y0_E2MID[7] _0061_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3108_ _0163_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[13\] _1413_ _1415_ _1416_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4088_ Tile_X0Y1_W2MID[0] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q _2260_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3039_ _1347_ _1348_ _1349_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_12_Left_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_127_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_21_Left_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_46_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Left_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2410_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q _0744_ _0732_
+ _0745_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3390_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[4\]
+ _1679_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2341_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q _0677_ _0678_
+ _0679_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5060_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2272_ _0069_ _0613_ _0614_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4011_ _2192_ _2191_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ Tile_X0Y1_W6END[5] net359 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4913_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5893_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 net288 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4844_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4775_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3726_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2
+ _1969_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q _1970_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3657_ _0162_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X
+ _1918_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2608_ _0776_ _0907_ _0929_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3588_ _1854_ _1855_ _1856_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_121_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2539_ _0863_ _0865_ _0861_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5327_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_87_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5258_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4209_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q _0113_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5189_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X
+ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[19\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2890_ _1139_ _1140_ _1201_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4560_ Tile_X0Y0_S1END[2] Tile_X0Y0_S2END[6] Tile_X0Y0_W1END[0] Tile_X0Y0_W1END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q
+ _0452_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_8_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3511_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1790_ _1791_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4491_ Tile_X0Y1_N2MID[3] _0056_ _0388_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3442_ _0187_ _1728_ _1729_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3373_ _0048_ _0181_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q
+ _1663_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5112_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_110_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2324_ Tile_X0Y1_W1END[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q _0664_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5043_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_83_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5945_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 net340 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5876_ Tile_X0Y1_FrameData[21] net263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4827_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_23_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_432 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4758_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_119_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3709_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 _0482_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3
+ _0468_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4689_ _0571_ _0572_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_421 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_432 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3991_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q _2168_ _2170_
+ _2172_ _2174_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5730_ Tile_X0Y1_N4END[12] net131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2942_ _1249_ _1251_ _1252_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5661_ Tile_X0Y0_FrameData[7] net78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2873_ Tile_X0Y1_N2MID[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q
+ _1185_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_88_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5592_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4612_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q _0500_ _0501_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4543_ Tile_X0Y1_NN4END[3] Tile_X0Y1_WW4END[0] Tile_X0Y0_S4END[7] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q
+ _0436_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_143_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4474_ Tile_X0Y0_E2MID[5] _0085_ _0086_ _0371_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3425_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q _1707_ _1712_
+ _1713_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3356_ _1646_ _1647_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3287_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4
+ _1581_ _1582_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2307_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0
+ _0647_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5026_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_57_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5928_ Tile_X0Y0_SS4END[13] net329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5859_ Tile_X0Y1_FrameData[4] net276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_128_1127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_1201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Left_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_113_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_326 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4190_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q _0094_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3210_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q _1511_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3141_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q _1442_ _1446_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q _1447_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_79_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3072_ _0598_ _0824_ _1382_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_93_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3974_ _2154_ _2157_ _2159_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5713_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 net108 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2925_ _0159_ _1235_ _0160_ _1236_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5644_ Tile_X0Y0_EE4END[10] net45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2856_ Tile_X0Y0_S2MID[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q _1168_ _1169_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2787_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q
+ _1102_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5575_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_116_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4526_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q _0218_ _0417_
+ _0420_ _0421_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4457_ Tile_X0Y1_W1END[2] _0078_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q
+ _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3408_ _0162_ Tile_X0Y1_DSP_bot.C3 _1696_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4388_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q _0287_ _0288_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3339_ Tile_X0Y1_W2MID[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q
+ _1631_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_134_Right_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_106 Tile_X0Y1_NN4END[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5009_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_56_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_287 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_101_Right_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_17_332 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2710_ _1020_ _1022_ _1025_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q
+ _1027_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3690_ _1945_ _1946_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2641_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q _0961_ _0962_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2572_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q _0895_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q
+ _0896_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5360_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput316 net316 Tile_X0Y1_S4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput305 net305 Tile_X0Y1_S4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4311_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 _0215_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput349 net349 Tile_X0Y1_W2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput327 net327 Tile_X0Y1_SS4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput338 net338 Tile_X0Y1_W2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5291_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4242_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[1\] _0146_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4173_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q _0077_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3124_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q
+ _1431_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3055_ _1362_ _1364_ _1365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_55_449 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_53_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_324 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_122_1090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3957_ Tile_X0Y1_N1END[2] Tile_X0Y1_E1END[2] _0351_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q
+ _2145_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2908_ _1216_ _1217_ _1219_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_61_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3888_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 _0254_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3
+ _0231_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5627_ Tile_X0Y0_E6END[3] net24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2839_ _0927_ _1053_ _1152_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5558_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4509_ Tile_X0Y0_E6END[0] Tile_X0Y0_W2END[2] Tile_X0Y0_S2END[2] Tile_X0Y0_W6END[0]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q
+ _0405_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5489_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_18_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_1108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_85_Left_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Left_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_432 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4860_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3811_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q _0916_ _2036_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_39 Tile_X0Y1_FrameStrobe[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4791_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_28 Tile_X0Y1_EE4END[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_17 net197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_3742_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q _1974_ _1976_
+ _1977_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_15_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3673_ _1884_ _1929_ _1931_ _1933_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5412_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2624_ _0939_ _0943_ _0945_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput113 net113 Tile_X0Y0_N2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput124 net124 Tile_X0Y0_N4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput102 net102 Tile_X0Y0_N1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5343_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput135 net135 Tile_X0Y0_N4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput146 net146 Tile_X0Y0_NN4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2555_ _0879_ _0880_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_443 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput157 net157 Tile_X0Y0_W1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput168 net168 Tile_X0Y0_W2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2486_ _0815_ _0816_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5274_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput179 net179 Tile_X0Y0_W6BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4225_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q _0129_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4156_ Tile_X0Y1_W1END[0] _0060_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3107_ _0163_ _1414_ _1415_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4087_ Tile_X0Y1_N2MID[6] Tile_X0Y1_E2MID[0] Tile_X0Y1_E2MID[6] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q
+ _2259_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3038_ _1328_ _1332_ _1348_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_70_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4989_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_105_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2340_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[6\]
+ _0678_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2271_ Tile_X0Y1_N2MID[4] Tile_X0Y0_E2END[4] Tile_X0Y0_E1END[2] Tile_X0Y0_E6END[0]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ _0613_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4010_ Tile_X0Y1_N1END[2] Tile_X0Y1_E1END[2] Tile_X0Y1_W1END[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q
+ _2192_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5961_ Tile_X0Y1_W6END[4] net358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4912_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5892_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 net287 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4843_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4774_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_20_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3725_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q _0408_ _1969_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3656_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[19\]
+ _1917_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2607_ _0882_ _0927_ _0928_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3587_ _1399_ _1779_ _1833_ _1832_ _1855_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2538_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q _0864_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q
+ _0865_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5326_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5257_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2469_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ _0800_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4208_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q _0112_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5188_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X
+ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[18\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4139_ Tile_X0Y1_E2END[3] _0043_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_86_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_385 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3510_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[3\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ _1791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4490_ _0273_ _0277_ _0305_ _0056_ _0387_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3441_ Tile_X0Y1_N2MID[2] Tile_X0Y1_E2MID[2] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q _1728_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3372_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q _1659_ _1660_
+ _1661_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q _1662_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5111_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_110_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2323_ Tile_X0Y1_W1END[3] _0098_ _0663_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5042_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5944_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 net339 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5875_ Tile_X0Y1_FrameData[20] net262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4826_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4757_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3708_ Tile_X0Y1_N2MID[1] Tile_X0Y0_W6END[0] Tile_X0Y1_N4END[4] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_119_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4688_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 Tile_X0Y0_S2MID[1] Tile_X0Y0_E2MID[1]
+ Tile_X0Y0_W2MID[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q
+ _0571_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3639_ _1895_ _1901_ _1902_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q
+ _1903_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_99_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_363 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_399 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_433 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3990_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q _2173_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q
+ _2174_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2941_ _1250_ _1251_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5660_ Tile_X0Y0_FrameData[6] net77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2872_ Tile_X0Y1_W2MID[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q _1184_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4611_ Tile_X0Y1_N1END[0] Tile_X0Y1_E1END[0] Tile_X0Y1_N2END[0] Tile_X0Y1_EE4END[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q
+ _0500_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_100_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5591_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_128_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4542_ _0428_ _0435_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4473_ _0356_ _0359_ _0365_ _0368_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q
+ _0370_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_143_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3424_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q _1711_ _1710_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q _1712_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_89_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_115_Right_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3355_ Tile_X0Y1_N2END[3] Tile_X0Y1_E2END[3] Tile_X0Y0_SS4END[4] Tile_X0Y1_W2END[3]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q
+ _1646_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2306_ _0644_ _0646_ _0642_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3286_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q _0672_ _0171_
+ _1581_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_96_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5025_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_36_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5927_ Tile_X0Y0_SS4END[12] net328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_449 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5858_ Tile_X0Y1_FrameData[3] net275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5789_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 net175 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4809_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_17_Right_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_119_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Right_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_1128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_1202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_35_Right_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_42_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Right_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3140_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q _1445_ _1446_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_105_Left_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3071_ _0940_ _1072_ _1076_ _1381_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_93_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_322 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5712_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 net107 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_53_Right_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3973_ _2158_ _2159_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_114_Left_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2924_ Tile_X0Y1_N2MID[7] Tile_X0Y1_E2MID[7] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7
+ Tile_X0Y1_W2MID[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q
+ _1235_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5643_ Tile_X0Y0_EE4END[9] net44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2855_ _0096_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q _1168_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5574_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2786_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q _1100_ _1098_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q _1101_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4525_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q _0419_ _0420_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_116_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_62_Right_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4456_ Tile_X0Y1_W1END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ _0354_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_123_Left_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4387_ _0286_ _0287_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3407_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q _1691_ _1693_
+ _1695_ Tile_X0Y1_DSP_bot.C3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3338_ Tile_X0Y1_N2MID[5] Tile_X0Y1_E2MID[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q
+ _1630_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3269_ Tile_X0Y1_E1END[3] _0172_ _1565_ _1566_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_107 net373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_5008_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_56_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_71_Right_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_132_Left_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_139_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_80_Right_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_141_Left_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_134_1165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2640_ Tile_X0Y1_N1END[0] Tile_X0Y1_N2END[2] Tile_X0Y1_N4END[2] Tile_X0Y1_E2END[2]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q
+ _0961_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2571_ Tile_X0Y0_E6END[0] Tile_X0Y0_S2END[4] Tile_X0Y0_W2END[4] Tile_X0Y0_W6END[0]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q
+ _0895_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput317 net317 Tile_X0Y1_S4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput306 net306 Tile_X0Y1_S4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4310_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 _0214_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput339 net339 Tile_X0Y1_W2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput328 net328 Tile_X0Y1_SS4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5290_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_141_433 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4241_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q _0145_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4172_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q _0076_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3123_ _1429_ _1430_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3054_ _1333_ _1334_ _1364_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_1091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3956_ _2141_ _2143_ _2144_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2907_ _1216_ _1217_ _1218_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5626_ Tile_X0Y0_E6END[2] net21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3887_ Tile_X0Y1_N2END[1] Tile_X0Y1_N4END[0] Tile_X0Y1_W6END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q
+ Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2838_ _1149_ _1150_ _1151_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5557_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2769_ _1081_ _1082_ _1084_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4508_ _0087_ _0403_ _0404_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5488_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4439_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q
+ _0338_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_76_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_1109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3810_ _2030_ _2035_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4790_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_29 Tile_X0Y1_FrameStrobe[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_3741_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q _0875_ _1975_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q _1976_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_32_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_18 net199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3672_ _1884_ _1931_ _1932_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5411_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_63_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2623_ _0939_ _0943_ _0944_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput125 net125 Tile_X0Y0_N4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput103 net103 Tile_X0Y0_N1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput114 net114 Tile_X0Y0_N2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2554_ Tile_X0Y1_N2MID[2] Tile_X0Y0_S2END[2] Tile_X0Y0_E2END[2] Tile_X0Y0_WW4END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q
+ _0879_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5342_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput147 net147 Tile_X0Y0_NN4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput136 net136 Tile_X0Y0_N4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput158 net158 Tile_X0Y0_W2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5273_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2485_ _0812_ _0814_ _0811_ _0815_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput169 net169 Tile_X0Y0_W2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4224_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q _0128_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4155_ Tile_X0Y0_W2END[3] _0059_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3106_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[13\]
+ _1414_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4086_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q _0204_ _2258_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3037_ _1346_ _1347_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4988_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3939_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q _1725_ _2130_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5609_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_1146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_447 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_142_1220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_431 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2270_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q _0609_ _0070_
+ _0612_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5960_ Tile_X0Y1_W6END[3] net357 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4911_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5891_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 net286 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4842_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4773_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_9_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3724_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 _0346_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1
+ _0321_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3655_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q _1910_ _1916_
+ _1904_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2606_ _0926_ _0927_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3586_ _1836_ _1852_ _1854_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2537_ Tile_X0Y0_S1END[1] Tile_X0Y0_S2END[5] Tile_X0Y0_S1END[3] Tile_X0Y0_W1END[1]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q
+ _0864_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5325_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2468_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ _0798_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q _0799_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5256_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_87_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4207_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q _0111_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2399_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q
+ _0735_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5187_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X
+ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[17\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4138_ Tile_X0Y1_N4END[3] _0042_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4069_ _0202_ _2242_ _2243_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_129_Right_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_105_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_364 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3440_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q _1721_ _1726_
+ _1727_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3371_ Tile_X0Y1_E2MID[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q _1661_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5110_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_111_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2322_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q _0660_ _0662_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5041_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_57_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5943_ Tile_X0Y1_W2END[0] net338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_103_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5874_ Tile_X0Y1_FrameData[19] net260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4825_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4756_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3707_ Tile_X0Y1_N2MID[0] Tile_X0Y1_N4END[7] Tile_X0Y0_W6END[1] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4687_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 Tile_X0Y0_E2MID[0] Tile_X0Y0_S2MID[0]
+ _0561_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q
+ _0570_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3638_ _0190_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 _1902_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3569_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4
+ _1838_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5308_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_142_391 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5239_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_102_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_1185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_2_3__f_Tile_X0Y1_UserCLK_regs clknet_0_Tile_X0Y1_UserCLK_regs clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_18_Left_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_66_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_27_Left_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2940_ _1160_ _1161_ _1197_ _1250_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2871_ _1171_ _1174_ _1178_ _1181_ _0154_ _1183_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_30_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4610_ _0490_ _0494_ _0495_ _0496_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q
+ _0499_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_100_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5590_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4541_ _0024_ _0434_ _0433_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q
+ _0435_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_128_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Left_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4472_ _0360_ _0369_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3423_ Tile_X0Y1_N2MID[5] Tile_X0Y1_E2MID[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q
+ _1711_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3354_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q _1644_ _1643_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q _1645_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2305_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q _0645_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q
+ _0646_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3285_ _0171_ _1579_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q
+ _1580_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_96_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_57_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5926_ Tile_X0Y0_SS4END[11] net327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5857_ Tile_X0Y1_FrameData[2] net272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5788_ Tile_X0Y0_W6END[11] net185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4808_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4739_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_107_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_1129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_59_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_1203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_441 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3070_ _1083_ _1086_ _1380_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5711_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 net106 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_33_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3972_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 _1651_ _1730_ _1222_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q _2158_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_93_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2923_ _1226_ _1228_ _1232_ _1234_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5642_ Tile_X0Y0_EE4END[8] net43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2854_ _0632_ _0633_ _0654_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ _1167_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5573_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2785_ Tile_X0Y1_N2MID[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q
+ _1099_ _1100_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4524_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q _0418_ _0419_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4455_ _0078_ Tile_X0Y0_S2MID[6] _0079_ _0353_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4386_ Tile_X0Y1_N4END[1] Tile_X0Y0_SS4END[5] Tile_X0Y1_W2END[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q
+ _0286_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3406_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q _1694_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q
+ _1695_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3337_ Tile_X0Y1_E2MID[4] Tile_X0Y1_W2MID[4] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q _1629_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3268_ Tile_X0Y1_E2END[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ _1565_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3199_ Tile_X0Y1_W1END[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q
+ _1500_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5007_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_108 net374 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5909_ Tile_X0Y0_S4END[10] net310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_134_1166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_47_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2570_ _0089_ _0893_ _0894_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput307 net307 Tile_X0Y1_S4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput329 net329 Tile_X0Y1_SS4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput318 net318 Tile_X0Y1_SS4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4240_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q _0144_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4171_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q _0075_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3122_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 Tile_X0Y0_E2MID[3] Tile_X0Y0_S2MID[3]
+ Tile_X0Y0_W2MID[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q _1429_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_67_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3053_ _1333_ _1334_ _1363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_23_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3955_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q _1188_ _2142_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q _2143_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_122_1092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2906_ _1149_ _1150_ _1157_ _1217_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_61_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5625_ Tile_X0Y0_E2MID[7] net20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3886_ Tile_X0Y1_N2END[0] Tile_X0Y1_N4END[3] Tile_X0Y1_W6END[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q
+ Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2837_ _1124_ _1125_ _1150_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5556_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2768_ _1079_ _1080_ _1082_ _1083_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4507_ Tile_X0Y1_N2MID[2] Tile_X0Y0_E1END[0] Tile_X0Y1_N4END[6] Tile_X0Y0_E2END[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q
+ _0403_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5487_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2699_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q _1016_ _1015_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q _1017_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4438_ _0322_ _0336_ _0337_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4369_ _0032_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q _0270_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_307 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3740_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q _1825_ _1975_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_19 Tile_X0Y1_E6END[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3671_ _1854_ _1855_ _1883_ _1836_ _1853_ _1931_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5410_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2622_ _0929_ _0941_ _0943_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput115 net115 Tile_X0Y0_N2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput104 net104 Tile_X0Y0_N1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2553_ _0114_ _0468_ _0878_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5341_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_141_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput137 net137 Tile_X0Y0_NN4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput126 net126 Tile_X0Y0_N4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput148 net148 Tile_X0Y0_NN4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput159 net159 Tile_X0Y0_W2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5272_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2484_ _0813_ _0814_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4223_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q _0127_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4154_ Tile_X0Y0_E6END[1] _0058_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4085_ _2250_ _2257_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3105_ _0162_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X
+ _1413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3036_ _1340_ _1343_ _1337_ _1346_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4987_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3938_ _2129_ _2128_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q
+ Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3869_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q _2079_ _2081_
+ _2083_ _2085_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5608_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5539_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_131_1147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_1221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_426 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4910_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5890_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 net285 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4841_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_60_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4772_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_20_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3723_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 _0630_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0
+ _0653_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3654_ _0190_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 _1915_ _0191_ _1916_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2605_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[5\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q
+ _0925_ _0926_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3585_ _1836_ _1852_ _1853_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2536_ _0113_ _0862_ _0863_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5324_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2467_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q _0208_ _0798_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5255_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4206_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q _0110_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2398_ _0135_ _0733_ _0734_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_3_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5186_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X
+ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[16\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4137_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q _0041_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_332 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4068_ _0955_ _1188_ _1730_ _1651_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q _2242_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3019_ _1326_ _1327_ _1329_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_106_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3370_ Tile_X0Y1_N2MID[6] _0180_ _1660_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2321_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q _0660_ _0661_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5040_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5942_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 net337 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5873_ Tile_X0Y1_FrameData[18] net259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_91_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4824_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_103_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4755_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3706_ Tile_X0Y1_N2MID[3] Tile_X0Y1_N4END[6] Tile_X0Y0_E6END[0] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4686_ _0563_ _0565_ _0567_ _0569_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_31_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3637_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q _1900_ _1901_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3568_ _0163_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[16\] _1837_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5307_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2519_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q _0843_ _0845_
+ _0846_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3499_ _1752_ _1753_ _1783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_99_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5238_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_102_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5169_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X
+ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[7\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_446 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_1186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2870_ _1175_ _1182_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_100_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4540_ Tile_X0Y1_N2END[2] Tile_X0Y1_N4END[2] Tile_X0Y1_E1END[0] Tile_X0Y1_E2END[2]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q
+ _0434_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_143_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4471_ _0365_ _0368_ _0369_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3422_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q _0454_ _1709_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q _1710_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_143_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3353_ Tile_X0Y1_N4END[2] Tile_X0Y0_SS4END[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q
+ _1644_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2304_ Tile_X0Y0_E6END[1] Tile_X0Y0_S2END[1] Tile_X0Y0_W2END[1] Tile_X0Y0_W6END[1]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q
+ _0645_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3284_ _0177_ _1578_ _1569_ _1579_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5023_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_96_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5925_ Tile_X0Y0_SS4END[10] net326 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5856_ Tile_X0Y1_FrameData[1] net261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4807_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_3_Right_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5787_ Tile_X0Y0_W6END[10] net184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2999_ _0907_ _1238_ _1241_ _1309_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_119_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4738_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_119_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4669_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q
+ _0553_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_135_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_0__f_Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK clknet_1_0__leaf_Tile_X0Y1_UserCLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3971_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q _2156_ _2157_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5710_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 net105 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_33_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2922_ _1227_ _1229_ _1231_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q
+ _1233_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5641_ Tile_X0Y0_EE4END[7] net42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2853_ _0375_ _0377_ _0410_ _0155_ _1166_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5572_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2784_ _0032_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q _1099_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4523_ Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[7] Tile_X0Y1_E1END[3] Tile_X0Y1_E2END[7]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ _0418_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_104_307 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4454_ _0322_ _0336_ _0350_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ _0352_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_131_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4385_ _0279_ _0281_ _0283_ _0285_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3405_ Tile_X0Y1_N2MID[1] Tile_X0Y1_E2MID[1] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1
+ Tile_X0Y1_W2MID[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q _1694_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3336_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q _1626_ _1625_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q _1628_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_0_Left_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3267_ Tile_X0Y1_N2END[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q _1564_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5006_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_38_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3198_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q _0488_ _1498_
+ _1499_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_109 net380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5908_ Tile_X0Y0_S4END[9] net309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5839_ Tile_X0Y1_EE4END[4] net234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_1167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_55_Left_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_76_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_441 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput308 net308 Tile_X0Y1_S4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput319 net319 Tile_X0Y1_SS4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4170_ Tile_X0Y0_W2MID[3] _0074_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3121_ _0163_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[11\] _1428_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3052_ _1358_ _1359_ _1350_ _1362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3954_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q _1676_ _2142_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_122_1093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3885_ Tile_X0Y1_N2END[3] Tile_X0Y1_E6END[0] Tile_X0Y1_N4END[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q
+ Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2905_ _1209_ _1215_ _1216_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5624_ Tile_X0Y0_E2MID[6] net19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2836_ _0990_ _1148_ _1149_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5555_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2767_ _0600_ _0948_ _0946_ _1082_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4506_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q _0401_ _0088_
+ _0402_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5486_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2698_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q
+ _1016_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4437_ _0082_ _0335_ _0336_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4368_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q _0262_ _0267_
+ _0268_ _0269_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4299_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q _0203_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3319_ Tile_X0Y1_W2MID[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q
+ _1611_ _1612_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_63_Left_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_72_Left_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3670_ _1929_ _1930_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2621_ _0929_ _0941_ _0942_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput116 net116 Tile_X0Y0_N2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput105 net105 Tile_X0Y0_N2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2552_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q _0874_ _0876_
+ _0877_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5340_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput149 net149 Tile_X0Y0_NN4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput127 net127 Tile_X0Y0_N4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput138 net138 Tile_X0Y0_NN4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5271_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_49_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_81_Left_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4222_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q _0126_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2483_ _0103_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q
+ _0813_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4153_ Tile_X0Y0_E2END[3] _0057_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4084_ _2252_ _2255_ _2256_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q _2257_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3104_ _1411_ _1410_ _1401_ _1412_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_95_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_385 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_1100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3035_ _1324_ _1329_ _1344_ _1345_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_66_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_90_Left_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4986_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3937_ Tile_X0Y1_N1END[2] Tile_X0Y1_E1END[2] Tile_X0Y1_W1END[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q
+ _2129_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3868_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q _2084_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q
+ _2085_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5607_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3799_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q _0816_ _2024_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q _2025_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2819_ _0719_ _0720_ _0907_ _1132_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5538_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_105_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_1148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5469_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_78_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_449 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_129_Left_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_142_1222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_138_Left_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4840_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_28_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4771_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3722_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q _1968_ _1963_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3653_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7
+ _1915_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2604_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q _0924_ _0925_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5323_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3584_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q _1851_ _1837_
+ _1852_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2535_ _0306_ Tile_X0Y0_E1END[1] Tile_X0Y1_N2MID[5] Tile_X0Y0_E2END[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q _0862_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_143_Right_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2466_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q
+ _0797_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5254_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_87_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4205_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q _0109_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5185_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X
+ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[15\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4136_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q _0040_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_3_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2397_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q
+ _0733_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4067_ _0202_ _2240_ _2241_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3018_ _1326_ _1327_ _1328_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_106_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_433 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4969_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_138_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_110_Right_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_85_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_425 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2320_ Tile_X0Y0_S2MID[5] _0098_ _0660_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5941_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 net336 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5872_ Tile_X0Y1_FrameData[17] net258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_91_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4823_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4754_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3705_ Tile_X0Y1_N2MID[2] Tile_X0Y1_N4END[5] Tile_X0Y0_E6END[1] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4685_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q _0568_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q
+ _0569_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_31_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3636_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q _1897_ _1899_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q _1900_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3567_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q _1811_ _1836_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5306_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2518_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[2\]
+ _0845_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5237_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3498_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1781_ _1782_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_99_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2449_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ _0780_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q _0781_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_68_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5168_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X
+ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[6\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4119_ Tile_X0Y1_W2END[2] _0023_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_39_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5099_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_17_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_1187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4470_ _0084_ _0367_ _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3421_ Tile_X0Y1_W2MID[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q
+ _1709_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3352_ _0023_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q
+ _1642_ _1643_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2303_ _0101_ _0643_ _0644_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3283_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 _1578_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5022_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_96_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5924_ Tile_X0Y0_SS4END[9] net325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5855_ Tile_X0Y1_FrameData[0] net250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4806_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2998_ _1282_ _1307_ _1308_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5786_ Tile_X0Y0_W6END[9] net183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4737_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_119_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4668_ _0551_ _0552_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3619_ _1836_ _1883_ _1884_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4599_ _0470_ _0480_ _0486_ _0488_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Right_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3970_ _0021_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q
+ _2155_ _2156_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2921_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q _1231_ _1232_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5640_ Tile_X0Y0_EE4END[6] net41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2852_ _0231_ _1164_ _0157_ _1165_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_22_Right_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5571_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2783_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7
+ _1097_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q _1098_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_79_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4522_ _0413_ _0414_ _0415_ _0416_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q
+ _0417_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4453_ _0337_ _0349_ _0351_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3404_ _0184_ _1692_ _1693_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4384_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q _0284_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q
+ _0285_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3335_ _1626_ _1627_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_31_Right_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3266_ Tile_X0Y1_N1END[3] _0172_ _1563_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5005_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_85_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_1120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3197_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q _0351_ _1498_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5907_ Tile_X0Y0_S4END[8] net302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5838_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 net224 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_40_Right_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5769_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 net164 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_101_Left_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_135_400 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_1168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_110_Left_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_49_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput309 net309 Tile_X0Y1_S4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3120_ _1425_ _1426_ _1427_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3051_ _1357_ _1360_ _1349_ _1361_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3953_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ _2140_ _2141_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3884_ Tile_X0Y1_N2END[2] Tile_X0Y1_E6END[1] Tile_X0Y1_N4END[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q
+ Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2904_ _1153_ _1210_ _1211_ _1215_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5623_ Tile_X0Y0_E2MID[5] net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2835_ _0882_ _1121_ _1148_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5554_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2766_ _1079_ _1080_ _1081_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4505_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q
+ _0401_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5485_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2697_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q _1014_ _1015_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4436_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1
+ _0335_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4367_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q _0048_ _0049_
+ _0268_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3318_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q _1578_ _1611_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4298_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q _0202_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_69_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3249_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[9\]
+ _1546_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2620_ _0825_ _0926_ _0941_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_124_Right_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput106 net106 Tile_X0Y0_N2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2551_ _0114_ _0875_ _0876_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
Xoutput139 net139 Tile_X0Y0_NN4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput117 net117 Tile_X0Y0_N2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput128 net128 Tile_X0Y0_N4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5270_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2482_ _0667_ _0670_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q
+ _0621_ _0812_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4221_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q _0125_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4152_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q _0056_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4083_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q
+ _2256_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3103_ Tile_X0Y0_EE4END[3] Tile_X0Y0_WW4END[1] Tile_X0Y0_S4END[0] _0561_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q _1412_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3034_ _1327_ _1338_ _1341_ _1306_ _1344_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_55_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4985_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_23_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3936_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q _2125_ _2127_
+ _2128_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3867_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q
+ _2084_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3798_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q _0674_ _2024_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5606_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2818_ _0552_ _0907_ _1131_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5537_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2749_ _0935_ _0936_ _1064_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_1149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5468_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_6_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5399_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4419_ Tile_X0Y1_NN4END[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q
+ _0319_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_1223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_88_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_389 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3721_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q _1967_ _1966_
+ _1968_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3652_ _1913_ _1914_ _1911_ _1912_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_9_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2603_ _0924_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3583_ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[16\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X
+ _0162_ _1851_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2534_ _0113_ _0854_ _0860_ _0861_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5322_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5253_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2465_ _0790_ _0793_ _0795_ _0116_ _0117_ _0796_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4204_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q _0108_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2396_ _0727_ _0730_ _0731_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q _0732_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5184_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X
+ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[14\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4135_ Tile_X0Y0_S2MID[4] _0039_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_3_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_364 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4066_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q
+ _2240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3017_ _0847_ _1192_ _1193_ _1327_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_106_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4968_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4899_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3919_ Tile_X0Y0_S2MID[1] Tile_X0Y0_S4END[5] Tile_X0Y1_W2END[1] Tile_X0Y1_W6END[1]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q
+ _2115_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_11_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_69_Right_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_25_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_78_Right_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5940_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 net335 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_87_Right_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5871_ Tile_X0Y1_FrameData[16] net257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_91_888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4822_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4753_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3704_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 _0374_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2
+ _0407_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4684_ Tile_X0Y1_E6END[1] Tile_X0Y1_W2END[1] Tile_X0Y0_SS4END[5] Tile_X0Y1_W6END[1]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q
+ _0568_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_31_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3635_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q _1898_ _1899_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_96_Right_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3566_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1834_ _1835_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5305_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2517_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q _0843_ _0844_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3497_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[14\]
+ _1782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2448_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q _0215_ _0780_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5236_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_102_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2379_ _0715_ _0716_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5167_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X
+ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[5\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4118_ Tile_X0Y1_E6END[0] _0022_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5098_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_140_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4049_ Tile_X0Y1_W1END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q
+ _2225_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_1188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_100_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3420_ _1707_ _1708_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3351_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4
+ _1642_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2302_ _0456_ Tile_X0Y1_N4END[5] Tile_X0Y1_N2MID[1] Tile_X0Y0_EE4END[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q _0643_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_97_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3282_ _1571_ _1573_ _1576_ _1577_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5021_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_97_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5923_ Tile_X0Y0_SS4END[8] net318 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5854_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 net240 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4805_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_21_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2997_ _0989_ _1049_ _1052_ _1307_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5785_ Tile_X0Y0_W6END[8] net182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4736_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_119_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4667_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q _0549_ _0550_
+ _0551_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3618_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q _1882_ _1859_
+ _1883_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4598_ _0026_ _0482_ _0485_ _0487_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3549_ _0035_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q
+ _1819_ _1820_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5219_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_28_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2920_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q _1113_ _1230_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q _1231_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2851_ Tile_X0Y1_N2END[2] Tile_X0Y1_E2END[2] Tile_X0Y0_S2MID[2] Tile_X0Y1_WW4END[2]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q
+ _1164_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5570_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2782_ _0048_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q _1097_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4521_ _0094_ Tile_X0Y1_W1END[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ _0416_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4452_ _0349_ _0350_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3403_ Tile_X0Y1_E2MID[0] Tile_X0Y1_W2MID[0] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q _1692_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_131_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4383_ Tile_X0Y0_S2MID[4] Tile_X0Y0_S4END[4] Tile_X0Y1_W2END[4] Tile_X0Y1_WW4END[2]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q
+ _0284_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3334_ Tile_X0Y1_NN4END[1] Tile_X0Y1_E2END[5] Tile_X0Y0_S2MID[5] Tile_X0Y1_W2END[5]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q
+ _1626_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3265_ _0412_ _0657_ Tile_X0Y1_W1END[3] Tile_X0Y0_S2MID[7] _0172_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q
+ _1562_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5004_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_127_1121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3196_ _1495_ _1497_ _1494_ _1496_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_138_Right_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5906_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 net301 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5837_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 net223 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5768_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 net163 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_412 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4719_ _0551_ _0598_ _0600_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5699_ Tile_X0Y1_FrameStrobe[13] net85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_134_1169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_364 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_105_Right_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_426 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3050_ _1347_ _1348_ _1360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_48_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3952_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q _0956_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q
+ _2140_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3883_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 _0482_ _0561_ _0468_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2903_ _0551_ _0747_ _1213_ _1214_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5622_ Tile_X0Y0_E2MID[4] net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2834_ _1090_ _1145_ _1147_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5553_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4504_ _0087_ _0399_ _0400_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2765_ _0942_ _0944_ _1077_ _1080_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5484_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2696_ _1013_ _1014_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4435_ _0332_ _0334_ _0330_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4366_ _0262_ _0267_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3317_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q _1604_ _1609_
+ _1610_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4297_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q _0201_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_69_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3248_ _1545_ Tile_X0Y1_DSP_bot.C9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3179_ _1207_ _1375_ _1479_ _1482_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_41_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput107 net107 Tile_X0Y0_N2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2550_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 Tile_X0Y0_E2MID[3] Tile_X0Y0_S2MID[3]
+ Tile_X0Y0_W2MID[3] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q _0875_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_141_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput129 net129 Tile_X0Y0_N4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput118 net118 Tile_X0Y0_N2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2481_ Tile_X0Y0_S2MID[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q _0810_ _0811_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4220_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q _0124_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4151_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q _0055_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4082_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q _2254_ _2255_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3102_ Tile_X0Y0_E2MID[0] Tile_X0Y0_W2MID[0] Tile_X0Y0_S2MID[0] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q
+ _1411_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3033_ _1054_ _1122_ _1342_ _1343_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_66_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4984_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_74_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3935_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q _1188_ _2126_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q _2127_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3866_ _0195_ _2082_ _2083_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5605_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3797_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q _2017_ _2019_
+ _2021_ _2023_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2817_ _0679_ _1053_ _1130_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5536_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2748_ _0997_ _1062_ _1063_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_415 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5467_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2679_ _0995_ _0996_ _0997_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4418_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q Tile_X0Y0_W2END[0]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q _0318_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5398_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_143_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4349_ _0249_ _0251_ _0252_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_6_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Left_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_139_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_443 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_71_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3720_ Tile_X0Y1_N2MID[1] Tile_X0Y1_N4END[5] Tile_X0Y0_E1END[3] Tile_X0Y0_E2END[1]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q
+ _1967_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3651_ Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[2] Tile_X0Y0_SS4END[0] Tile_X0Y0_WW4END[0]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q
+ _1914_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_9_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2602_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q _0923_ _0919_
+ _0924_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_11_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3582_ _1842_ _1845_ _1847_ _1850_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2533_ _0856_ _0859_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q
+ _0860_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5321_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_114_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2464_ _0794_ _0795_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5252_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4203_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q _0107_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2395_ _0033_ _0034_ _0253_ _0038_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q _0731_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5183_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X
+ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[13\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_3_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4134_ Tile_X0Y1_W2MID[1] _0038_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4065_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q _2238_ _2239_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3016_ _0747_ _1239_ _1240_ _1326_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_106_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_446 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4967_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4898_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3918_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q _2113_ _2112_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q _2114_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3849_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q _0346_ _2067_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q _2068_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5519_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_105_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_110_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_69_Left_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5870_ Tile_X0Y1_FrameData[15] net256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4821_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_91_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_78_Left_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4752_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4683_ _0106_ _0566_ _0567_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3703_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 _0346_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1
+ _0321_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3634_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q
+ _1898_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_31_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3565_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[15\]
+ _1835_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_351 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5304_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2516_ _0843_ Tile_X0Y1_DSP_bot.A2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3496_ _1779_ _1780_ _1781_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5235_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2447_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ _0778_ _0779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_87_Left_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2378_ Tile_X0Y1_N2END[0] Tile_X0Y0_S2MID[0] Tile_X0Y1_EE4END[1] Tile_X0Y1_W2END[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q
+ _0715_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5166_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X
+ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[4\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5097_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_56_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4117_ Tile_X0Y1_E1END[0] _0021_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4048_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q _0488_ _2223_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q _2224_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_17_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_96_Left_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_137_1189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_449 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput290 net290 Tile_X0Y1_S2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3350_ _1639_ _1640_ _1641_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2301_ _0101_ _0635_ _0641_ _0642_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3281_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q _1574_ _0176_
+ _1577_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5020_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_119_Right_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5922_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 net308 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5853_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 net239 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4804_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5784_ Tile_X0Y0_W6END[7] net181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_44_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4735_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2996_ _1049_ _1052_ _1122_ _1306_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4666_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[4\]
+ _0550_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4597_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q _0483_ _0484_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q _0486_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3617_ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[17\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X
+ _0162_ _1882_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3548_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4
+ _1819_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3479_ _1762_ _1763_ _1764_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5218_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_88_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5149_ _0015_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[15\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_443 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2850_ _0926_ _1054_ _1156_ _1155_ _1163_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_41_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2781_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q _1094_ _1095_
+ _1096_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4520_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q Tile_X0Y1_W1END[1]
+ _0415_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4451_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ _0348_ _0082_ _0349_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_116_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3402_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q _1685_ _1690_
+ _1691_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4382_ _0054_ _0282_ _0283_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3333_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q _1624_ _1625_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_7_Right_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3264_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q _1560_ _1559_
+ _1561_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5003_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_78_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_127_1122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3195_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q
+ _1497_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_93_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5905_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 net300 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5836_ Tile_X0Y1_E6END[11] net233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2979_ _0926_ _1238_ _1241_ _1289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5767_ Tile_X0Y0_W2END[4] net162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5698_ Tile_X0Y1_FrameStrobe[12] net84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4718_ _0598_ _0599_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4649_ _0091_ _0534_ _0535_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_15_Left_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_49_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_24_Left_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_17_316 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_33_Left_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_141_449 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_42_Left_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3951_ _2139_ _2138_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q
+ Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2902_ _0719_ _0720_ _0847_ _1213_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3882_ _2090_ _2097_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5621_ Tile_X0Y0_E2MID[3] net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_51_Left_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2833_ _1090_ _1145_ _1146_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5552_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2764_ _1071_ _1078_ _1079_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4503_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q
+ _0399_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5483_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2695_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q
+ _1013_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_104_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4434_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q _0333_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q
+ _0334_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4365_ _0264_ _0266_ _0267_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3316_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q _1608_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q
+ _1609_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4296_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q _0200_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_69_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3247_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q _1541_ _1544_
+ _1545_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3178_ _1376_ _1479_ _1480_ _1481_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_26_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5819_ Tile_X0Y1_E2MID[0] net214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_9_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput119 net119 Tile_X0Y0_N2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput108 net108 Tile_X0Y0_N2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_113_1029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2480_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q _0809_ _0810_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4150_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q _0054_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput90 net90 Tile_X0Y0_FrameStrobe_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3101_ Tile_X0Y1_NN4END[6] Tile_X0Y0_E2END[1] Tile_X0Y0_S2END[1] Tile_X0Y0_W2END[1]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q
+ _1410_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4081_ _0203_ _1629_ _2253_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q
+ _2254_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3032_ _1327_ _1338_ _1341_ _1342_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_66_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4983_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3934_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q _1647_ _2126_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3865_ _0915_ _1429_ _0875_ _0346_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q _2082_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_14_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5604_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2816_ _1126_ _1127_ _1129_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3796_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q _2022_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q
+ _2023_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5535_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2747_ _0998_ _1061_ _1062_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5466_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2678_ _0853_ _0908_ _0996_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4417_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q _0222_ _0311_
+ _0314_ _0075_ _0317_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5397_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4348_ _0036_ _0250_ _0037_ _0251_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_6_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4279_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[3\] _0183_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_107_Left_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_399 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_116_Left_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_45_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3650_ _0255_ Tile_X0Y1_N2MID[0] Tile_X0Y0_E1END[0] Tile_X0Y0_E2END[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q _1913_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2601_ _0921_ _0920_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q
+ _0923_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3581_ _0128_ _1848_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q
+ _1850_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2532_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q _0858_ _0859_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5320_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5251_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_130_1140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2463_ Tile_X0Y1_N2MID[4] Tile_X0Y0_E2END[4] Tile_X0Y0_SS4END[2] Tile_X0Y0_W2END[4]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q
+ _0794_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4202_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q _0106_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2394_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q _0729_ _0730_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5182_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X
+ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[12\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4133_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q _0037_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4064_ Tile_X0Y1_E1END[3] Tile_X0Y1_W1END[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q _2238_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3015_ _0846_ _1239_ _1240_ _1325_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_336 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4966_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3917_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q
+ _2113_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4897_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_137_316 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3848_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q _0795_ _2067_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3779_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q _2008_ _2009_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5518_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_105_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5449_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_120_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_439 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_351 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4820_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_103_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4751_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3702_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 _0630_ _1956_ _0653_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4682_ Tile_X0Y1_N2END[1] Tile_X0Y1_N4END[1] Tile_X0Y1_E1END[3] Tile_X0Y1_E2END[1]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q
+ _0566_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3633_ _1896_ _1897_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3564_ _1808_ _1811_ _1831_ _1834_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2515_ _0841_ _0842_ _0843_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5303_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3495_ _1418_ _1778_ _1400_ _1780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5234_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2446_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q _0209_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q
+ _0778_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5165_ Tile_X0Y1_DSP_bot.B3 clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[3\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2377_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q _0711_ _0713_
+ _0714_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4116_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q _0020_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5096_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_110_293 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4047_ Tile_X0Y1_N1END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q
+ _2223_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4949_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput280 net280 Tile_X0Y1_FrameData_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput291 net291 Tile_X0Y1_S2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2300_ _0637_ _0640_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q
+ _0641_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3280_ _0175_ _1575_ _1576_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5921_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 net307 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5852_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 net238 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4803_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_44_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5783_ Tile_X0Y0_W6END[6] net180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4734_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2995_ _0748_ _1194_ _1305_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4665_ _0549_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4596_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q _0484_ _0485_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3616_ _1874_ _1881_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3547_ _0126_ _1816_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q
+ _1818_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3478_ _1366_ _1368_ _1639_ _1763_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5217_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_76_409 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2429_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q _0759_ _0762_
+ _0763_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5148_ _0014_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[14\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5079_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_56_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2780_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q _0436_ _1095_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4450_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q _0347_ _0348_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_116_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4381_ Tile_X0Y1_N2END[4] Tile_X0Y1_E2END[4] Tile_X0Y1_E1END[2] Tile_X0Y1_E6END[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q
+ _0282_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3401_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q _1689_ _1690_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3332_ _1623_ _1624_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3263_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q
+ _1560_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5002_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3194_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q
+ _1496_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_127_1123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5904_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 net299 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5835_ Tile_X0Y1_E6END[10] net232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2978_ _1285_ _1286_ _1287_ _1288_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5766_ Tile_X0Y0_W2END[3] net161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5697_ Tile_X0Y1_FrameStrobe[11] net83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4717_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q _0596_ _0597_
+ _0598_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4648_ Tile_X0Y0_E6END[1] Tile_X0Y0_S2END[3] Tile_X0Y0_W2END[3] Tile_X0Y0_WW4END[1]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q
+ _0534_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_1_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4579_ _0465_ _0467_ _0026_ _0462_ _0469_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_32_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3950_ Tile_X0Y1_N1END[1] Tile_X0Y1_W1END[1] Tile_X0Y1_E1END[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q
+ _2139_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2901_ _0721_ _0747_ _1211_ _1212_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3881_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q _2096_ _2095_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q _2097_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5620_ Tile_X0Y0_E2MID[2] net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2832_ _1143_ _1144_ _1145_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5551_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_77_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2763_ _1077_ _1078_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4502_ _0393_ _0398_ _0384_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5482_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2694_ _1011_ _1012_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4433_ Tile_X0Y0_E6END[0] Tile_X0Y0_W2END[2] Tile_X0Y0_S2END[2] Tile_X0Y0_WW4END[3]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q
+ _0333_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_133_1160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4364_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q _0265_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q
+ _0266_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3315_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q _1605_ _1607_
+ _1608_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4295_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q _0199_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3246_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q _1543_ _1544_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3177_ _1257_ _1374_ _1207_ _1480_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5818_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 net213 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5749_ Tile_X0Y1_NN4END[15] net150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_60_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_386 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput109 net109 Tile_X0Y0_N2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput1 net1 Tile_X0Y0_E1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput80 net80 Tile_X0Y0_FrameData_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput91 net91 Tile_X0Y0_FrameStrobe_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3100_ _1403_ _1405_ _1407_ _1409_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4080_ _0203_ _1707_ _2253_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3031_ _0989_ _1192_ _1193_ _1238_ _1241_ _0847_ _1341_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai33_1
XTAP_TAPCELL_ROW_66_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4982_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3933_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ _2124_ _2125_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3864_ _0195_ _2080_ _2081_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5603_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2815_ _1126_ _1127_ _1128_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3795_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q
+ _2022_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5534_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2746_ _0722_ _1055_ _1057_ _1061_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_117_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5465_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2677_ _0851_ _0990_ _0994_ _0748_ _0995_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4416_ _0315_ _0316_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5396_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4347_ Tile_X0Y0_S4END[2] Tile_X0Y0_SS4END[2] Tile_X0Y0_W2END[2] Tile_X0Y0_W6END[0]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q
+ _0250_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_6_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4278_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q _0182_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3229_ _0166_ _1528_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q
+ _1529_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3580_ _1848_ _1849_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2600_ _0921_ _0922_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2531_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q _0211_ _0857_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q _0858_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5250_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_130_1141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4201_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q _0105_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2462_ _0116_ _0792_ _0793_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2393_ _0133_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q
+ _0728_ _0729_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_68_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5181_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X
+ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[11\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4132_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q _0036_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4063_ _2237_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_3_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3014_ _1282_ _1307_ _1324_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4965_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_106_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3916_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q _2111_ _2112_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4896_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3847_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ _2065_ _2066_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3778_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q _0815_ _2007_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q _2008_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2729_ Tile_X0Y1_N2END[4] Tile_X0Y1_E2END[4] Tile_X0Y0_SS4END[6] Tile_X0Y1_W2END[4]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q
+ _1045_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5517_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_105_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5448_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5379_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_59_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_29_Right_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_38_Right_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_136_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_47_Right_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4750_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_56_Right_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3701_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q _1951_ _1953_
+ _1955_ _1956_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4681_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q _0564_ _0107_
+ _0565_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3632_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q
+ _1896_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_119_1069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5302_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3563_ _1811_ _1831_ _1833_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2514_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q _0839_ _0837_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q _0842_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3494_ _1400_ _1418_ _1778_ _1779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_65_Right_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5233_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2445_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q
+ _0777_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5164_ Tile_X0Y1_DSP_bot.B2 clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[2\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2376_ Tile_X0Y1_N4END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q
+ _0712_ _0713_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4115_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1936_ _0019_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5095_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4046_ _0201_ _2221_ _2222_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_74_Right_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_135_Left_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4948_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_90_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4879_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_30_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_83_Right_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput270 net270 Tile_X0Y1_FrameData_O[28] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput292 net292 Tile_X0Y1_S2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput281 net281 Tile_X0Y1_FrameData_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_92_Right_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_133_Right_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5920_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 net306 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5851_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 net237 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4802_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_44_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2994_ _1277_ _1302_ _1303_ _1304_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5782_ Tile_X0Y0_W6END[5] net179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_100_Right_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4733_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_9_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4664_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q _0540_ _0545_
+ _0548_ _0549_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4595_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ _0484_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3615_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q _0321_ _1880_
+ _1881_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_136_1180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3546_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q _0346_ _1817_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5216_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3477_ _1365_ _1656_ _1657_ _1760_ _1761_ _1762_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2428_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q _0761_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q
+ _0762_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5147_ _0013_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[13\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2359_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q _0696_ _0697_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5078_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4029_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ _2207_ _2208_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_425 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_375 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_432 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4380_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q _0280_ _0055_
+ _0281_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3400_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q _1686_ _1688_
+ _1689_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3331_ Tile_X0Y1_E6END[1] Tile_X0Y0_S4END[5] Tile_X0Y1_WW4END[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q
+ _1623_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3262_ _1555_ _1556_ _1558_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q _1559_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_85_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5001_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3193_ Tile_X0Y1_N1END[2] Tile_X0Y1_E1END[2] Tile_X0Y1_N2END[6] Tile_X0Y1_E2END[6]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q
+ _1495_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_127_1124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5903_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 net298 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5834_ Tile_X0Y1_E6END[9] net231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2977_ _0846_ _1050_ _1051_ _1287_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5765_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 net160 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5696_ Tile_X0Y1_FrameStrobe[10] net82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4716_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[7\]
+ _0597_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_437 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4647_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q _0532_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q
+ _0533_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4578_ _0464_ _0466_ _0463_ _0468_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3529_ _1772_ _1773_ _1803_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_130_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2900_ _0552_ _0847_ _1211_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_122_1087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3880_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q
+ _2096_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2831_ _1066_ _1067_ _1144_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5550_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2762_ _1074_ _1075_ _1077_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5481_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4501_ _0397_ _0398_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2693_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q _1010_ _1011_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4432_ _0081_ _0331_ _0332_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_133_1161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4363_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ _0265_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4294_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q _0198_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3314_ _0025_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q
+ _1606_ _1607_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_58_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3245_ _1542_ _1543_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_69_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3176_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q _0164_ _1477_
+ _1478_ _1479_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_446 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5817_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 net212 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5748_ Tile_X0Y1_NN4END[14] net149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5679_ Tile_X0Y0_FrameData[25] net66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_9_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput2 net2 Tile_X0Y0_E1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput70 net70 Tile_X0Y0_FrameData_O[29] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput81 net81 Tile_X0Y0_FrameStrobe_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput92 net92 Tile_X0Y0_FrameStrobe_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3030_ _1327_ _1338_ _1340_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_66_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4981_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_63_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3932_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q _0956_ _2124_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3863_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q
+ _2080_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_31_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5602_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2814_ _0992_ _0993_ _1127_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3794_ _0194_ _2020_ _2021_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5533_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_117_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2745_ _0723_ _1059_ _1060_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5464_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2676_ _0882_ _0992_ _0994_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5395_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4415_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q _0222_ _0311_
+ _0314_ _0315_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4346_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q _0248_ _0249_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_6_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4277_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q _0181_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_357 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3228_ Tile_X0Y1_N1END[2] Tile_X0Y1_E1END[2] Tile_X0Y1_N2END[6] Tile_X0Y1_E2END[6]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q
+ _1528_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_86_379 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3159_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q _0421_ _1463_
+ _1464_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_63_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2530_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ _0857_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2461_ _0100_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q
+ _0791_ _0792_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_39_Left_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4200_ Tile_X0Y0_W2MID[4] _0104_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_130_1142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2392_ Tile_X0Y1_N2MID[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q
+ _0728_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5180_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X
+ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[10\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4131_ Tile_X0Y0_W2END[2] _0035_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4062_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q _2231_ _2236_
+ _2237_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3013_ _1282_ _1307_ _1323_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_48_Left_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4964_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3915_ _2110_ _2111_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4895_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3846_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q _1430_ _2065_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3777_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q _1460_ _2007_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5516_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2728_ Tile_X0Y1_NN4END[1] Tile_X0Y1_EE4END[1] Tile_X0Y0_S4END[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q
+ _1044_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_105_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5447_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2659_ Tile_X0Y1_NN4END[0] Tile_X0Y0_S2MID[2] Tile_X0Y1_E2END[2] Tile_X0Y1_W2END[2]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q
+ _0978_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5378_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4329_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q
+ _0232_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_101_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_114_Right_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_281 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ _0067_ _1954_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q
+ _1955_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4680_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q
+ _0564_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_41_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3631_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q _1894_ _1893_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q _1895_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3562_ _1811_ _1831_ _1832_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_142_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2513_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q _0827_ _0840_
+ _0841_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5301_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3493_ _1416_ _1417_ _1774_ _1775_ _1427_ _1778_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_142_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5232_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2444_ _0775_ _0776_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2375_ _0140_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q
+ _0712_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5163_ Tile_X0Y1_DSP_bot.B1 clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4114_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1940_ _0018_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5094_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4045_ _0201_ _2220_ _2222_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_56_Left_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4947_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_90_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4878_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3829_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q _1420_ _2050_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q _2051_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_30_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput260 net260 Tile_X0Y1_FrameData_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput271 net271 Tile_X0Y1_FrameData_O[29] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput282 net282 Tile_X0Y1_S1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput293 net293 Tile_X0Y1_S2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5850_ Tile_X0Y1_EE4END[15] net236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4801_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_44_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2993_ _1275_ _1276_ _1303_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5781_ Tile_X0Y0_W6END[4] net178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4732_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4663_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q _0547_ _0548_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3614_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q _1879_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q
+ _1880_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4594_ _0482_ _0483_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_136_1181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3545_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 Tile_X0Y0_W2MID[2] Tile_X0Y0_S2MID[2]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q _1816_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3476_ _1362_ _1364_ _1656_ _1761_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5215_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2427_ _0760_ _0761_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5146_ _0012_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[12\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2358_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q
+ _0696_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2289_ _0623_ _0626_ _0628_ _0630_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5077_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4028_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q _1707_ _2207_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5979_ Tile_X0Y1_WW4END[12] net380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3330_ _1620_ _1621_ _1622_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5000_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3261_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ _1557_ _1558_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3192_ _0489_ _0351_ Tile_X0Y0_S2MID[6] Tile_X0Y1_W1END[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q _1494_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_127_1125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5902_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 net297 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5833_ Tile_X0Y1_E6END[8] net230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2976_ _0719_ _0720_ _0989_ _1283_ _1286_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_5764_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 net159 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5695_ Tile_X0Y1_FrameStrobe[9] net100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4715_ _0596_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4646_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q
+ _0532_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4577_ _0466_ _0467_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3528_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1801_ _1802_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3459_ _1744_ _0272_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q
+ _1745_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5129_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_29_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_400 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Left_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_122_1088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_322 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2830_ _1142_ _1143_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2761_ _0598_ _0882_ _1074_ _1076_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5480_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2692_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q _1009_ _1010_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4500_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q _0396_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q
+ _0397_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_1 Tile_X0Y0_E6END[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4431_ _0255_ Tile_X0Y1_N2MID[2] Tile_X0Y1_N4END[6] Tile_X0Y0_E2END[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q _0331_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_20_Left_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_133_1162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4362_ _0047_ _0263_ _0264_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4293_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q _0197_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3313_ Tile_X0Y1_W2END[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q
+ _1606_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3244_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q
+ _1542_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_100_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3175_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[10\]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q _1478_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5816_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 net211 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5747_ Tile_X0Y1_NN4END[13] net148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2959_ _0679_ _1242_ _1269_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5678_ Tile_X0Y0_FrameData[24] net65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4629_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q _0516_ _0517_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_128_Right_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput3 net3 Tile_X0Y0_E1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput60 net60 Tile_X0Y0_FrameData_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_441 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput93 net93 Tile_X0Y0_FrameStrobe_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput82 net82 Tile_X0Y0_FrameStrobe_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput71 net71 Tile_X0Y0_FrameData_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_124_1106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4980_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_51_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3931_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 _0455_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2
+ _0436_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3862_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q _2078_ _2079_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2813_ _0990_ _1123_ _1124_ _1125_ _1126_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_82_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5601_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3793_ _0915_ _1429_ _0875_ _0346_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q _2020_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5532_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_31_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2744_ _0721_ _0927_ _1059_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5463_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2675_ _0747_ _0882_ _0993_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5394_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4414_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q _0313_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q
+ _0314_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4345_ Tile_X0Y1_NN4END[6] Tile_X0Y0_E1END[0] Tile_X0Y0_EE4END[2] Tile_X0Y0_E6END[0]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q
+ _0248_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_98_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4276_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q _0180_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3227_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q _1526_ _1527_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3158_ Tile_X0Y0_E2MID[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q _1463_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_142_1217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3089_ _0529_ _1398_ _1399_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2460_ Tile_X0Y1_NN4END[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q
+ _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_130_1143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2391_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0
+ _0726_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q _0727_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4130_ Tile_X0Y1_E2MID[1] _0034_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_79_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4061_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q _2235_ _2233_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q _2236_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3012_ _1320_ _1321_ _1322_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_19_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4963_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_51_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3914_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q
+ _2110_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4894_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3845_ _2064_ _2063_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3776_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q _0673_ _2005_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q _2006_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5515_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2727_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q _1041_ _1043_
+ _1037_ _1039_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5446_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2658_ _0971_ _0973_ _0975_ _0977_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2589_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3
+ _0911_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5377_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4328_ Tile_X0Y1_N4END[2] Tile_X0Y1_E2END[2] Tile_X0Y1_W2END[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q
+ _0231_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4259_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q _0163_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_2_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3630_ Tile_X0Y0_S1END[0] Tile_X0Y0_S2END[0] Tile_X0Y0_S1END[2] Tile_X0Y0_W1END[0]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q
+ _1894_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3561_ _1830_ _1831_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2512_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q _0455_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q
+ _0840_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5300_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_5_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3492_ _1427_ _1776_ _1777_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5231_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2443_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q _0773_ _0774_
+ _0775_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2374_ Tile_X0Y1_W6END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q _0710_ _0711_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5162_ Tile_X0Y1_DSP_bot.B0 clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[0\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_99_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5093_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4113_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1885_ _0017_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4044_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q _2217_ _2219_
+ _2221_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_3_Left_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_39_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4946_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_90_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4877_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_22_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3828_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ _2050_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3759_ _1991_ _1990_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_30_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput261 net261 Tile_X0Y1_FrameData_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5429_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput250 net250 Tile_X0Y1_FrameData_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput294 net294 Tile_X0Y1_S2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput283 net283 Tile_X0Y1_S1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput272 net272 Tile_X0Y1_FrameData_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_44_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2992_ _1300_ _1301_ _1299_ _1302_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5780_ Tile_X0Y0_W6END[3] net177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4731_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4662_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q _0546_ _0547_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3613_ _1876_ _1878_ _1879_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4593_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 Tile_X0Y0_S2MID[1] Tile_X0Y0_E2MID[1]
+ Tile_X0Y0_W2MID[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q _0482_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_136_1182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3544_ _1814_ _1815_ _1812_ _1813_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3475_ _1758_ _1759_ _1683_ _1760_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_388 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5214_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2426_ Tile_X0Y0_S2END[3] Tile_X0Y0_W2END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_W6END[1]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q
+ _0760_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2357_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q Tile_X0Y1_W2MID[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q _0695_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5145_ _0011_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[11\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2288_ _0628_ _0629_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5076_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4027_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q _1629_ _2205_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q _2206_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5978_ Tile_X0Y1_WW4END[11] net379 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4929_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_100_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_449 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_109_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_75_Left_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_84_Left_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3260_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q _0212_ _1557_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3191_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q _1486_ _1491_
+ _1493_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5901_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 net296 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_93_Left_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5832_ Tile_X0Y1_E6END[7] net229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5763_ Tile_X0Y0_W2END[0] net158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2975_ _0719_ _0720_ _0989_ _1283_ _1285_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4714_ _0574_ _0595_ _0596_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5694_ Tile_X0Y1_FrameStrobe[8] net99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4645_ _0091_ _0530_ _0531_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4576_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q Tile_X0Y0_W2END[7]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q _0466_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_450 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_408 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3527_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[10\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ _1802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3458_ Tile_X0Y1_N2MID[6] Tile_X0Y1_W2MID[6] Tile_X0Y1_E2MID[6] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q
+ _1744_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_130_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2409_ _0742_ _0741_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q
+ _0744_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3389_ _1678_ Tile_X0Y1_DSP_bot.C4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5128_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_72_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5059_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_55_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_109_Right_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_96_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_1089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2760_ _0598_ _0882_ _1075_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2691_ Tile_X0Y1_N1END[1] Tile_X0Y1_N2END[5] Tile_X0Y1_E1END[1] Tile_X0Y1_E2END[5]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q
+ _1009_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_2 Tile_X0Y0_E6END[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4430_ _0081_ _0323_ _0329_ _0330_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_133_1163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4361_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q
+ _0263_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_98_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4292_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q _0196_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3312_ Tile_X0Y1_N2END[1] Tile_X0Y1_EE4END[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q
+ _1605_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3243_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 _1521_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q _1541_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_39_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3174_ _0162_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X
+ _1477_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5815_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 net210 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_52_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5746_ Tile_X0Y1_NN4END[12] net147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2958_ _1258_ _1260_ _1261_ _1268_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5677_ Tile_X0Y0_FrameData[23] net64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4628_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q _0513_ _0515_
+ _0516_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2889_ _1199_ _1200_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4559_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y0_E1END[2] Tile_X0Y1_N2MID[6]
+ Tile_X0Y0_E2END[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q _0451_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_103_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput4 net4 Tile_X0Y0_E1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput61 net61 Tile_X0Y0_FrameData_O[20] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput50 net50 Tile_X0Y0_FrameData_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput72 net72 Tile_X0Y0_FrameData_O[30] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput94 net94 Tile_X0Y0_FrameStrobe_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput83 net83 Tile_X0Y0_FrameStrobe_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3930_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1
+ _1651_ _1604_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3861_ Tile_X0Y0_E1END[3] Tile_X0Y0_W1END[3] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q _2078_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_31_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3792_ _0194_ _2018_ _2019_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5600_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2812_ _0846_ _0882_ _1125_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5531_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2743_ _0552_ _0926_ _0722_ _1058_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5462_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2674_ _0848_ _0991_ _0992_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5393_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4413_ _0312_ _0313_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4344_ _0037_ _0244_ _0246_ _0247_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_140_283 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4275_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q _0179_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3226_ _0351_ Tile_X0Y0_S2MID[6] Tile_X0Y1_W1END[0] Tile_X0Y1_W1END[2] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q _1526_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3157_ _0121_ _1459_ _1461_ _1462_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_142_1218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3088_ _1389_ _1397_ _1398_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_42_429 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5729_ Tile_X0Y1_N4END[11] net130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_112_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_130_1144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2390_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q _0241_ _0726_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_79_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4060_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ _2234_ _2235_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3011_ _1300_ _1301_ _1321_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_19_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4962_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4893_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3913_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 _0254_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3
+ _0231_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3844_ _0456_ Tile_X0Y0_W1END[3] Tile_X0Y0_S1END[3] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q
+ _2064_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3775_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ _2005_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5514_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2726_ _0151_ _1042_ _1043_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2657_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q _0976_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q
+ _0977_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5445_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_120_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5376_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2588_ _0852_ _0909_ _0910_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4327_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q _0228_ _0230_
+ _0224_ _0226_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4258_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q _0162_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3209_ _0169_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 _1510_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_85_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4189_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q _0093_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_105_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_399 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_16_Right_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_16_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_25_Right_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3560_ _0163_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[15\] _1829_ _1830_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2511_ _0838_ _0839_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5230_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3491_ _1774_ _1775_ _1776_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2442_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[7\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q
+ _0774_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2373_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q _0445_ _0710_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5161_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X
+ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[7\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_99_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5092_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_68_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4112_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1856_ _0016_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4043_ Tile_X0Y1_N1END[3] Tile_X0Y1_W1END[3] _0412_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q
+ _2220_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_34_Right_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_39_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_370 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4945_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_90_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4876_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_22_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_421 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_43_Right_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3827_ _2049_ _2048_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3758_ _0255_ Tile_X0Y0_W1END[0] Tile_X0Y0_E1END[0] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q
+ _1991_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_104_Left_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_30_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2709_ _1019_ _1021_ _1024_ _1026_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3689_ _1768_ _1944_ _1945_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput240 net240 Tile_X0Y1_EE4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput251 net251 Tile_X0Y1_FrameData_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5428_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput262 net262 Tile_X0Y1_FrameData_O[20] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput284 net284 Tile_X0Y1_S1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput295 net295 Tile_X0Y1_S2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5359_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput273 net273 Tile_X0Y1_FrameData_O[30] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_307 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_52_Right_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_59_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_113_Left_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Right_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_122_Left_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_70_Right_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_131_Left_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_65_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2991_ _1297_ _1298_ _1301_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_140_Left_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_44_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_398 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4730_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4661_ Tile_X0Y0_E2MID[6] Tile_X0Y0_W2MID[6] Tile_X0Y0_S2MID[6] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q
+ _0546_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3612_ _0066_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q
+ _1877_ _1878_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4592_ _0480_ _0481_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_136_1183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3543_ Tile_X0Y0_S1END[1] Tile_X0Y0_S2END[7] Tile_X0Y0_S1END[3] Tile_X0Y0_W1END[3]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q
+ _1815_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3474_ _1681_ _1682_ _1759_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5213_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2425_ _0306_ Tile_X0Y0_E2END[3] Tile_X0Y1_N2MID[3] Tile_X0Y0_E6END[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q _0759_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5144_ _0010_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[10\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2356_ _0686_ _0689_ _0692_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q
+ _0137_ _0694_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_56_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2287_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q Tile_X0Y0_S2MID[7]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q _0627_ _0628_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5075_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4026_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q _0743_ _2205_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5977_ Tile_X0Y1_WW4END[10] net378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4928_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4859_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_133_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3190_ _0165_ _1492_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q
+ _1493_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5900_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 net295 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_332 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5831_ Tile_X0Y1_E6END[6] net228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2974_ _1259_ _1282_ _1284_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5762_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 net157 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4713_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q _0593_ _0592_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q _0595_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5693_ Tile_X0Y1_FrameStrobe[7] net98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4644_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q
+ _0530_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4575_ _0393_ _0398_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q
+ _0384_ _0465_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3526_ _1482_ _1771_ _1801_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3457_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q _1742_ _1740_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q _1743_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2408_ _0742_ _0743_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3388_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q _1662_ _1667_
+ _1672_ _1677_ _1678_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_111_370 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2339_ _0677_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5127_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_2_Right_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_57_446 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5058_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4009_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q _2188_ _2190_
+ _2191_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_115_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2690_ _0999_ _1003_ _1004_ _1005_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q
+ _1008_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_77_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_3 Tile_X0Y0_E6END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4360_ _0257_ _0259_ _0261_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q
+ _0262_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_133_1164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3311_ _1603_ _1604_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4291_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q _0195_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3242_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q _1533_ _1538_
+ _1540_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_307 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3173_ _1475_ _1476_ _1462_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5814_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 net209 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5745_ Tile_X0Y1_NN4END[11] net146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2957_ _0926_ _1194_ _1267_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5676_ Tile_X0Y0_FrameData[22] net63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2888_ _1197_ _1198_ _1162_ _1199_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4627_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q _0211_ _0514_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q _0515_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4558_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q _0447_ _0449_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q _0450_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3509_ _1755_ _1756_ _1790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4489_ _0274_ _0276_ _0304_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ _0386_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_89_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_142_Right_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_408 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_324 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_390 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput5 net5 Tile_X0Y0_E2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput51 net51 Tile_X0Y0_FrameData_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_281 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput40 net40 Tile_X0Y0_EE4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput73 net73 Tile_X0Y0_FrameData_O[31] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput84 net84 Tile_X0Y0_FrameStrobe_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput62 net62 Tile_X0Y0_FrameData_O[21] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_443 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput95 net95 Tile_X0Y0_FrameStrobe_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3860_ _2077_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3791_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q
+ _2018_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2811_ _0990_ _1123_ _1124_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_14_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5530_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_31_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2742_ _0552_ _0926_ _1057_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5461_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_117_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2673_ _0775_ _0988_ _0991_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4412_ Tile_X0Y0_S1END[1] Tile_X0Y0_S2END[5] Tile_X0Y0_S1END[3] Tile_X0Y0_W1END[1]
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ _0312_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5392_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4343_ _0036_ _0245_ _0246_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_99_Right_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4274_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q _0178_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3225_ _0166_ _1522_ _0167_ _1525_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3156_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q _1458_ _1461_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_142_1219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3087_ _1395_ _1396_ _1397_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5728_ Tile_X0Y1_N4END[10] net129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3989_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q
+ _2173_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5659_ Tile_X0Y0_FrameData[5] net76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_1145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3010_ _1318_ _1319_ _1317_ _1320_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_19_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4961_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4892_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3912_ Tile_X0Y0_S2MID[1] Tile_X0Y0_S4END[4] Tile_X0Y1_W6END[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_17_Left_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3843_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 _0674_ _0815_ _1419_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q
+ _2063_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xclkbuf_0_Tile_X0Y1_UserCLK Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3774_ _2004_ _2003_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5513_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2725_ Tile_X0Y0_S2MID[3] Tile_X0Y1_W2END[3] Tile_X0Y0_S4END[7] Tile_X0Y1_W6END[1]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q
+ _1042_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2656_ Tile_X0Y1_E6END[0] Tile_X0Y0_S2MID[4] Tile_X0Y1_W2END[4] Tile_X0Y1_W6END[0]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q
+ _0976_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5444_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_5375_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2587_ _0853_ _0908_ _0909_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_26_Left_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4326_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q _0229_ _0230_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4257_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[12\] _0161_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_2_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3208_ _0169_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 _1508_ _1509_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4188_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q _0092_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3139_ Tile_X0Y1_NN4END[6] Tile_X0Y0_S4END[2] Tile_X0Y0_E2END[2] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q
+ _1445_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_85_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2510_ Tile_X0Y1_N2END[4] Tile_X0Y0_S2MID[4] Tile_X0Y1_EE4END[0] Tile_X0Y1_W2END[4]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q
+ _0838_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3490_ _1425_ _1426_ _1775_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_5_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2441_ _0773_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2372_ _0706_ _0708_ _0709_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5160_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X
+ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[6\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5091_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4111_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr _1834_ _0015_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4042_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q _0827_ _2218_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q _2219_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_82_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4944_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_90_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4875_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_102_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3826_ _0255_ Tile_X0Y0_W1END[0] Tile_X0Y0_E1END[0] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q
+ _2049_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3757_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q _1989_ _1987_
+ _1990_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_332 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2708_ _1024_ _1025_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3688_ _1622_ _1766_ _1767_ _1944_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xoutput230 net230 Tile_X0Y1_E6BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput241 net241 Tile_X0Y1_EE4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2639_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q _0959_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q
+ _0960_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5427_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput252 net252 Tile_X0Y1_FrameData_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput285 net285 Tile_X0Y1_S1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5358_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput263 net263 Tile_X0Y1_FrameData_O[21] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput274 net274 Tile_X0Y1_FrameData_O[31] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput296 net296 Tile_X0Y1_S2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4309_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 _0213_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5289_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_101_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_118_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2990_ _1290_ _1295_ _1300_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_44_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4660_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q _0542_ _0544_
+ _0545_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3611_ Tile_X0Y0_W2END[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q
+ _1877_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4591_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q _0479_ _0480_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_136_1184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3542_ _0456_ Tile_X0Y0_E1END[3] Tile_X0Y1_N2MID[7] Tile_X0Y0_E2END[7] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q _1814_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_115_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3473_ _1699_ _1757_ _1758_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5212_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2424_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q _0752_ _0757_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q _0758_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2355_ _0686_ _0689_ _0692_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q
+ _0693_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5143_ _0009_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[9\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_433 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5074_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2286_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q _0064_ _0627_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4025_ _2204_ _2203_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5976_ Tile_X0Y1_WW4END[9] net377 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4927_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_100_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4858_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_20_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3809_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q _2031_ _2034_
+ _2035_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4789_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_87_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5830_ Tile_X0Y1_E6END[5] net227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2973_ _0552_ _1122_ _1283_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5761_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 net156 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4712_ _0593_ _0594_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5692_ Tile_X0Y1_FrameStrobe[6] net97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_408 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4643_ _0163_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[14\] _0528_ _0529_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4574_ _0394_ _0397_ _0031_ _0385_ _0464_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_143_441 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3525_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1
+ _1651_ _1604_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_123_Right_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_115_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3456_ _1741_ _1742_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2407_ Tile_X0Y1_N2END[0] Tile_X0Y0_S2MID[0] Tile_X0Y1_E2END[0] Tile_X0Y1_WW4END[3]
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q
+ _0742_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3387_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q _1676_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q
+ _1677_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2338_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q _0608_ _0676_
+ _0677_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5126_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2269_ _0069_ _0610_ _0611_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5057_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_4008_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q _1188_ _2189_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q _2190_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_25_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_9_Left_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5959_ Tile_X0Y1_W6END[2] net354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_414 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_377 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_4 Tile_X0Y0_EE4END[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_3310_ _1600_ _1602_ _1603_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4290_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q _0194_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3241_ _0168_ _1539_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q
+ _1540_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3172_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q _0630_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q
+ _1476_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_13_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5813_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 net208 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5744_ Tile_X0Y1_NN4END[10] net145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2956_ _1209_ _1215_ _1263_ _1266_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5675_ Tile_X0Y0_FrameData[21] net62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_60_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2887_ _1151_ _1159_ _1161_ _1198_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4626_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ _0514_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4557_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q _0448_ _0449_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3508_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q _1788_ _1789_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4488_ _0384_ _0385_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3439_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q _1725_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q
+ _1726_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5109_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_68_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput6 net6 Tile_X0Y0_E2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput52 net52 Tile_X0Y0_FrameData_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput30 net30 Tile_X0Y0_E6BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput41 net41 Tile_X0Y0_EE4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput74 net74 Tile_X0Y0_FrameData_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput63 net63 Tile_X0Y0_FrameData_O[22] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput85 net85 Tile_X0Y0_FrameStrobe_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_8_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput96 net96 Tile_X0Y0_FrameStrobe_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3790_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q _2016_ _2017_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2810_ _0775_ _1121_ _1123_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2741_ _1055_ _1056_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5460_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_8_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2672_ _0822_ _0823_ _0989_ _0990_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4411_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q _0307_ _0308_
+ _0310_ _0311_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5391_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_125_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4342_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q
+ _0245_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_98_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4273_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q _0177_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3224_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q _1523_ _1524_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
.ends

