`default_nettype none

module fabric_wrapper #(
    	parameter FrameBitsPerRow = 32,
	parameter MaxFramesPerCol = 20,
	
	parameter NumColumns = 12,
	parameter NumRows = 18,
	
    parameter FABRIC_NUM_IO_WEST = 32
)(
    input clk_i,
    
    // Configuration
    input  logic [(FrameBitsPerRow*NumRows)-1:0]    FrameData_i,
    input  logic [(MaxFramesPerCol*NumColumns)-1:0] FrameStrobe_i,
    
    // Fabric is configured
    input                                 configured_i,

    // I/Os West
    input  [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_in_i,
    output [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_out_o,
    output [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_oe_o,

    // WARMBOOT
    output        fabric_warmboot_boot_o,
    output  [3:0] fabric_warmboot_slot_o,
    input         fabric_warmboot_reset_i,

    // CPU_IRQ
    output  [3:0] fabric_irq_o,
    
    // CUSTOM_INSTRUCTION
    output logic        fabric_issue_ready_o,
    output logic        fabric_issue_accept_o,
    input  logic        fabric_issue_valid_i,
    input  logic [31:0] fabric_issue_instr_i,
    input  logic [31:0] fabric_issue_op0_i,
    input  logic [31:0] fabric_issue_op1_i,
    input  logic [3 :0] fabric_issue_id_i,
    
    output logic        fabric_result_valid_o,
    output logic [3 :0] fabric_result_id_o,
    output logic [4 :0] fabric_result_rd_o,
    output logic [31:0] fabric_result_o,

    // OBI_PERIPHERAL
    input          fabric_obi_req_i,
    input          fabric_obi_we_i,
    input   [3 :0] fabric_obi_be_i,
    input   [23:0] fabric_obi_addr_i,
    input   [31:0] fabric_obi_wdata_i,
    output         fabric_obi_gnt_o,
    output         fabric_obi_rvalid_o,
    output  [31:0] fabric_obi_rdata_o
);

    // SRAM 0
    logic [31:0] fabric_sram0_a_dout_i;
    logic [9 :0] fabric_sram0_a_addr_o;
    logic [31:0] fabric_sram0_a_bm_o;
    logic [31:0] fabric_sram0_a_din_o;
    logic        fabric_sram0_a_wen_o;
    logic        fabric_sram0_a_men_o;
    logic        fabric_sram0_a_ren_o;
    logic        fabric_sram0_a_clk_o;
    logic        fabric_sram0_a_tie_high_o;
    logic        fabric_sram0_a_tie_low_o;

    // SRAM 1
    logic [31:0] fabric_sram1_a_dout_i;
    logic [9 :0] fabric_sram1_a_addr_o;
    logic [31:0] fabric_sram1_a_bm_o;
    logic [31:0] fabric_sram1_a_din_o;
    logic        fabric_sram1_a_wen_o;
    logic        fabric_sram1_a_men_o;
    logic        fabric_sram1_a_ren_o;
    logic        fabric_sram1_a_clk_o;
    logic        fabric_sram1_a_tie_high_o;
    logic        fabric_sram1_a_tie_low_o;

    // SRAM 2
    logic [31:0] fabric_sram2_a_dout_i;
    logic [9 :0] fabric_sram2_a_addr_o;
    logic [31:0] fabric_sram2_a_bm_o;
    logic [31:0] fabric_sram2_a_din_o;
    logic        fabric_sram2_a_wen_o;
    logic        fabric_sram2_a_men_o;
    logic        fabric_sram2_a_ren_o;
    logic        fabric_sram2_a_clk_o;
    logic        fabric_sram2_a_tie_high_o;
    logic        fabric_sram2_a_tie_low_o;

    // SRAM 3
    logic [31:0] fabric_sram3_a_dout_i;
    logic [9 :0] fabric_sram3_a_addr_o;
    logic [31:0] fabric_sram3_a_bm_o;
    logic [31:0] fabric_sram3_a_din_o;
    logic        fabric_sram3_a_wen_o;
    logic        fabric_sram3_a_men_o;
    logic        fabric_sram3_a_ren_o;
    logic        fabric_sram3_a_clk_o;
    logic        fabric_sram3_a_tie_high_o;
    logic        fabric_sram3_a_tie_low_o;

    // BRAM 0
    logic [15:0] fabric_bram0_a_dout_i;
    logic [9 :0] fabric_bram0_a_addr_o;
    logic [15:0] fabric_bram0_a_bm_o;
    logic [15:0] fabric_bram0_a_din_o;
    logic        fabric_bram0_a_wen_o;
    logic        fabric_bram0_a_men_o;
    logic        fabric_bram0_a_ren_o;
    logic        fabric_bram0_a_clk_o;
    logic        fabric_bram0_a_tie_high_o;
    logic        fabric_bram0_a_tie_low_o;
    logic [15:0] fabric_bram0_b_dout_i;
    logic [9 :0] fabric_bram0_b_addr_o;
    logic [15:0] fabric_bram0_b_bm_o;
    logic [15:0] fabric_bram0_b_din_o;
    logic        fabric_bram0_b_wen_o;
    logic        fabric_bram0_b_men_o;
    logic        fabric_bram0_b_ren_o;
    logic        fabric_bram0_b_clk_o;
    logic        fabric_bram0_b_tie_high_o;
    logic        fabric_bram0_b_tie_low_o;

    // BRAM 1
    logic [15:0] fabric_bram1_a_dout_i;
    logic [9 :0] fabric_bram1_a_addr_o;
    logic [15:0] fabric_bram1_a_bm_o;
    logic [15:0] fabric_bram1_a_din_o;
    logic        fabric_bram1_a_wen_o;
    logic        fabric_bram1_a_men_o;
    logic        fabric_bram1_a_ren_o;
    logic        fabric_bram1_a_clk_o;
    logic        fabric_bram1_a_tie_high_o;
    logic        fabric_bram1_a_tie_low_o;
    logic [15:0] fabric_bram1_b_dout_i;
    logic [9 :0] fabric_bram1_b_addr_o;
    logic [15:0] fabric_bram1_b_bm_o;
    logic [15:0] fabric_bram1_b_din_o;
    logic        fabric_bram1_b_wen_o;
    logic        fabric_bram1_b_men_o;
    logic        fabric_bram1_b_ren_o;
    logic        fabric_bram1_b_clk_o;
    logic        fabric_bram1_b_tie_high_o;
    logic        fabric_bram1_b_tie_low_o;

    // BRAM 2
    logic [15:0] fabric_bram2_a_dout_i;
    logic [9 :0] fabric_bram2_a_addr_o;
    logic [15:0] fabric_bram2_a_bm_o;
    logic [15:0] fabric_bram2_a_din_o;
    logic        fabric_bram2_a_wen_o;
    logic        fabric_bram2_a_men_o;
    logic        fabric_bram2_a_ren_o;
    logic        fabric_bram2_a_clk_o;
    logic        fabric_bram2_a_tie_high_o;
    logic        fabric_bram2_a_tie_low_o;
    logic [15:0] fabric_bram2_b_dout_i;
    logic [9 :0] fabric_bram2_b_addr_o;
    logic [15:0] fabric_bram2_b_bm_o;
    logic [15:0] fabric_bram2_b_din_o;
    logic        fabric_bram2_b_wen_o;
    logic        fabric_bram2_b_men_o;
    logic        fabric_bram2_b_ren_o;
    logic        fabric_bram2_b_clk_o;
    logic        fabric_bram2_b_tie_high_o;
    logic        fabric_bram2_b_tie_low_o;

    // BRAM 3
    logic [15:0] fabric_bram3_a_dout_i;
    logic [9 :0] fabric_bram3_a_addr_o;
    logic [15:0] fabric_bram3_a_bm_o;
    logic [15:0] fabric_bram3_a_din_o;
    logic        fabric_bram3_a_wen_o;
    logic        fabric_bram3_a_men_o;
    logic        fabric_bram3_a_ren_o;
    logic        fabric_bram3_a_clk_o;
    logic        fabric_bram3_a_tie_high_o;
    logic        fabric_bram3_a_tie_low_o;
    logic [15:0] fabric_bram3_b_dout_i;
    logic [9 :0] fabric_bram3_b_addr_o;
    logic [15:0] fabric_bram3_b_bm_o;
    logic [15:0] fabric_bram3_b_din_o;
    logic        fabric_bram3_b_wen_o;
    logic        fabric_bram3_b_men_o;
    logic        fabric_bram3_b_ren_o;
    logic        fabric_bram3_b_clk_o;
    logic        fabric_bram3_b_tie_high_o;
    logic        fabric_bram3_b_tie_low_o;

    eFPGA
    //#(
    //    .MaxFramesPerCol(MaxFramesPerCol),
    //    .FrameBitsPerRow(FrameBitsPerRow)
    //)
    eFPGA
    (
        .FrameData      (FrameData_i),
        .FrameStrobe    (FrameStrobe_i),
        .UserCLK        (clk_i),

        // West I/Os
        .Tile_X0Y1_A_O_top(fabric_io_west_in_i[31]),
        .Tile_X0Y1_A_I_top(fabric_io_west_out_o[31]),
        .Tile_X0Y1_A_T_top(fabric_io_west_oe_o[31]),

        .Tile_X0Y1_B_O_top(fabric_io_west_in_i[30]),
        .Tile_X0Y1_B_I_top(fabric_io_west_out_o[30]),
        .Tile_X0Y1_B_T_top(fabric_io_west_oe_o[30]),

        .Tile_X0Y2_A_O_top(fabric_io_west_in_i[29]),
        .Tile_X0Y2_A_I_top(fabric_io_west_out_o[29]),
        .Tile_X0Y2_A_T_top(fabric_io_west_oe_o[29]),

        .Tile_X0Y2_B_O_top(fabric_io_west_in_i[28]),
        .Tile_X0Y2_B_I_top(fabric_io_west_out_o[28]),
        .Tile_X0Y2_B_T_top(fabric_io_west_oe_o[28]),

        .Tile_X0Y3_A_O_top(fabric_io_west_in_i[27]),
        .Tile_X0Y3_A_I_top(fabric_io_west_out_o[27]),
        .Tile_X0Y3_A_T_top(fabric_io_west_oe_o[27]),

        .Tile_X0Y3_B_O_top(fabric_io_west_in_i[26]),
        .Tile_X0Y3_B_I_top(fabric_io_west_out_o[26]),
        .Tile_X0Y3_B_T_top(fabric_io_west_oe_o[26]),

        .Tile_X0Y4_A_O_top(fabric_io_west_in_i[25]),
        .Tile_X0Y4_A_I_top(fabric_io_west_out_o[25]),
        .Tile_X0Y4_A_T_top(fabric_io_west_oe_o[25]),

        .Tile_X0Y4_B_O_top(fabric_io_west_in_i[24]),
        .Tile_X0Y4_B_I_top(fabric_io_west_out_o[24]),
        .Tile_X0Y4_B_T_top(fabric_io_west_oe_o[24]),

        .Tile_X0Y5_A_O_top(fabric_io_west_in_i[23]),
        .Tile_X0Y5_A_I_top(fabric_io_west_out_o[23]),
        .Tile_X0Y5_A_T_top(fabric_io_west_oe_o[23]),

        .Tile_X0Y5_B_O_top(fabric_io_west_in_i[22]),
        .Tile_X0Y5_B_I_top(fabric_io_west_out_o[22]),
        .Tile_X0Y5_B_T_top(fabric_io_west_oe_o[22]),

        .Tile_X0Y6_A_O_top(fabric_io_west_in_i[21]),
        .Tile_X0Y6_A_I_top(fabric_io_west_out_o[21]),
        .Tile_X0Y6_A_T_top(fabric_io_west_oe_o[21]),

        .Tile_X0Y6_B_O_top(fabric_io_west_in_i[20]),
        .Tile_X0Y6_B_I_top(fabric_io_west_out_o[20]),
        .Tile_X0Y6_B_T_top(fabric_io_west_oe_o[20]),

        .Tile_X0Y7_A_O_top(fabric_io_west_in_i[19]),
        .Tile_X0Y7_A_I_top(fabric_io_west_out_o[19]),
        .Tile_X0Y7_A_T_top(fabric_io_west_oe_o[19]),

        .Tile_X0Y7_B_O_top(fabric_io_west_in_i[18]),
        .Tile_X0Y7_B_I_top(fabric_io_west_out_o[18]),
        .Tile_X0Y7_B_T_top(fabric_io_west_oe_o[18]),

        .Tile_X0Y8_A_O_top(fabric_io_west_in_i[17]),
        .Tile_X0Y8_A_I_top(fabric_io_west_out_o[17]),
        .Tile_X0Y8_A_T_top(fabric_io_west_oe_o[17]),

        .Tile_X0Y8_B_O_top(fabric_io_west_in_i[16]),
        .Tile_X0Y8_B_I_top(fabric_io_west_out_o[16]),
        .Tile_X0Y8_B_T_top(fabric_io_west_oe_o[16]),

        .Tile_X0Y9_A_O_top(fabric_io_west_in_i[15]),
        .Tile_X0Y9_A_I_top(fabric_io_west_out_o[15]),
        .Tile_X0Y9_A_T_top(fabric_io_west_oe_o[15]),

        .Tile_X0Y9_B_O_top(fabric_io_west_in_i[14]),
        .Tile_X0Y9_B_I_top(fabric_io_west_out_o[14]),
        .Tile_X0Y9_B_T_top(fabric_io_west_oe_o[14]),

        .Tile_X0Y10_A_O_top(fabric_io_west_in_i[13]),
        .Tile_X0Y10_A_I_top(fabric_io_west_out_o[13]),
        .Tile_X0Y10_A_T_top(fabric_io_west_oe_o[13]),

        .Tile_X0Y10_B_O_top(fabric_io_west_in_i[12]),
        .Tile_X0Y10_B_I_top(fabric_io_west_out_o[12]),
        .Tile_X0Y10_B_T_top(fabric_io_west_oe_o[12]),

        .Tile_X0Y11_A_O_top(fabric_io_west_in_i[11]),
        .Tile_X0Y11_A_I_top(fabric_io_west_out_o[11]),
        .Tile_X0Y11_A_T_top(fabric_io_west_oe_o[11]),

        .Tile_X0Y11_B_O_top(fabric_io_west_in_i[10]),
        .Tile_X0Y11_B_I_top(fabric_io_west_out_o[10]),
        .Tile_X0Y11_B_T_top(fabric_io_west_oe_o[10]),

        .Tile_X0Y12_A_O_top(fabric_io_west_in_i[9]),
        .Tile_X0Y12_A_I_top(fabric_io_west_out_o[9]),
        .Tile_X0Y12_A_T_top(fabric_io_west_oe_o[9]),

        .Tile_X0Y12_B_O_top(fabric_io_west_in_i[8]),
        .Tile_X0Y12_B_I_top(fabric_io_west_out_o[8]),
        .Tile_X0Y12_B_T_top(fabric_io_west_oe_o[8]),

        .Tile_X0Y13_A_O_top(fabric_io_west_in_i[7]),
        .Tile_X0Y13_A_I_top(fabric_io_west_out_o[7]),
        .Tile_X0Y13_A_T_top(fabric_io_west_oe_o[7]),

        .Tile_X0Y13_B_O_top(fabric_io_west_in_i[6]),
        .Tile_X0Y13_B_I_top(fabric_io_west_out_o[6]),
        .Tile_X0Y13_B_T_top(fabric_io_west_oe_o[6]),

        .Tile_X0Y14_A_O_top(fabric_io_west_in_i[5]),
        .Tile_X0Y14_A_I_top(fabric_io_west_out_o[5]),
        .Tile_X0Y14_A_T_top(fabric_io_west_oe_o[5]),

        .Tile_X0Y14_B_O_top(fabric_io_west_in_i[4]),
        .Tile_X0Y14_B_I_top(fabric_io_west_out_o[4]),
        .Tile_X0Y14_B_T_top(fabric_io_west_oe_o[4]),

        .Tile_X0Y15_A_O_top(fabric_io_west_in_i[3]),
        .Tile_X0Y15_A_I_top(fabric_io_west_out_o[3]),
        .Tile_X0Y15_A_T_top(fabric_io_west_oe_o[3]),

        .Tile_X0Y15_B_O_top(fabric_io_west_in_i[2]),
        .Tile_X0Y15_B_I_top(fabric_io_west_out_o[2]),
        .Tile_X0Y15_B_T_top(fabric_io_west_oe_o[2]),

        .Tile_X0Y16_A_O_top(fabric_io_west_in_i[1]),
        .Tile_X0Y16_A_I_top(fabric_io_west_out_o[1]),
        .Tile_X0Y16_A_T_top(fabric_io_west_oe_o[1]),

        .Tile_X0Y16_B_O_top(fabric_io_west_in_i[0]),
        .Tile_X0Y16_B_I_top(fabric_io_west_out_o[0]),
        .Tile_X0Y16_B_T_top(fabric_io_west_oe_o[0]),

        // WARMBOOT
        .Tile_X1Y17_RESET_top(fabric_warmboot_reset_i),
        .Tile_X1Y17_BOOT_top(fabric_warmboot_boot_o),
        .Tile_X1Y17_SLOT_top0(fabric_warmboot_slot_o[0]),
        .Tile_X1Y17_SLOT_top1(fabric_warmboot_slot_o[1]),
        .Tile_X1Y17_SLOT_top2(fabric_warmboot_slot_o[2]),
        .Tile_X1Y17_SLOT_top3(fabric_warmboot_slot_o[3]),
        .Tile_X1Y17_CONFIGURED_top(configured_i),

        // IRQ
        .Tile_X2Y17_IRQ_top0(fabric_irq_o[0]),
        .Tile_X2Y17_IRQ_top1(fabric_irq_o[1]),
        .Tile_X2Y17_IRQ_top2(fabric_irq_o[2]),
        .Tile_X2Y17_IRQ_top3(fabric_irq_o[3]),
        .Tile_X2Y17_CONFIGURED_top(configured_i),

        // S_XIF 0
        .Tile_X9Y17_ISSUE_READY_top(fabric_issue_ready_o),
        .Tile_X9Y17_ISSUE_ACCEPT_top(fabric_issue_accept_o),
        .Tile_X9Y17_ISSUE_VALID_top(fabric_issue_valid_i),
        .Tile_X9Y17_ISSUE_INSTR_top0(fabric_issue_instr_i[0]),
        .Tile_X9Y17_ISSUE_INSTR_top1(fabric_issue_instr_i[1]),
        .Tile_X9Y17_ISSUE_INSTR_top2(fabric_issue_instr_i[2]),
        .Tile_X9Y17_ISSUE_INSTR_top3(fabric_issue_instr_i[3]),
        .Tile_X9Y17_ISSUE_INSTR_top4(fabric_issue_instr_i[4]),
        .Tile_X9Y17_ISSUE_INSTR_top5(fabric_issue_instr_i[5]),
        .Tile_X9Y17_ISSUE_INSTR_top6(fabric_issue_instr_i[6]),
        .Tile_X9Y17_ISSUE_INSTR_top7(fabric_issue_instr_i[7]),
        .Tile_X9Y17_ISSUE_INSTR_top8(fabric_issue_instr_i[8]),
        .Tile_X9Y17_ISSUE_INSTR_top9(fabric_issue_instr_i[9]),
        .Tile_X9Y17_ISSUE_INSTR_top10(fabric_issue_instr_i[10]),
        .Tile_X9Y17_ISSUE_INSTR_top11(fabric_issue_instr_i[11]),
        .Tile_X9Y17_ISSUE_INSTR_top12(fabric_issue_instr_i[12]),
        .Tile_X9Y17_ISSUE_INSTR_top13(fabric_issue_instr_i[13]),
        .Tile_X9Y17_ISSUE_INSTR_top14(fabric_issue_instr_i[14]),
        .Tile_X9Y17_ISSUE_INSTR_top15(fabric_issue_instr_i[15]),
        .Tile_X9Y17_ISSUE_INSTR_top16(fabric_issue_instr_i[16]),
        .Tile_X9Y17_ISSUE_INSTR_top17(fabric_issue_instr_i[17]),
        .Tile_X9Y17_ISSUE_INSTR_top18(fabric_issue_instr_i[18]),
        .Tile_X9Y17_ISSUE_INSTR_top19(fabric_issue_instr_i[19]),
        .Tile_X9Y17_ISSUE_INSTR_top20(fabric_issue_instr_i[20]),
        .Tile_X9Y17_ISSUE_INSTR_top21(fabric_issue_instr_i[21]),
        .Tile_X9Y17_ISSUE_INSTR_top22(fabric_issue_instr_i[22]),
        .Tile_X9Y17_ISSUE_INSTR_top23(fabric_issue_instr_i[23]),
        .Tile_X9Y17_ISSUE_INSTR_top24(fabric_issue_instr_i[24]),
        .Tile_X9Y17_ISSUE_INSTR_top25(fabric_issue_instr_i[25]),
        .Tile_X9Y17_ISSUE_INSTR_top26(fabric_issue_instr_i[26]),
        .Tile_X9Y17_ISSUE_INSTR_top27(fabric_issue_instr_i[27]),
        .Tile_X9Y17_ISSUE_INSTR_top28(fabric_issue_instr_i[28]),
        .Tile_X9Y17_ISSUE_INSTR_top29(fabric_issue_instr_i[29]),
        .Tile_X9Y17_ISSUE_INSTR_top30(fabric_issue_instr_i[30]),
        .Tile_X9Y17_ISSUE_INSTR_top31(fabric_issue_instr_i[31]),
        .Tile_X9Y17_ISSUE_OPA_top0(fabric_issue_op0_i[0]),
        .Tile_X9Y17_ISSUE_OPA_top1(fabric_issue_op0_i[1]),
        .Tile_X9Y17_ISSUE_OPA_top2(fabric_issue_op0_i[2]),
        .Tile_X9Y17_ISSUE_OPA_top3(fabric_issue_op0_i[3]),
        .Tile_X9Y17_ISSUE_OPA_top4(fabric_issue_op0_i[4]),
        .Tile_X9Y17_ISSUE_OPA_top5(fabric_issue_op0_i[5]),
        .Tile_X9Y17_ISSUE_OPA_top6(fabric_issue_op0_i[6]),
        .Tile_X9Y17_ISSUE_OPA_top7(fabric_issue_op0_i[7]),
        .Tile_X9Y17_ISSUE_OPA_top8(fabric_issue_op0_i[8]),
        .Tile_X9Y17_ISSUE_OPA_top9(fabric_issue_op0_i[9]),
        .Tile_X9Y17_ISSUE_OPA_top10(fabric_issue_op0_i[10]),
        .Tile_X9Y17_ISSUE_OPA_top11(fabric_issue_op0_i[11]),
        .Tile_X9Y17_ISSUE_OPA_top12(fabric_issue_op0_i[12]),
        .Tile_X9Y17_ISSUE_OPA_top13(fabric_issue_op0_i[13]),
        .Tile_X9Y17_ISSUE_OPA_top14(fabric_issue_op0_i[14]),
        .Tile_X9Y17_ISSUE_OPA_top15(fabric_issue_op0_i[15]),
        .Tile_X9Y17_ISSUE_OPA_top16(fabric_issue_op0_i[16]),
        .Tile_X9Y17_ISSUE_OPA_top17(fabric_issue_op0_i[17]),
        .Tile_X9Y17_ISSUE_OPA_top18(fabric_issue_op0_i[18]),
        .Tile_X9Y17_ISSUE_OPA_top19(fabric_issue_op0_i[19]),
        .Tile_X9Y17_ISSUE_OPA_top20(fabric_issue_op0_i[20]),
        .Tile_X9Y17_ISSUE_OPA_top21(fabric_issue_op0_i[21]),
        .Tile_X9Y17_ISSUE_OPA_top22(fabric_issue_op0_i[22]),
        .Tile_X9Y17_ISSUE_OPA_top23(fabric_issue_op0_i[23]),
        .Tile_X9Y17_ISSUE_OPA_top24(fabric_issue_op0_i[24]),
        .Tile_X9Y17_ISSUE_OPA_top25(fabric_issue_op0_i[25]),
        .Tile_X9Y17_ISSUE_OPA_top26(fabric_issue_op0_i[26]),
        .Tile_X9Y17_ISSUE_OPA_top27(fabric_issue_op0_i[27]),
        .Tile_X9Y17_ISSUE_OPA_top28(fabric_issue_op0_i[28]),
        .Tile_X9Y17_ISSUE_OPA_top29(fabric_issue_op0_i[29]),
        .Tile_X9Y17_ISSUE_OPA_top30(fabric_issue_op0_i[30]),
        .Tile_X9Y17_ISSUE_OPA_top31(fabric_issue_op0_i[31]),
        .Tile_X9Y17_ISSUE_OPB_top0(fabric_issue_op1_i[0]),
        .Tile_X9Y17_ISSUE_OPB_top1(fabric_issue_op1_i[1]),
        .Tile_X9Y17_ISSUE_OPB_top2(fabric_issue_op1_i[2]),
        .Tile_X9Y17_ISSUE_OPB_top3(fabric_issue_op1_i[3]),
        .Tile_X9Y17_ISSUE_OPB_top4(fabric_issue_op1_i[4]),
        .Tile_X9Y17_ISSUE_OPB_top5(fabric_issue_op1_i[5]),
        .Tile_X9Y17_ISSUE_OPB_top6(fabric_issue_op1_i[6]),
        .Tile_X9Y17_ISSUE_OPB_top7(fabric_issue_op1_i[7]),
        .Tile_X9Y17_ISSUE_OPB_top8(fabric_issue_op1_i[8]),
        .Tile_X9Y17_ISSUE_OPB_top9(fabric_issue_op1_i[9]),
        .Tile_X9Y17_ISSUE_OPB_top10(fabric_issue_op1_i[10]),
        .Tile_X9Y17_ISSUE_OPB_top11(fabric_issue_op1_i[11]),
        .Tile_X9Y17_ISSUE_OPB_top12(fabric_issue_op1_i[12]),
        .Tile_X9Y17_ISSUE_OPB_top13(fabric_issue_op1_i[13]),
        .Tile_X9Y17_ISSUE_OPB_top14(fabric_issue_op1_i[14]),
        .Tile_X9Y17_ISSUE_OPB_top15(fabric_issue_op1_i[15]),
        .Tile_X9Y17_ISSUE_OPB_top16(fabric_issue_op1_i[16]),
        .Tile_X9Y17_ISSUE_OPB_top17(fabric_issue_op1_i[17]),
        .Tile_X9Y17_ISSUE_OPB_top18(fabric_issue_op1_i[18]),
        .Tile_X9Y17_ISSUE_OPB_top19(fabric_issue_op1_i[19]),
        .Tile_X9Y17_ISSUE_OPB_top20(fabric_issue_op1_i[20]),
        .Tile_X9Y17_ISSUE_OPB_top21(fabric_issue_op1_i[21]),
        .Tile_X9Y17_ISSUE_OPB_top22(fabric_issue_op1_i[22]),
        .Tile_X9Y17_ISSUE_OPB_top23(fabric_issue_op1_i[23]),
        .Tile_X9Y17_ISSUE_OPB_top24(fabric_issue_op1_i[24]),
        .Tile_X9Y17_ISSUE_OPB_top25(fabric_issue_op1_i[25]),
        .Tile_X9Y17_ISSUE_OPB_top26(fabric_issue_op1_i[26]),
        .Tile_X9Y17_ISSUE_OPB_top27(fabric_issue_op1_i[27]),
        .Tile_X9Y17_ISSUE_OPB_top28(fabric_issue_op1_i[28]),
        .Tile_X9Y17_ISSUE_OPB_top29(fabric_issue_op1_i[29]),
        .Tile_X9Y17_ISSUE_OPB_top30(fabric_issue_op1_i[30]),
        .Tile_X9Y17_ISSUE_OPB_top31(fabric_issue_op1_i[31]),
        .Tile_X9Y17_ISSUE_ID_top0(fabric_issue_id_i[0]),
        .Tile_X9Y17_ISSUE_ID_top1(fabric_issue_id_i[1]),
        .Tile_X9Y17_ISSUE_ID_top2(fabric_issue_id_i[2]),
        .Tile_X9Y17_ISSUE_ID_top3(fabric_issue_id_i[3]),
        .Tile_X9Y17_RESULT_VALID_top(fabric_result_valid_o),
        .Tile_X9Y17_RESULT_ID_top0(fabric_result_id_o[0]),
        .Tile_X9Y17_RESULT_ID_top1(fabric_result_id_o[1]),
        .Tile_X9Y17_RESULT_ID_top2(fabric_result_id_o[2]),
        .Tile_X9Y17_RESULT_ID_top3(fabric_result_id_o[3]),
        .Tile_X9Y17_RESULT_RD_top0(fabric_result_rd_o[0]),
        .Tile_X9Y17_RESULT_RD_top1(fabric_result_rd_o[1]),
        .Tile_X9Y17_RESULT_RD_top2(fabric_result_rd_o[2]),
        .Tile_X9Y17_RESULT_RD_top3(fabric_result_rd_o[3]),
        .Tile_X9Y17_RESULT_RD_top4(fabric_result_rd_o[4]),
        .Tile_X9Y17_RESULT_top0(fabric_result_o[0]),
        .Tile_X9Y17_RESULT_top1(fabric_result_o[1]),
        .Tile_X9Y17_RESULT_top2(fabric_result_o[2]),
        .Tile_X9Y17_RESULT_top3(fabric_result_o[3]),
        .Tile_X9Y17_RESULT_top4(fabric_result_o[4]),
        .Tile_X9Y17_RESULT_top5(fabric_result_o[5]),
        .Tile_X9Y17_RESULT_top6(fabric_result_o[6]),
        .Tile_X9Y17_RESULT_top7(fabric_result_o[7]),
        .Tile_X9Y17_RESULT_top8(fabric_result_o[8]),
        .Tile_X9Y17_RESULT_top9(fabric_result_o[9]),
        .Tile_X9Y17_RESULT_top10(fabric_result_o[10]),
        .Tile_X9Y17_RESULT_top11(fabric_result_o[11]),
        .Tile_X9Y17_RESULT_top12(fabric_result_o[12]),
        .Tile_X9Y17_RESULT_top13(fabric_result_o[13]),
        .Tile_X9Y17_RESULT_top14(fabric_result_o[14]),
        .Tile_X9Y17_RESULT_top15(fabric_result_o[15]),
        .Tile_X9Y17_RESULT_top16(fabric_result_o[16]),
        .Tile_X9Y17_RESULT_top17(fabric_result_o[17]),
        .Tile_X9Y17_RESULT_top18(fabric_result_o[18]),
        .Tile_X9Y17_RESULT_top19(fabric_result_o[19]),
        .Tile_X9Y17_RESULT_top20(fabric_result_o[20]),
        .Tile_X9Y17_RESULT_top21(fabric_result_o[21]),
        .Tile_X9Y17_RESULT_top22(fabric_result_o[22]),
        .Tile_X9Y17_RESULT_top23(fabric_result_o[23]),
        .Tile_X9Y17_RESULT_top24(fabric_result_o[24]),
        .Tile_X9Y17_RESULT_top25(fabric_result_o[25]),
        .Tile_X9Y17_RESULT_top26(fabric_result_o[26]),
        .Tile_X9Y17_RESULT_top27(fabric_result_o[27]),
        .Tile_X9Y17_RESULT_top28(fabric_result_o[28]),
        .Tile_X9Y17_RESULT_top29(fabric_result_o[29]),
        .Tile_X9Y17_RESULT_top30(fabric_result_o[30]),
        .Tile_X9Y17_RESULT_top31(fabric_result_o[31]),

        // S_OBI 0
        .Tile_X5Y17_REQ_top(fabric_obi_req_i),
        .Tile_X5Y17_WE_top(fabric_obi_we_i),
        .Tile_X5Y17_BE_top0(fabric_obi_be_i[0]),
        .Tile_X5Y17_BE_top1(fabric_obi_be_i[1]),
        .Tile_X5Y17_BE_top2(fabric_obi_be_i[2]),
        .Tile_X5Y17_BE_top3(fabric_obi_be_i[3]),
        .Tile_X5Y17_ADDR_top0(fabric_obi_addr_i[0]),
        .Tile_X5Y17_ADDR_top1(fabric_obi_addr_i[1]),
        .Tile_X5Y17_ADDR_top2(fabric_obi_addr_i[2]),
        .Tile_X5Y17_ADDR_top3(fabric_obi_addr_i[3]),
        .Tile_X5Y17_ADDR_top4(fabric_obi_addr_i[4]),
        .Tile_X5Y17_ADDR_top5(fabric_obi_addr_i[5]),
        .Tile_X5Y17_ADDR_top6(fabric_obi_addr_i[6]),
        .Tile_X5Y17_ADDR_top7(fabric_obi_addr_i[7]),
        .Tile_X5Y17_ADDR_top8(fabric_obi_addr_i[8]),
        .Tile_X5Y17_ADDR_top9(fabric_obi_addr_i[9]),
        .Tile_X5Y17_ADDR_top10(fabric_obi_addr_i[10]),
        .Tile_X5Y17_ADDR_top11(fabric_obi_addr_i[11]),
        .Tile_X5Y17_ADDR_top12(fabric_obi_addr_i[12]),
        .Tile_X5Y17_ADDR_top13(fabric_obi_addr_i[13]),
        .Tile_X5Y17_ADDR_top14(fabric_obi_addr_i[14]),
        .Tile_X5Y17_ADDR_top15(fabric_obi_addr_i[15]),
        .Tile_X5Y17_ADDR_top16(fabric_obi_addr_i[16]),
        .Tile_X5Y17_ADDR_top17(fabric_obi_addr_i[17]),
        .Tile_X5Y17_ADDR_top18(fabric_obi_addr_i[18]),
        .Tile_X5Y17_ADDR_top19(fabric_obi_addr_i[19]),
        .Tile_X5Y17_ADDR_top20(fabric_obi_addr_i[20]),
        .Tile_X5Y17_ADDR_top21(fabric_obi_addr_i[21]),
        .Tile_X5Y17_ADDR_top22(fabric_obi_addr_i[22]),
        .Tile_X5Y17_ADDR_top23(fabric_obi_addr_i[23]),
        .Tile_X5Y17_WDATA_top0(fabric_obi_wdata_i[0]),
        .Tile_X5Y17_WDATA_top1(fabric_obi_wdata_i[1]),
        .Tile_X5Y17_WDATA_top2(fabric_obi_wdata_i[2]),
        .Tile_X5Y17_WDATA_top3(fabric_obi_wdata_i[3]),
        .Tile_X5Y17_WDATA_top4(fabric_obi_wdata_i[4]),
        .Tile_X5Y17_WDATA_top5(fabric_obi_wdata_i[5]),
        .Tile_X5Y17_WDATA_top6(fabric_obi_wdata_i[6]),
        .Tile_X5Y17_WDATA_top7(fabric_obi_wdata_i[7]),
        .Tile_X5Y17_WDATA_top8(fabric_obi_wdata_i[8]),
        .Tile_X5Y17_WDATA_top9(fabric_obi_wdata_i[9]),
        .Tile_X5Y17_WDATA_top10(fabric_obi_wdata_i[10]),
        .Tile_X5Y17_WDATA_top11(fabric_obi_wdata_i[11]),
        .Tile_X5Y17_WDATA_top12(fabric_obi_wdata_i[12]),
        .Tile_X5Y17_WDATA_top13(fabric_obi_wdata_i[13]),
        .Tile_X5Y17_WDATA_top14(fabric_obi_wdata_i[14]),
        .Tile_X5Y17_WDATA_top15(fabric_obi_wdata_i[15]),
        .Tile_X5Y17_WDATA_top16(fabric_obi_wdata_i[16]),
        .Tile_X5Y17_WDATA_top17(fabric_obi_wdata_i[17]),
        .Tile_X5Y17_WDATA_top18(fabric_obi_wdata_i[18]),
        .Tile_X5Y17_WDATA_top19(fabric_obi_wdata_i[19]),
        .Tile_X5Y17_WDATA_top20(fabric_obi_wdata_i[20]),
        .Tile_X5Y17_WDATA_top21(fabric_obi_wdata_i[21]),
        .Tile_X5Y17_WDATA_top22(fabric_obi_wdata_i[22]),
        .Tile_X5Y17_WDATA_top23(fabric_obi_wdata_i[23]),
        .Tile_X5Y17_WDATA_top24(fabric_obi_wdata_i[24]),
        .Tile_X5Y17_WDATA_top25(fabric_obi_wdata_i[25]),
        .Tile_X5Y17_WDATA_top26(fabric_obi_wdata_i[26]),
        .Tile_X5Y17_WDATA_top27(fabric_obi_wdata_i[27]),
        .Tile_X5Y17_WDATA_top28(fabric_obi_wdata_i[28]),
        .Tile_X5Y17_WDATA_top29(fabric_obi_wdata_i[29]),
        .Tile_X5Y17_WDATA_top30(fabric_obi_wdata_i[30]),
        .Tile_X5Y17_WDATA_top31(fabric_obi_wdata_i[31]),
        .Tile_X5Y17_GNT_top(fabric_obi_gnt_o),
        .Tile_X5Y17_RVALID_top(fabric_obi_rvalid_o),
        .Tile_X5Y17_RDATA_top0(fabric_obi_rdata_o[0]),
        .Tile_X5Y17_RDATA_top1(fabric_obi_rdata_o[1]),
        .Tile_X5Y17_RDATA_top2(fabric_obi_rdata_o[2]),
        .Tile_X5Y17_RDATA_top3(fabric_obi_rdata_o[3]),
        .Tile_X5Y17_RDATA_top4(fabric_obi_rdata_o[4]),
        .Tile_X5Y17_RDATA_top5(fabric_obi_rdata_o[5]),
        .Tile_X5Y17_RDATA_top6(fabric_obi_rdata_o[6]),
        .Tile_X5Y17_RDATA_top7(fabric_obi_rdata_o[7]),
        .Tile_X5Y17_RDATA_top8(fabric_obi_rdata_o[8]),
        .Tile_X5Y17_RDATA_top9(fabric_obi_rdata_o[9]),
        .Tile_X5Y17_RDATA_top10(fabric_obi_rdata_o[10]),
        .Tile_X5Y17_RDATA_top11(fabric_obi_rdata_o[11]),
        .Tile_X5Y17_RDATA_top12(fabric_obi_rdata_o[12]),
        .Tile_X5Y17_RDATA_top13(fabric_obi_rdata_o[13]),
        .Tile_X5Y17_RDATA_top14(fabric_obi_rdata_o[14]),
        .Tile_X5Y17_RDATA_top15(fabric_obi_rdata_o[15]),
        .Tile_X5Y17_RDATA_top16(fabric_obi_rdata_o[16]),
        .Tile_X5Y17_RDATA_top17(fabric_obi_rdata_o[17]),
        .Tile_X5Y17_RDATA_top18(fabric_obi_rdata_o[18]),
        .Tile_X5Y17_RDATA_top19(fabric_obi_rdata_o[19]),
        .Tile_X5Y17_RDATA_top20(fabric_obi_rdata_o[20]),
        .Tile_X5Y17_RDATA_top21(fabric_obi_rdata_o[21]),
        .Tile_X5Y17_RDATA_top22(fabric_obi_rdata_o[22]),
        .Tile_X5Y17_RDATA_top23(fabric_obi_rdata_o[23]),
        .Tile_X5Y17_RDATA_top24(fabric_obi_rdata_o[24]),
        .Tile_X5Y17_RDATA_top25(fabric_obi_rdata_o[25]),
        .Tile_X5Y17_RDATA_top26(fabric_obi_rdata_o[26]),
        .Tile_X5Y17_RDATA_top27(fabric_obi_rdata_o[27]),
        .Tile_X5Y17_RDATA_top28(fabric_obi_rdata_o[28]),
        .Tile_X5Y17_RDATA_top29(fabric_obi_rdata_o[29]),
        .Tile_X5Y17_RDATA_top30(fabric_obi_rdata_o[30]),
        .Tile_X5Y17_RDATA_top31(fabric_obi_rdata_o[31]),

        // SRAM 0
        .Tile_X11Y10_A_DOUT_SRAM0(fabric_sram0_a_dout_i[0]),
        .Tile_X11Y10_A_DOUT_SRAM1(fabric_sram0_a_dout_i[1]),
        .Tile_X11Y10_A_DOUT_SRAM2(fabric_sram0_a_dout_i[2]),
        .Tile_X11Y10_A_DOUT_SRAM3(fabric_sram0_a_dout_i[3]),
        .Tile_X11Y10_A_DOUT_SRAM4(fabric_sram0_a_dout_i[4]),
        .Tile_X11Y10_A_DOUT_SRAM5(fabric_sram0_a_dout_i[5]),
        .Tile_X11Y10_A_DOUT_SRAM6(fabric_sram0_a_dout_i[6]),
        .Tile_X11Y10_A_DOUT_SRAM7(fabric_sram0_a_dout_i[7]),
        .Tile_X11Y10_A_DOUT_SRAM8(fabric_sram0_a_dout_i[8]),
        .Tile_X11Y10_A_DOUT_SRAM9(fabric_sram0_a_dout_i[9]),
        .Tile_X11Y10_A_DOUT_SRAM10(fabric_sram0_a_dout_i[10]),
        .Tile_X11Y10_A_DOUT_SRAM11(fabric_sram0_a_dout_i[11]),
        .Tile_X11Y10_A_DOUT_SRAM12(fabric_sram0_a_dout_i[12]),
        .Tile_X11Y10_A_DOUT_SRAM13(fabric_sram0_a_dout_i[13]),
        .Tile_X11Y10_A_DOUT_SRAM14(fabric_sram0_a_dout_i[14]),
        .Tile_X11Y10_A_DOUT_SRAM15(fabric_sram0_a_dout_i[15]),
        .Tile_X11Y10_A_DOUT_SRAM16(fabric_sram0_a_dout_i[16]),
        .Tile_X11Y10_A_DOUT_SRAM17(fabric_sram0_a_dout_i[17]),
        .Tile_X11Y10_A_DOUT_SRAM18(fabric_sram0_a_dout_i[18]),
        .Tile_X11Y10_A_DOUT_SRAM19(fabric_sram0_a_dout_i[19]),
        .Tile_X11Y10_A_DOUT_SRAM20(fabric_sram0_a_dout_i[20]),
        .Tile_X11Y10_A_DOUT_SRAM21(fabric_sram0_a_dout_i[21]),
        .Tile_X11Y10_A_DOUT_SRAM22(fabric_sram0_a_dout_i[22]),
        .Tile_X11Y10_A_DOUT_SRAM23(fabric_sram0_a_dout_i[23]),
        .Tile_X11Y10_A_DOUT_SRAM24(fabric_sram0_a_dout_i[24]),
        .Tile_X11Y10_A_DOUT_SRAM25(fabric_sram0_a_dout_i[25]),
        .Tile_X11Y10_A_DOUT_SRAM26(fabric_sram0_a_dout_i[26]),
        .Tile_X11Y10_A_DOUT_SRAM27(fabric_sram0_a_dout_i[27]),
        .Tile_X11Y10_A_DOUT_SRAM28(fabric_sram0_a_dout_i[28]),
        .Tile_X11Y10_A_DOUT_SRAM29(fabric_sram0_a_dout_i[29]),
        .Tile_X11Y10_A_DOUT_SRAM30(fabric_sram0_a_dout_i[30]),
        .Tile_X11Y10_A_DOUT_SRAM31(fabric_sram0_a_dout_i[31]),
        .Tile_X11Y10_A_ADDR_SRAM0(fabric_sram0_a_addr_o[0]),
        .Tile_X11Y10_A_ADDR_SRAM1(fabric_sram0_a_addr_o[1]),
        .Tile_X11Y10_A_ADDR_SRAM2(fabric_sram0_a_addr_o[2]),
        .Tile_X11Y10_A_ADDR_SRAM3(fabric_sram0_a_addr_o[3]),
        .Tile_X11Y10_A_ADDR_SRAM4(fabric_sram0_a_addr_o[4]),
        .Tile_X11Y10_A_ADDR_SRAM5(fabric_sram0_a_addr_o[5]),
        .Tile_X11Y10_A_ADDR_SRAM6(fabric_sram0_a_addr_o[6]),
        .Tile_X11Y10_A_ADDR_SRAM7(fabric_sram0_a_addr_o[7]),
        .Tile_X11Y10_A_ADDR_SRAM8(fabric_sram0_a_addr_o[8]),
        .Tile_X11Y10_A_ADDR_SRAM9(fabric_sram0_a_addr_o[9]),
        .Tile_X11Y10_A_BM_SRAM0(fabric_sram0_a_bm_o[0]),
        .Tile_X11Y10_A_BM_SRAM1(fabric_sram0_a_bm_o[1]),
        .Tile_X11Y10_A_BM_SRAM2(fabric_sram0_a_bm_o[2]),
        .Tile_X11Y10_A_BM_SRAM3(fabric_sram0_a_bm_o[3]),
        .Tile_X11Y10_A_BM_SRAM4(fabric_sram0_a_bm_o[4]),
        .Tile_X11Y10_A_BM_SRAM5(fabric_sram0_a_bm_o[5]),
        .Tile_X11Y10_A_BM_SRAM6(fabric_sram0_a_bm_o[6]),
        .Tile_X11Y10_A_BM_SRAM7(fabric_sram0_a_bm_o[7]),
        .Tile_X11Y10_A_BM_SRAM8(fabric_sram0_a_bm_o[8]),
        .Tile_X11Y10_A_BM_SRAM9(fabric_sram0_a_bm_o[9]),
        .Tile_X11Y10_A_BM_SRAM10(fabric_sram0_a_bm_o[10]),
        .Tile_X11Y10_A_BM_SRAM11(fabric_sram0_a_bm_o[11]),
        .Tile_X11Y10_A_BM_SRAM12(fabric_sram0_a_bm_o[12]),
        .Tile_X11Y10_A_BM_SRAM13(fabric_sram0_a_bm_o[13]),
        .Tile_X11Y10_A_BM_SRAM14(fabric_sram0_a_bm_o[14]),
        .Tile_X11Y10_A_BM_SRAM15(fabric_sram0_a_bm_o[15]),
        .Tile_X11Y10_A_BM_SRAM16(fabric_sram0_a_bm_o[16]),
        .Tile_X11Y10_A_BM_SRAM17(fabric_sram0_a_bm_o[17]),
        .Tile_X11Y10_A_BM_SRAM18(fabric_sram0_a_bm_o[18]),
        .Tile_X11Y10_A_BM_SRAM19(fabric_sram0_a_bm_o[19]),
        .Tile_X11Y10_A_BM_SRAM20(fabric_sram0_a_bm_o[20]),
        .Tile_X11Y10_A_BM_SRAM21(fabric_sram0_a_bm_o[21]),
        .Tile_X11Y10_A_BM_SRAM22(fabric_sram0_a_bm_o[22]),
        .Tile_X11Y10_A_BM_SRAM23(fabric_sram0_a_bm_o[23]),
        .Tile_X11Y10_A_BM_SRAM24(fabric_sram0_a_bm_o[24]),
        .Tile_X11Y10_A_BM_SRAM25(fabric_sram0_a_bm_o[25]),
        .Tile_X11Y10_A_BM_SRAM26(fabric_sram0_a_bm_o[26]),
        .Tile_X11Y10_A_BM_SRAM27(fabric_sram0_a_bm_o[27]),
        .Tile_X11Y10_A_BM_SRAM28(fabric_sram0_a_bm_o[28]),
        .Tile_X11Y10_A_BM_SRAM29(fabric_sram0_a_bm_o[29]),
        .Tile_X11Y10_A_BM_SRAM30(fabric_sram0_a_bm_o[30]),
        .Tile_X11Y10_A_BM_SRAM31(fabric_sram0_a_bm_o[31]),
        .Tile_X11Y10_A_DIN_SRAM0(fabric_sram0_a_din_o[0]),
        .Tile_X11Y10_A_DIN_SRAM1(fabric_sram0_a_din_o[1]),
        .Tile_X11Y10_A_DIN_SRAM2(fabric_sram0_a_din_o[2]),
        .Tile_X11Y10_A_DIN_SRAM3(fabric_sram0_a_din_o[3]),
        .Tile_X11Y10_A_DIN_SRAM4(fabric_sram0_a_din_o[4]),
        .Tile_X11Y10_A_DIN_SRAM5(fabric_sram0_a_din_o[5]),
        .Tile_X11Y10_A_DIN_SRAM6(fabric_sram0_a_din_o[6]),
        .Tile_X11Y10_A_DIN_SRAM7(fabric_sram0_a_din_o[7]),
        .Tile_X11Y10_A_DIN_SRAM8(fabric_sram0_a_din_o[8]),
        .Tile_X11Y10_A_DIN_SRAM9(fabric_sram0_a_din_o[9]),
        .Tile_X11Y10_A_DIN_SRAM10(fabric_sram0_a_din_o[10]),
        .Tile_X11Y10_A_DIN_SRAM11(fabric_sram0_a_din_o[11]),
        .Tile_X11Y10_A_DIN_SRAM12(fabric_sram0_a_din_o[12]),
        .Tile_X11Y10_A_DIN_SRAM13(fabric_sram0_a_din_o[13]),
        .Tile_X11Y10_A_DIN_SRAM14(fabric_sram0_a_din_o[14]),
        .Tile_X11Y10_A_DIN_SRAM15(fabric_sram0_a_din_o[15]),
        .Tile_X11Y10_A_DIN_SRAM16(fabric_sram0_a_din_o[16]),
        .Tile_X11Y10_A_DIN_SRAM17(fabric_sram0_a_din_o[17]),
        .Tile_X11Y10_A_DIN_SRAM18(fabric_sram0_a_din_o[18]),
        .Tile_X11Y10_A_DIN_SRAM19(fabric_sram0_a_din_o[19]),
        .Tile_X11Y10_A_DIN_SRAM20(fabric_sram0_a_din_o[20]),
        .Tile_X11Y10_A_DIN_SRAM21(fabric_sram0_a_din_o[21]),
        .Tile_X11Y10_A_DIN_SRAM22(fabric_sram0_a_din_o[22]),
        .Tile_X11Y10_A_DIN_SRAM23(fabric_sram0_a_din_o[23]),
        .Tile_X11Y10_A_DIN_SRAM24(fabric_sram0_a_din_o[24]),
        .Tile_X11Y10_A_DIN_SRAM25(fabric_sram0_a_din_o[25]),
        .Tile_X11Y10_A_DIN_SRAM26(fabric_sram0_a_din_o[26]),
        .Tile_X11Y10_A_DIN_SRAM27(fabric_sram0_a_din_o[27]),
        .Tile_X11Y10_A_DIN_SRAM28(fabric_sram0_a_din_o[28]),
        .Tile_X11Y10_A_DIN_SRAM29(fabric_sram0_a_din_o[29]),
        .Tile_X11Y10_A_DIN_SRAM30(fabric_sram0_a_din_o[30]),
        .Tile_X11Y10_A_DIN_SRAM31(fabric_sram0_a_din_o[31]),
        .Tile_X11Y10_A_WEN_SRAM(fabric_sram0_a_wen_o),
        .Tile_X11Y10_A_MEN_SRAM(fabric_sram0_a_men_o),
        .Tile_X11Y10_A_REN_SRAM(fabric_sram0_a_ren_o),
        .Tile_X11Y10_A_CLK_SRAM(fabric_sram0_a_clk_o),
        .Tile_X11Y10_A_TIE_HIGH_SRAM(fabric_sram0_a_tie_high_o),
        .Tile_X11Y10_A_TIE_LOW_SRAM(fabric_sram0_a_tie_low_o),
        .Tile_X11Y10_CONFIGURED_top(configured_i),

        // SRAM 1
        .Tile_X11Y12_A_DOUT_SRAM0(fabric_sram1_a_dout_i[0]),
        .Tile_X11Y12_A_DOUT_SRAM1(fabric_sram1_a_dout_i[1]),
        .Tile_X11Y12_A_DOUT_SRAM2(fabric_sram1_a_dout_i[2]),
        .Tile_X11Y12_A_DOUT_SRAM3(fabric_sram1_a_dout_i[3]),
        .Tile_X11Y12_A_DOUT_SRAM4(fabric_sram1_a_dout_i[4]),
        .Tile_X11Y12_A_DOUT_SRAM5(fabric_sram1_a_dout_i[5]),
        .Tile_X11Y12_A_DOUT_SRAM6(fabric_sram1_a_dout_i[6]),
        .Tile_X11Y12_A_DOUT_SRAM7(fabric_sram1_a_dout_i[7]),
        .Tile_X11Y12_A_DOUT_SRAM8(fabric_sram1_a_dout_i[8]),
        .Tile_X11Y12_A_DOUT_SRAM9(fabric_sram1_a_dout_i[9]),
        .Tile_X11Y12_A_DOUT_SRAM10(fabric_sram1_a_dout_i[10]),
        .Tile_X11Y12_A_DOUT_SRAM11(fabric_sram1_a_dout_i[11]),
        .Tile_X11Y12_A_DOUT_SRAM12(fabric_sram1_a_dout_i[12]),
        .Tile_X11Y12_A_DOUT_SRAM13(fabric_sram1_a_dout_i[13]),
        .Tile_X11Y12_A_DOUT_SRAM14(fabric_sram1_a_dout_i[14]),
        .Tile_X11Y12_A_DOUT_SRAM15(fabric_sram1_a_dout_i[15]),
        .Tile_X11Y12_A_DOUT_SRAM16(fabric_sram1_a_dout_i[16]),
        .Tile_X11Y12_A_DOUT_SRAM17(fabric_sram1_a_dout_i[17]),
        .Tile_X11Y12_A_DOUT_SRAM18(fabric_sram1_a_dout_i[18]),
        .Tile_X11Y12_A_DOUT_SRAM19(fabric_sram1_a_dout_i[19]),
        .Tile_X11Y12_A_DOUT_SRAM20(fabric_sram1_a_dout_i[20]),
        .Tile_X11Y12_A_DOUT_SRAM21(fabric_sram1_a_dout_i[21]),
        .Tile_X11Y12_A_DOUT_SRAM22(fabric_sram1_a_dout_i[22]),
        .Tile_X11Y12_A_DOUT_SRAM23(fabric_sram1_a_dout_i[23]),
        .Tile_X11Y12_A_DOUT_SRAM24(fabric_sram1_a_dout_i[24]),
        .Tile_X11Y12_A_DOUT_SRAM25(fabric_sram1_a_dout_i[25]),
        .Tile_X11Y12_A_DOUT_SRAM26(fabric_sram1_a_dout_i[26]),
        .Tile_X11Y12_A_DOUT_SRAM27(fabric_sram1_a_dout_i[27]),
        .Tile_X11Y12_A_DOUT_SRAM28(fabric_sram1_a_dout_i[28]),
        .Tile_X11Y12_A_DOUT_SRAM29(fabric_sram1_a_dout_i[29]),
        .Tile_X11Y12_A_DOUT_SRAM30(fabric_sram1_a_dout_i[30]),
        .Tile_X11Y12_A_DOUT_SRAM31(fabric_sram1_a_dout_i[31]),
        .Tile_X11Y12_A_ADDR_SRAM0(fabric_sram1_a_addr_o[0]),
        .Tile_X11Y12_A_ADDR_SRAM1(fabric_sram1_a_addr_o[1]),
        .Tile_X11Y12_A_ADDR_SRAM2(fabric_sram1_a_addr_o[2]),
        .Tile_X11Y12_A_ADDR_SRAM3(fabric_sram1_a_addr_o[3]),
        .Tile_X11Y12_A_ADDR_SRAM4(fabric_sram1_a_addr_o[4]),
        .Tile_X11Y12_A_ADDR_SRAM5(fabric_sram1_a_addr_o[5]),
        .Tile_X11Y12_A_ADDR_SRAM6(fabric_sram1_a_addr_o[6]),
        .Tile_X11Y12_A_ADDR_SRAM7(fabric_sram1_a_addr_o[7]),
        .Tile_X11Y12_A_ADDR_SRAM8(fabric_sram1_a_addr_o[8]),
        .Tile_X11Y12_A_ADDR_SRAM9(fabric_sram1_a_addr_o[9]),
        .Tile_X11Y12_A_BM_SRAM0(fabric_sram1_a_bm_o[0]),
        .Tile_X11Y12_A_BM_SRAM1(fabric_sram1_a_bm_o[1]),
        .Tile_X11Y12_A_BM_SRAM2(fabric_sram1_a_bm_o[2]),
        .Tile_X11Y12_A_BM_SRAM3(fabric_sram1_a_bm_o[3]),
        .Tile_X11Y12_A_BM_SRAM4(fabric_sram1_a_bm_o[4]),
        .Tile_X11Y12_A_BM_SRAM5(fabric_sram1_a_bm_o[5]),
        .Tile_X11Y12_A_BM_SRAM6(fabric_sram1_a_bm_o[6]),
        .Tile_X11Y12_A_BM_SRAM7(fabric_sram1_a_bm_o[7]),
        .Tile_X11Y12_A_BM_SRAM8(fabric_sram1_a_bm_o[8]),
        .Tile_X11Y12_A_BM_SRAM9(fabric_sram1_a_bm_o[9]),
        .Tile_X11Y12_A_BM_SRAM10(fabric_sram1_a_bm_o[10]),
        .Tile_X11Y12_A_BM_SRAM11(fabric_sram1_a_bm_o[11]),
        .Tile_X11Y12_A_BM_SRAM12(fabric_sram1_a_bm_o[12]),
        .Tile_X11Y12_A_BM_SRAM13(fabric_sram1_a_bm_o[13]),
        .Tile_X11Y12_A_BM_SRAM14(fabric_sram1_a_bm_o[14]),
        .Tile_X11Y12_A_BM_SRAM15(fabric_sram1_a_bm_o[15]),
        .Tile_X11Y12_A_BM_SRAM16(fabric_sram1_a_bm_o[16]),
        .Tile_X11Y12_A_BM_SRAM17(fabric_sram1_a_bm_o[17]),
        .Tile_X11Y12_A_BM_SRAM18(fabric_sram1_a_bm_o[18]),
        .Tile_X11Y12_A_BM_SRAM19(fabric_sram1_a_bm_o[19]),
        .Tile_X11Y12_A_BM_SRAM20(fabric_sram1_a_bm_o[20]),
        .Tile_X11Y12_A_BM_SRAM21(fabric_sram1_a_bm_o[21]),
        .Tile_X11Y12_A_BM_SRAM22(fabric_sram1_a_bm_o[22]),
        .Tile_X11Y12_A_BM_SRAM23(fabric_sram1_a_bm_o[23]),
        .Tile_X11Y12_A_BM_SRAM24(fabric_sram1_a_bm_o[24]),
        .Tile_X11Y12_A_BM_SRAM25(fabric_sram1_a_bm_o[25]),
        .Tile_X11Y12_A_BM_SRAM26(fabric_sram1_a_bm_o[26]),
        .Tile_X11Y12_A_BM_SRAM27(fabric_sram1_a_bm_o[27]),
        .Tile_X11Y12_A_BM_SRAM28(fabric_sram1_a_bm_o[28]),
        .Tile_X11Y12_A_BM_SRAM29(fabric_sram1_a_bm_o[29]),
        .Tile_X11Y12_A_BM_SRAM30(fabric_sram1_a_bm_o[30]),
        .Tile_X11Y12_A_BM_SRAM31(fabric_sram1_a_bm_o[31]),
        .Tile_X11Y12_A_DIN_SRAM0(fabric_sram1_a_din_o[0]),
        .Tile_X11Y12_A_DIN_SRAM1(fabric_sram1_a_din_o[1]),
        .Tile_X11Y12_A_DIN_SRAM2(fabric_sram1_a_din_o[2]),
        .Tile_X11Y12_A_DIN_SRAM3(fabric_sram1_a_din_o[3]),
        .Tile_X11Y12_A_DIN_SRAM4(fabric_sram1_a_din_o[4]),
        .Tile_X11Y12_A_DIN_SRAM5(fabric_sram1_a_din_o[5]),
        .Tile_X11Y12_A_DIN_SRAM6(fabric_sram1_a_din_o[6]),
        .Tile_X11Y12_A_DIN_SRAM7(fabric_sram1_a_din_o[7]),
        .Tile_X11Y12_A_DIN_SRAM8(fabric_sram1_a_din_o[8]),
        .Tile_X11Y12_A_DIN_SRAM9(fabric_sram1_a_din_o[9]),
        .Tile_X11Y12_A_DIN_SRAM10(fabric_sram1_a_din_o[10]),
        .Tile_X11Y12_A_DIN_SRAM11(fabric_sram1_a_din_o[11]),
        .Tile_X11Y12_A_DIN_SRAM12(fabric_sram1_a_din_o[12]),
        .Tile_X11Y12_A_DIN_SRAM13(fabric_sram1_a_din_o[13]),
        .Tile_X11Y12_A_DIN_SRAM14(fabric_sram1_a_din_o[14]),
        .Tile_X11Y12_A_DIN_SRAM15(fabric_sram1_a_din_o[15]),
        .Tile_X11Y12_A_DIN_SRAM16(fabric_sram1_a_din_o[16]),
        .Tile_X11Y12_A_DIN_SRAM17(fabric_sram1_a_din_o[17]),
        .Tile_X11Y12_A_DIN_SRAM18(fabric_sram1_a_din_o[18]),
        .Tile_X11Y12_A_DIN_SRAM19(fabric_sram1_a_din_o[19]),
        .Tile_X11Y12_A_DIN_SRAM20(fabric_sram1_a_din_o[20]),
        .Tile_X11Y12_A_DIN_SRAM21(fabric_sram1_a_din_o[21]),
        .Tile_X11Y12_A_DIN_SRAM22(fabric_sram1_a_din_o[22]),
        .Tile_X11Y12_A_DIN_SRAM23(fabric_sram1_a_din_o[23]),
        .Tile_X11Y12_A_DIN_SRAM24(fabric_sram1_a_din_o[24]),
        .Tile_X11Y12_A_DIN_SRAM25(fabric_sram1_a_din_o[25]),
        .Tile_X11Y12_A_DIN_SRAM26(fabric_sram1_a_din_o[26]),
        .Tile_X11Y12_A_DIN_SRAM27(fabric_sram1_a_din_o[27]),
        .Tile_X11Y12_A_DIN_SRAM28(fabric_sram1_a_din_o[28]),
        .Tile_X11Y12_A_DIN_SRAM29(fabric_sram1_a_din_o[29]),
        .Tile_X11Y12_A_DIN_SRAM30(fabric_sram1_a_din_o[30]),
        .Tile_X11Y12_A_DIN_SRAM31(fabric_sram1_a_din_o[31]),
        .Tile_X11Y12_A_WEN_SRAM(fabric_sram1_a_wen_o),
        .Tile_X11Y12_A_MEN_SRAM(fabric_sram1_a_men_o),
        .Tile_X11Y12_A_REN_SRAM(fabric_sram1_a_ren_o),
        .Tile_X11Y12_A_CLK_SRAM(fabric_sram1_a_clk_o),
        .Tile_X11Y12_A_TIE_HIGH_SRAM(fabric_sram1_a_tie_high_o),
        .Tile_X11Y12_A_TIE_LOW_SRAM(fabric_sram1_a_tie_low_o),
        .Tile_X11Y12_CONFIGURED_top(configured_i),

        // SRAM 2
        .Tile_X11Y14_A_DOUT_SRAM0(fabric_sram2_a_dout_i[0]),
        .Tile_X11Y14_A_DOUT_SRAM1(fabric_sram2_a_dout_i[1]),
        .Tile_X11Y14_A_DOUT_SRAM2(fabric_sram2_a_dout_i[2]),
        .Tile_X11Y14_A_DOUT_SRAM3(fabric_sram2_a_dout_i[3]),
        .Tile_X11Y14_A_DOUT_SRAM4(fabric_sram2_a_dout_i[4]),
        .Tile_X11Y14_A_DOUT_SRAM5(fabric_sram2_a_dout_i[5]),
        .Tile_X11Y14_A_DOUT_SRAM6(fabric_sram2_a_dout_i[6]),
        .Tile_X11Y14_A_DOUT_SRAM7(fabric_sram2_a_dout_i[7]),
        .Tile_X11Y14_A_DOUT_SRAM8(fabric_sram2_a_dout_i[8]),
        .Tile_X11Y14_A_DOUT_SRAM9(fabric_sram2_a_dout_i[9]),
        .Tile_X11Y14_A_DOUT_SRAM10(fabric_sram2_a_dout_i[10]),
        .Tile_X11Y14_A_DOUT_SRAM11(fabric_sram2_a_dout_i[11]),
        .Tile_X11Y14_A_DOUT_SRAM12(fabric_sram2_a_dout_i[12]),
        .Tile_X11Y14_A_DOUT_SRAM13(fabric_sram2_a_dout_i[13]),
        .Tile_X11Y14_A_DOUT_SRAM14(fabric_sram2_a_dout_i[14]),
        .Tile_X11Y14_A_DOUT_SRAM15(fabric_sram2_a_dout_i[15]),
        .Tile_X11Y14_A_DOUT_SRAM16(fabric_sram2_a_dout_i[16]),
        .Tile_X11Y14_A_DOUT_SRAM17(fabric_sram2_a_dout_i[17]),
        .Tile_X11Y14_A_DOUT_SRAM18(fabric_sram2_a_dout_i[18]),
        .Tile_X11Y14_A_DOUT_SRAM19(fabric_sram2_a_dout_i[19]),
        .Tile_X11Y14_A_DOUT_SRAM20(fabric_sram2_a_dout_i[20]),
        .Tile_X11Y14_A_DOUT_SRAM21(fabric_sram2_a_dout_i[21]),
        .Tile_X11Y14_A_DOUT_SRAM22(fabric_sram2_a_dout_i[22]),
        .Tile_X11Y14_A_DOUT_SRAM23(fabric_sram2_a_dout_i[23]),
        .Tile_X11Y14_A_DOUT_SRAM24(fabric_sram2_a_dout_i[24]),
        .Tile_X11Y14_A_DOUT_SRAM25(fabric_sram2_a_dout_i[25]),
        .Tile_X11Y14_A_DOUT_SRAM26(fabric_sram2_a_dout_i[26]),
        .Tile_X11Y14_A_DOUT_SRAM27(fabric_sram2_a_dout_i[27]),
        .Tile_X11Y14_A_DOUT_SRAM28(fabric_sram2_a_dout_i[28]),
        .Tile_X11Y14_A_DOUT_SRAM29(fabric_sram2_a_dout_i[29]),
        .Tile_X11Y14_A_DOUT_SRAM30(fabric_sram2_a_dout_i[30]),
        .Tile_X11Y14_A_DOUT_SRAM31(fabric_sram2_a_dout_i[31]),
        .Tile_X11Y14_A_ADDR_SRAM0(fabric_sram2_a_addr_o[0]),
        .Tile_X11Y14_A_ADDR_SRAM1(fabric_sram2_a_addr_o[1]),
        .Tile_X11Y14_A_ADDR_SRAM2(fabric_sram2_a_addr_o[2]),
        .Tile_X11Y14_A_ADDR_SRAM3(fabric_sram2_a_addr_o[3]),
        .Tile_X11Y14_A_ADDR_SRAM4(fabric_sram2_a_addr_o[4]),
        .Tile_X11Y14_A_ADDR_SRAM5(fabric_sram2_a_addr_o[5]),
        .Tile_X11Y14_A_ADDR_SRAM6(fabric_sram2_a_addr_o[6]),
        .Tile_X11Y14_A_ADDR_SRAM7(fabric_sram2_a_addr_o[7]),
        .Tile_X11Y14_A_ADDR_SRAM8(fabric_sram2_a_addr_o[8]),
        .Tile_X11Y14_A_ADDR_SRAM9(fabric_sram2_a_addr_o[9]),
        .Tile_X11Y14_A_BM_SRAM0(fabric_sram2_a_bm_o[0]),
        .Tile_X11Y14_A_BM_SRAM1(fabric_sram2_a_bm_o[1]),
        .Tile_X11Y14_A_BM_SRAM2(fabric_sram2_a_bm_o[2]),
        .Tile_X11Y14_A_BM_SRAM3(fabric_sram2_a_bm_o[3]),
        .Tile_X11Y14_A_BM_SRAM4(fabric_sram2_a_bm_o[4]),
        .Tile_X11Y14_A_BM_SRAM5(fabric_sram2_a_bm_o[5]),
        .Tile_X11Y14_A_BM_SRAM6(fabric_sram2_a_bm_o[6]),
        .Tile_X11Y14_A_BM_SRAM7(fabric_sram2_a_bm_o[7]),
        .Tile_X11Y14_A_BM_SRAM8(fabric_sram2_a_bm_o[8]),
        .Tile_X11Y14_A_BM_SRAM9(fabric_sram2_a_bm_o[9]),
        .Tile_X11Y14_A_BM_SRAM10(fabric_sram2_a_bm_o[10]),
        .Tile_X11Y14_A_BM_SRAM11(fabric_sram2_a_bm_o[11]),
        .Tile_X11Y14_A_BM_SRAM12(fabric_sram2_a_bm_o[12]),
        .Tile_X11Y14_A_BM_SRAM13(fabric_sram2_a_bm_o[13]),
        .Tile_X11Y14_A_BM_SRAM14(fabric_sram2_a_bm_o[14]),
        .Tile_X11Y14_A_BM_SRAM15(fabric_sram2_a_bm_o[15]),
        .Tile_X11Y14_A_BM_SRAM16(fabric_sram2_a_bm_o[16]),
        .Tile_X11Y14_A_BM_SRAM17(fabric_sram2_a_bm_o[17]),
        .Tile_X11Y14_A_BM_SRAM18(fabric_sram2_a_bm_o[18]),
        .Tile_X11Y14_A_BM_SRAM19(fabric_sram2_a_bm_o[19]),
        .Tile_X11Y14_A_BM_SRAM20(fabric_sram2_a_bm_o[20]),
        .Tile_X11Y14_A_BM_SRAM21(fabric_sram2_a_bm_o[21]),
        .Tile_X11Y14_A_BM_SRAM22(fabric_sram2_a_bm_o[22]),
        .Tile_X11Y14_A_BM_SRAM23(fabric_sram2_a_bm_o[23]),
        .Tile_X11Y14_A_BM_SRAM24(fabric_sram2_a_bm_o[24]),
        .Tile_X11Y14_A_BM_SRAM25(fabric_sram2_a_bm_o[25]),
        .Tile_X11Y14_A_BM_SRAM26(fabric_sram2_a_bm_o[26]),
        .Tile_X11Y14_A_BM_SRAM27(fabric_sram2_a_bm_o[27]),
        .Tile_X11Y14_A_BM_SRAM28(fabric_sram2_a_bm_o[28]),
        .Tile_X11Y14_A_BM_SRAM29(fabric_sram2_a_bm_o[29]),
        .Tile_X11Y14_A_BM_SRAM30(fabric_sram2_a_bm_o[30]),
        .Tile_X11Y14_A_BM_SRAM31(fabric_sram2_a_bm_o[31]),
        .Tile_X11Y14_A_DIN_SRAM0(fabric_sram2_a_din_o[0]),
        .Tile_X11Y14_A_DIN_SRAM1(fabric_sram2_a_din_o[1]),
        .Tile_X11Y14_A_DIN_SRAM2(fabric_sram2_a_din_o[2]),
        .Tile_X11Y14_A_DIN_SRAM3(fabric_sram2_a_din_o[3]),
        .Tile_X11Y14_A_DIN_SRAM4(fabric_sram2_a_din_o[4]),
        .Tile_X11Y14_A_DIN_SRAM5(fabric_sram2_a_din_o[5]),
        .Tile_X11Y14_A_DIN_SRAM6(fabric_sram2_a_din_o[6]),
        .Tile_X11Y14_A_DIN_SRAM7(fabric_sram2_a_din_o[7]),
        .Tile_X11Y14_A_DIN_SRAM8(fabric_sram2_a_din_o[8]),
        .Tile_X11Y14_A_DIN_SRAM9(fabric_sram2_a_din_o[9]),
        .Tile_X11Y14_A_DIN_SRAM10(fabric_sram2_a_din_o[10]),
        .Tile_X11Y14_A_DIN_SRAM11(fabric_sram2_a_din_o[11]),
        .Tile_X11Y14_A_DIN_SRAM12(fabric_sram2_a_din_o[12]),
        .Tile_X11Y14_A_DIN_SRAM13(fabric_sram2_a_din_o[13]),
        .Tile_X11Y14_A_DIN_SRAM14(fabric_sram2_a_din_o[14]),
        .Tile_X11Y14_A_DIN_SRAM15(fabric_sram2_a_din_o[15]),
        .Tile_X11Y14_A_DIN_SRAM16(fabric_sram2_a_din_o[16]),
        .Tile_X11Y14_A_DIN_SRAM17(fabric_sram2_a_din_o[17]),
        .Tile_X11Y14_A_DIN_SRAM18(fabric_sram2_a_din_o[18]),
        .Tile_X11Y14_A_DIN_SRAM19(fabric_sram2_a_din_o[19]),
        .Tile_X11Y14_A_DIN_SRAM20(fabric_sram2_a_din_o[20]),
        .Tile_X11Y14_A_DIN_SRAM21(fabric_sram2_a_din_o[21]),
        .Tile_X11Y14_A_DIN_SRAM22(fabric_sram2_a_din_o[22]),
        .Tile_X11Y14_A_DIN_SRAM23(fabric_sram2_a_din_o[23]),
        .Tile_X11Y14_A_DIN_SRAM24(fabric_sram2_a_din_o[24]),
        .Tile_X11Y14_A_DIN_SRAM25(fabric_sram2_a_din_o[25]),
        .Tile_X11Y14_A_DIN_SRAM26(fabric_sram2_a_din_o[26]),
        .Tile_X11Y14_A_DIN_SRAM27(fabric_sram2_a_din_o[27]),
        .Tile_X11Y14_A_DIN_SRAM28(fabric_sram2_a_din_o[28]),
        .Tile_X11Y14_A_DIN_SRAM29(fabric_sram2_a_din_o[29]),
        .Tile_X11Y14_A_DIN_SRAM30(fabric_sram2_a_din_o[30]),
        .Tile_X11Y14_A_DIN_SRAM31(fabric_sram2_a_din_o[31]),
        .Tile_X11Y14_A_WEN_SRAM(fabric_sram2_a_wen_o),
        .Tile_X11Y14_A_MEN_SRAM(fabric_sram2_a_men_o),
        .Tile_X11Y14_A_REN_SRAM(fabric_sram2_a_ren_o),
        .Tile_X11Y14_A_CLK_SRAM(fabric_sram2_a_clk_o),
        .Tile_X11Y14_A_TIE_HIGH_SRAM(fabric_sram2_a_tie_high_o),
        .Tile_X11Y14_A_TIE_LOW_SRAM(fabric_sram2_a_tie_low_o),
        .Tile_X11Y14_CONFIGURED_top(configured_i),

        // SRAM 3
        .Tile_X11Y16_A_DOUT_SRAM0(fabric_sram3_a_dout_i[0]),
        .Tile_X11Y16_A_DOUT_SRAM1(fabric_sram3_a_dout_i[1]),
        .Tile_X11Y16_A_DOUT_SRAM2(fabric_sram3_a_dout_i[2]),
        .Tile_X11Y16_A_DOUT_SRAM3(fabric_sram3_a_dout_i[3]),
        .Tile_X11Y16_A_DOUT_SRAM4(fabric_sram3_a_dout_i[4]),
        .Tile_X11Y16_A_DOUT_SRAM5(fabric_sram3_a_dout_i[5]),
        .Tile_X11Y16_A_DOUT_SRAM6(fabric_sram3_a_dout_i[6]),
        .Tile_X11Y16_A_DOUT_SRAM7(fabric_sram3_a_dout_i[7]),
        .Tile_X11Y16_A_DOUT_SRAM8(fabric_sram3_a_dout_i[8]),
        .Tile_X11Y16_A_DOUT_SRAM9(fabric_sram3_a_dout_i[9]),
        .Tile_X11Y16_A_DOUT_SRAM10(fabric_sram3_a_dout_i[10]),
        .Tile_X11Y16_A_DOUT_SRAM11(fabric_sram3_a_dout_i[11]),
        .Tile_X11Y16_A_DOUT_SRAM12(fabric_sram3_a_dout_i[12]),
        .Tile_X11Y16_A_DOUT_SRAM13(fabric_sram3_a_dout_i[13]),
        .Tile_X11Y16_A_DOUT_SRAM14(fabric_sram3_a_dout_i[14]),
        .Tile_X11Y16_A_DOUT_SRAM15(fabric_sram3_a_dout_i[15]),
        .Tile_X11Y16_A_DOUT_SRAM16(fabric_sram3_a_dout_i[16]),
        .Tile_X11Y16_A_DOUT_SRAM17(fabric_sram3_a_dout_i[17]),
        .Tile_X11Y16_A_DOUT_SRAM18(fabric_sram3_a_dout_i[18]),
        .Tile_X11Y16_A_DOUT_SRAM19(fabric_sram3_a_dout_i[19]),
        .Tile_X11Y16_A_DOUT_SRAM20(fabric_sram3_a_dout_i[20]),
        .Tile_X11Y16_A_DOUT_SRAM21(fabric_sram3_a_dout_i[21]),
        .Tile_X11Y16_A_DOUT_SRAM22(fabric_sram3_a_dout_i[22]),
        .Tile_X11Y16_A_DOUT_SRAM23(fabric_sram3_a_dout_i[23]),
        .Tile_X11Y16_A_DOUT_SRAM24(fabric_sram3_a_dout_i[24]),
        .Tile_X11Y16_A_DOUT_SRAM25(fabric_sram3_a_dout_i[25]),
        .Tile_X11Y16_A_DOUT_SRAM26(fabric_sram3_a_dout_i[26]),
        .Tile_X11Y16_A_DOUT_SRAM27(fabric_sram3_a_dout_i[27]),
        .Tile_X11Y16_A_DOUT_SRAM28(fabric_sram3_a_dout_i[28]),
        .Tile_X11Y16_A_DOUT_SRAM29(fabric_sram3_a_dout_i[29]),
        .Tile_X11Y16_A_DOUT_SRAM30(fabric_sram3_a_dout_i[30]),
        .Tile_X11Y16_A_DOUT_SRAM31(fabric_sram3_a_dout_i[31]),
        .Tile_X11Y16_A_ADDR_SRAM0(fabric_sram3_a_addr_o[0]),
        .Tile_X11Y16_A_ADDR_SRAM1(fabric_sram3_a_addr_o[1]),
        .Tile_X11Y16_A_ADDR_SRAM2(fabric_sram3_a_addr_o[2]),
        .Tile_X11Y16_A_ADDR_SRAM3(fabric_sram3_a_addr_o[3]),
        .Tile_X11Y16_A_ADDR_SRAM4(fabric_sram3_a_addr_o[4]),
        .Tile_X11Y16_A_ADDR_SRAM5(fabric_sram3_a_addr_o[5]),
        .Tile_X11Y16_A_ADDR_SRAM6(fabric_sram3_a_addr_o[6]),
        .Tile_X11Y16_A_ADDR_SRAM7(fabric_sram3_a_addr_o[7]),
        .Tile_X11Y16_A_ADDR_SRAM8(fabric_sram3_a_addr_o[8]),
        .Tile_X11Y16_A_ADDR_SRAM9(fabric_sram3_a_addr_o[9]),
        .Tile_X11Y16_A_BM_SRAM0(fabric_sram3_a_bm_o[0]),
        .Tile_X11Y16_A_BM_SRAM1(fabric_sram3_a_bm_o[1]),
        .Tile_X11Y16_A_BM_SRAM2(fabric_sram3_a_bm_o[2]),
        .Tile_X11Y16_A_BM_SRAM3(fabric_sram3_a_bm_o[3]),
        .Tile_X11Y16_A_BM_SRAM4(fabric_sram3_a_bm_o[4]),
        .Tile_X11Y16_A_BM_SRAM5(fabric_sram3_a_bm_o[5]),
        .Tile_X11Y16_A_BM_SRAM6(fabric_sram3_a_bm_o[6]),
        .Tile_X11Y16_A_BM_SRAM7(fabric_sram3_a_bm_o[7]),
        .Tile_X11Y16_A_BM_SRAM8(fabric_sram3_a_bm_o[8]),
        .Tile_X11Y16_A_BM_SRAM9(fabric_sram3_a_bm_o[9]),
        .Tile_X11Y16_A_BM_SRAM10(fabric_sram3_a_bm_o[10]),
        .Tile_X11Y16_A_BM_SRAM11(fabric_sram3_a_bm_o[11]),
        .Tile_X11Y16_A_BM_SRAM12(fabric_sram3_a_bm_o[12]),
        .Tile_X11Y16_A_BM_SRAM13(fabric_sram3_a_bm_o[13]),
        .Tile_X11Y16_A_BM_SRAM14(fabric_sram3_a_bm_o[14]),
        .Tile_X11Y16_A_BM_SRAM15(fabric_sram3_a_bm_o[15]),
        .Tile_X11Y16_A_BM_SRAM16(fabric_sram3_a_bm_o[16]),
        .Tile_X11Y16_A_BM_SRAM17(fabric_sram3_a_bm_o[17]),
        .Tile_X11Y16_A_BM_SRAM18(fabric_sram3_a_bm_o[18]),
        .Tile_X11Y16_A_BM_SRAM19(fabric_sram3_a_bm_o[19]),
        .Tile_X11Y16_A_BM_SRAM20(fabric_sram3_a_bm_o[20]),
        .Tile_X11Y16_A_BM_SRAM21(fabric_sram3_a_bm_o[21]),
        .Tile_X11Y16_A_BM_SRAM22(fabric_sram3_a_bm_o[22]),
        .Tile_X11Y16_A_BM_SRAM23(fabric_sram3_a_bm_o[23]),
        .Tile_X11Y16_A_BM_SRAM24(fabric_sram3_a_bm_o[24]),
        .Tile_X11Y16_A_BM_SRAM25(fabric_sram3_a_bm_o[25]),
        .Tile_X11Y16_A_BM_SRAM26(fabric_sram3_a_bm_o[26]),
        .Tile_X11Y16_A_BM_SRAM27(fabric_sram3_a_bm_o[27]),
        .Tile_X11Y16_A_BM_SRAM28(fabric_sram3_a_bm_o[28]),
        .Tile_X11Y16_A_BM_SRAM29(fabric_sram3_a_bm_o[29]),
        .Tile_X11Y16_A_BM_SRAM30(fabric_sram3_a_bm_o[30]),
        .Tile_X11Y16_A_BM_SRAM31(fabric_sram3_a_bm_o[31]),
        .Tile_X11Y16_A_DIN_SRAM0(fabric_sram3_a_din_o[0]),
        .Tile_X11Y16_A_DIN_SRAM1(fabric_sram3_a_din_o[1]),
        .Tile_X11Y16_A_DIN_SRAM2(fabric_sram3_a_din_o[2]),
        .Tile_X11Y16_A_DIN_SRAM3(fabric_sram3_a_din_o[3]),
        .Tile_X11Y16_A_DIN_SRAM4(fabric_sram3_a_din_o[4]),
        .Tile_X11Y16_A_DIN_SRAM5(fabric_sram3_a_din_o[5]),
        .Tile_X11Y16_A_DIN_SRAM6(fabric_sram3_a_din_o[6]),
        .Tile_X11Y16_A_DIN_SRAM7(fabric_sram3_a_din_o[7]),
        .Tile_X11Y16_A_DIN_SRAM8(fabric_sram3_a_din_o[8]),
        .Tile_X11Y16_A_DIN_SRAM9(fabric_sram3_a_din_o[9]),
        .Tile_X11Y16_A_DIN_SRAM10(fabric_sram3_a_din_o[10]),
        .Tile_X11Y16_A_DIN_SRAM11(fabric_sram3_a_din_o[11]),
        .Tile_X11Y16_A_DIN_SRAM12(fabric_sram3_a_din_o[12]),
        .Tile_X11Y16_A_DIN_SRAM13(fabric_sram3_a_din_o[13]),
        .Tile_X11Y16_A_DIN_SRAM14(fabric_sram3_a_din_o[14]),
        .Tile_X11Y16_A_DIN_SRAM15(fabric_sram3_a_din_o[15]),
        .Tile_X11Y16_A_DIN_SRAM16(fabric_sram3_a_din_o[16]),
        .Tile_X11Y16_A_DIN_SRAM17(fabric_sram3_a_din_o[17]),
        .Tile_X11Y16_A_DIN_SRAM18(fabric_sram3_a_din_o[18]),
        .Tile_X11Y16_A_DIN_SRAM19(fabric_sram3_a_din_o[19]),
        .Tile_X11Y16_A_DIN_SRAM20(fabric_sram3_a_din_o[20]),
        .Tile_X11Y16_A_DIN_SRAM21(fabric_sram3_a_din_o[21]),
        .Tile_X11Y16_A_DIN_SRAM22(fabric_sram3_a_din_o[22]),
        .Tile_X11Y16_A_DIN_SRAM23(fabric_sram3_a_din_o[23]),
        .Tile_X11Y16_A_DIN_SRAM24(fabric_sram3_a_din_o[24]),
        .Tile_X11Y16_A_DIN_SRAM25(fabric_sram3_a_din_o[25]),
        .Tile_X11Y16_A_DIN_SRAM26(fabric_sram3_a_din_o[26]),
        .Tile_X11Y16_A_DIN_SRAM27(fabric_sram3_a_din_o[27]),
        .Tile_X11Y16_A_DIN_SRAM28(fabric_sram3_a_din_o[28]),
        .Tile_X11Y16_A_DIN_SRAM29(fabric_sram3_a_din_o[29]),
        .Tile_X11Y16_A_DIN_SRAM30(fabric_sram3_a_din_o[30]),
        .Tile_X11Y16_A_DIN_SRAM31(fabric_sram3_a_din_o[31]),
        .Tile_X11Y16_A_WEN_SRAM(fabric_sram3_a_wen_o),
        .Tile_X11Y16_A_MEN_SRAM(fabric_sram3_a_men_o),
        .Tile_X11Y16_A_REN_SRAM(fabric_sram3_a_ren_o),
        .Tile_X11Y16_A_CLK_SRAM(fabric_sram3_a_clk_o),
        .Tile_X11Y16_A_TIE_HIGH_SRAM(fabric_sram3_a_tie_high_o),
        .Tile_X11Y16_A_TIE_LOW_SRAM(fabric_sram3_a_tie_low_o),
        .Tile_X11Y16_CONFIGURED_top(configured_i),

        // BRAM 0
        // Port A
        .Tile_X11Y2_A_DOUT_BRAM0(fabric_bram0_a_dout_i[0]),
        .Tile_X11Y2_A_DOUT_BRAM1(fabric_bram0_a_dout_i[1]),
        .Tile_X11Y2_A_DOUT_BRAM2(fabric_bram0_a_dout_i[2]),
        .Tile_X11Y2_A_DOUT_BRAM3(fabric_bram0_a_dout_i[3]),
        .Tile_X11Y2_A_DOUT_BRAM4(fabric_bram0_a_dout_i[4]),
        .Tile_X11Y2_A_DOUT_BRAM5(fabric_bram0_a_dout_i[5]),
        .Tile_X11Y2_A_DOUT_BRAM6(fabric_bram0_a_dout_i[6]),
        .Tile_X11Y2_A_DOUT_BRAM7(fabric_bram0_a_dout_i[7]),
        .Tile_X11Y2_A_DOUT_BRAM8(fabric_bram0_a_dout_i[8]),
        .Tile_X11Y2_A_DOUT_BRAM9(fabric_bram0_a_dout_i[9]),
        .Tile_X11Y2_A_DOUT_BRAM10(fabric_bram0_a_dout_i[10]),
        .Tile_X11Y2_A_DOUT_BRAM11(fabric_bram0_a_dout_i[11]),
        .Tile_X11Y2_A_DOUT_BRAM12(fabric_bram0_a_dout_i[12]),
        .Tile_X11Y2_A_DOUT_BRAM13(fabric_bram0_a_dout_i[13]),
        .Tile_X11Y2_A_DOUT_BRAM14(fabric_bram0_a_dout_i[14]),
        .Tile_X11Y2_A_DOUT_BRAM15(fabric_bram0_a_dout_i[15]),
        .Tile_X11Y2_A_ADDR_BRAM0(fabric_bram0_a_addr_o[0]),
        .Tile_X11Y2_A_ADDR_BRAM1(fabric_bram0_a_addr_o[1]),
        .Tile_X11Y2_A_ADDR_BRAM2(fabric_bram0_a_addr_o[2]),
        .Tile_X11Y2_A_ADDR_BRAM3(fabric_bram0_a_addr_o[3]),
        .Tile_X11Y2_A_ADDR_BRAM4(fabric_bram0_a_addr_o[4]),
        .Tile_X11Y2_A_ADDR_BRAM5(fabric_bram0_a_addr_o[5]),
        .Tile_X11Y2_A_ADDR_BRAM6(fabric_bram0_a_addr_o[6]),
        .Tile_X11Y2_A_ADDR_BRAM7(fabric_bram0_a_addr_o[7]),
        .Tile_X11Y2_A_ADDR_BRAM8(fabric_bram0_a_addr_o[8]),
        .Tile_X11Y2_A_ADDR_BRAM9(fabric_bram0_a_addr_o[9]),
        .Tile_X11Y2_A_BM_BRAM0(fabric_bram0_a_bm_o[0]),
        .Tile_X11Y2_A_BM_BRAM1(fabric_bram0_a_bm_o[1]),
        .Tile_X11Y2_A_BM_BRAM2(fabric_bram0_a_bm_o[2]),
        .Tile_X11Y2_A_BM_BRAM3(fabric_bram0_a_bm_o[3]),
        .Tile_X11Y2_A_BM_BRAM4(fabric_bram0_a_bm_o[4]),
        .Tile_X11Y2_A_BM_BRAM5(fabric_bram0_a_bm_o[5]),
        .Tile_X11Y2_A_BM_BRAM6(fabric_bram0_a_bm_o[6]),
        .Tile_X11Y2_A_BM_BRAM7(fabric_bram0_a_bm_o[7]),
        .Tile_X11Y2_A_BM_BRAM8(fabric_bram0_a_bm_o[8]),
        .Tile_X11Y2_A_BM_BRAM9(fabric_bram0_a_bm_o[9]),
        .Tile_X11Y2_A_BM_BRAM10(fabric_bram0_a_bm_o[10]),
        .Tile_X11Y2_A_BM_BRAM11(fabric_bram0_a_bm_o[11]),
        .Tile_X11Y2_A_BM_BRAM12(fabric_bram0_a_bm_o[12]),
        .Tile_X11Y2_A_BM_BRAM13(fabric_bram0_a_bm_o[13]),
        .Tile_X11Y2_A_BM_BRAM14(fabric_bram0_a_bm_o[14]),
        .Tile_X11Y2_A_BM_BRAM15(fabric_bram0_a_bm_o[15]),
        .Tile_X11Y2_A_DIN_BRAM0(fabric_bram0_a_din_o[0]),
        .Tile_X11Y2_A_DIN_BRAM1(fabric_bram0_a_din_o[1]),
        .Tile_X11Y2_A_DIN_BRAM2(fabric_bram0_a_din_o[2]),
        .Tile_X11Y2_A_DIN_BRAM3(fabric_bram0_a_din_o[3]),
        .Tile_X11Y2_A_DIN_BRAM4(fabric_bram0_a_din_o[4]),
        .Tile_X11Y2_A_DIN_BRAM5(fabric_bram0_a_din_o[5]),
        .Tile_X11Y2_A_DIN_BRAM6(fabric_bram0_a_din_o[6]),
        .Tile_X11Y2_A_DIN_BRAM7(fabric_bram0_a_din_o[7]),
        .Tile_X11Y2_A_DIN_BRAM8(fabric_bram0_a_din_o[8]),
        .Tile_X11Y2_A_DIN_BRAM9(fabric_bram0_a_din_o[9]),
        .Tile_X11Y2_A_DIN_BRAM10(fabric_bram0_a_din_o[10]),
        .Tile_X11Y2_A_DIN_BRAM11(fabric_bram0_a_din_o[11]),
        .Tile_X11Y2_A_DIN_BRAM12(fabric_bram0_a_din_o[12]),
        .Tile_X11Y2_A_DIN_BRAM13(fabric_bram0_a_din_o[13]),
        .Tile_X11Y2_A_DIN_BRAM14(fabric_bram0_a_din_o[14]),
        .Tile_X11Y2_A_DIN_BRAM15(fabric_bram0_a_din_o[15]),
        .Tile_X11Y2_A_WEN_BRAM(fabric_bram0_a_wen_o),
        .Tile_X11Y2_A_MEN_BRAM(fabric_bram0_a_men_o),
        .Tile_X11Y2_A_REN_BRAM(fabric_bram0_a_ren_o),
        .Tile_X11Y2_A_CLK_BRAM(fabric_bram0_a_clk_o),
        .Tile_X11Y2_A_TIE_HIGH_BRAM(fabric_bram0_a_tie_high_o),
        .Tile_X11Y2_A_TIE_LOW_BRAM(fabric_bram0_a_tie_low_o),

        // Port B
        .Tile_X11Y2_B_DOUT_BRAM0(fabric_bram0_b_dout_i[0]),
        .Tile_X11Y2_B_DOUT_BRAM1(fabric_bram0_b_dout_i[1]),
        .Tile_X11Y2_B_DOUT_BRAM2(fabric_bram0_b_dout_i[2]),
        .Tile_X11Y2_B_DOUT_BRAM3(fabric_bram0_b_dout_i[3]),
        .Tile_X11Y2_B_DOUT_BRAM4(fabric_bram0_b_dout_i[4]),
        .Tile_X11Y2_B_DOUT_BRAM5(fabric_bram0_b_dout_i[5]),
        .Tile_X11Y2_B_DOUT_BRAM6(fabric_bram0_b_dout_i[6]),
        .Tile_X11Y2_B_DOUT_BRAM7(fabric_bram0_b_dout_i[7]),
        .Tile_X11Y2_B_DOUT_BRAM8(fabric_bram0_b_dout_i[8]),
        .Tile_X11Y2_B_DOUT_BRAM9(fabric_bram0_b_dout_i[9]),
        .Tile_X11Y2_B_DOUT_BRAM10(fabric_bram0_b_dout_i[10]),
        .Tile_X11Y2_B_DOUT_BRAM11(fabric_bram0_b_dout_i[11]),
        .Tile_X11Y2_B_DOUT_BRAM12(fabric_bram0_b_dout_i[12]),
        .Tile_X11Y2_B_DOUT_BRAM13(fabric_bram0_b_dout_i[13]),
        .Tile_X11Y2_B_DOUT_BRAM14(fabric_bram0_b_dout_i[14]),
        .Tile_X11Y2_B_DOUT_BRAM15(fabric_bram0_b_dout_i[15]),
        .Tile_X11Y2_B_ADDR_BRAM0(fabric_bram0_b_addr_o[0]),
        .Tile_X11Y2_B_ADDR_BRAM1(fabric_bram0_b_addr_o[1]),
        .Tile_X11Y2_B_ADDR_BRAM2(fabric_bram0_b_addr_o[2]),
        .Tile_X11Y2_B_ADDR_BRAM3(fabric_bram0_b_addr_o[3]),
        .Tile_X11Y2_B_ADDR_BRAM4(fabric_bram0_b_addr_o[4]),
        .Tile_X11Y2_B_ADDR_BRAM5(fabric_bram0_b_addr_o[5]),
        .Tile_X11Y2_B_ADDR_BRAM6(fabric_bram0_b_addr_o[6]),
        .Tile_X11Y2_B_ADDR_BRAM7(fabric_bram0_b_addr_o[7]),
        .Tile_X11Y2_B_ADDR_BRAM8(fabric_bram0_b_addr_o[8]),
        .Tile_X11Y2_B_ADDR_BRAM9(fabric_bram0_b_addr_o[9]),
        .Tile_X11Y2_B_BM_BRAM0(fabric_bram0_b_bm_o[0]),
        .Tile_X11Y2_B_BM_BRAM1(fabric_bram0_b_bm_o[1]),
        .Tile_X11Y2_B_BM_BRAM2(fabric_bram0_b_bm_o[2]),
        .Tile_X11Y2_B_BM_BRAM3(fabric_bram0_b_bm_o[3]),
        .Tile_X11Y2_B_BM_BRAM4(fabric_bram0_b_bm_o[4]),
        .Tile_X11Y2_B_BM_BRAM5(fabric_bram0_b_bm_o[5]),
        .Tile_X11Y2_B_BM_BRAM6(fabric_bram0_b_bm_o[6]),
        .Tile_X11Y2_B_BM_BRAM7(fabric_bram0_b_bm_o[7]),
        .Tile_X11Y2_B_BM_BRAM8(fabric_bram0_b_bm_o[8]),
        .Tile_X11Y2_B_BM_BRAM9(fabric_bram0_b_bm_o[9]),
        .Tile_X11Y2_B_BM_BRAM10(fabric_bram0_b_bm_o[10]),
        .Tile_X11Y2_B_BM_BRAM11(fabric_bram0_b_bm_o[11]),
        .Tile_X11Y2_B_BM_BRAM12(fabric_bram0_b_bm_o[12]),
        .Tile_X11Y2_B_BM_BRAM13(fabric_bram0_b_bm_o[13]),
        .Tile_X11Y2_B_BM_BRAM14(fabric_bram0_b_bm_o[14]),
        .Tile_X11Y2_B_BM_BRAM15(fabric_bram0_b_bm_o[15]),
        .Tile_X11Y2_B_DIN_BRAM0(fabric_bram0_b_din_o[0]),
        .Tile_X11Y2_B_DIN_BRAM1(fabric_bram0_b_din_o[1]),
        .Tile_X11Y2_B_DIN_BRAM2(fabric_bram0_b_din_o[2]),
        .Tile_X11Y2_B_DIN_BRAM3(fabric_bram0_b_din_o[3]),
        .Tile_X11Y2_B_DIN_BRAM4(fabric_bram0_b_din_o[4]),
        .Tile_X11Y2_B_DIN_BRAM5(fabric_bram0_b_din_o[5]),
        .Tile_X11Y2_B_DIN_BRAM6(fabric_bram0_b_din_o[6]),
        .Tile_X11Y2_B_DIN_BRAM7(fabric_bram0_b_din_o[7]),
        .Tile_X11Y2_B_DIN_BRAM8(fabric_bram0_b_din_o[8]),
        .Tile_X11Y2_B_DIN_BRAM9(fabric_bram0_b_din_o[9]),
        .Tile_X11Y2_B_DIN_BRAM10(fabric_bram0_b_din_o[10]),
        .Tile_X11Y2_B_DIN_BRAM11(fabric_bram0_b_din_o[11]),
        .Tile_X11Y2_B_DIN_BRAM12(fabric_bram0_b_din_o[12]),
        .Tile_X11Y2_B_DIN_BRAM13(fabric_bram0_b_din_o[13]),
        .Tile_X11Y2_B_DIN_BRAM14(fabric_bram0_b_din_o[14]),
        .Tile_X11Y2_B_DIN_BRAM15(fabric_bram0_b_din_o[15]),
        .Tile_X11Y2_B_WEN_BRAM(fabric_bram0_b_wen_o),
        .Tile_X11Y2_B_MEN_BRAM(fabric_bram0_b_men_o),
        .Tile_X11Y2_B_REN_BRAM(fabric_bram0_b_ren_o),
        .Tile_X11Y2_B_CLK_BRAM(fabric_bram0_b_clk_o),
        .Tile_X11Y2_B_TIE_HIGH_BRAM(fabric_bram0_b_tie_high_o),
        .Tile_X11Y2_B_TIE_LOW_BRAM(fabric_bram0_b_tie_low_o),

        .Tile_X11Y2_CONFIGURED_top(configured_i),

        // BRAM 1
        // Port A
        .Tile_X11Y4_A_DOUT_BRAM0(fabric_bram1_a_dout_i[0]),
        .Tile_X11Y4_A_DOUT_BRAM1(fabric_bram1_a_dout_i[1]),
        .Tile_X11Y4_A_DOUT_BRAM2(fabric_bram1_a_dout_i[2]),
        .Tile_X11Y4_A_DOUT_BRAM3(fabric_bram1_a_dout_i[3]),
        .Tile_X11Y4_A_DOUT_BRAM4(fabric_bram1_a_dout_i[4]),
        .Tile_X11Y4_A_DOUT_BRAM5(fabric_bram1_a_dout_i[5]),
        .Tile_X11Y4_A_DOUT_BRAM6(fabric_bram1_a_dout_i[6]),
        .Tile_X11Y4_A_DOUT_BRAM7(fabric_bram1_a_dout_i[7]),
        .Tile_X11Y4_A_DOUT_BRAM8(fabric_bram1_a_dout_i[8]),
        .Tile_X11Y4_A_DOUT_BRAM9(fabric_bram1_a_dout_i[9]),
        .Tile_X11Y4_A_DOUT_BRAM10(fabric_bram1_a_dout_i[10]),
        .Tile_X11Y4_A_DOUT_BRAM11(fabric_bram1_a_dout_i[11]),
        .Tile_X11Y4_A_DOUT_BRAM12(fabric_bram1_a_dout_i[12]),
        .Tile_X11Y4_A_DOUT_BRAM13(fabric_bram1_a_dout_i[13]),
        .Tile_X11Y4_A_DOUT_BRAM14(fabric_bram1_a_dout_i[14]),
        .Tile_X11Y4_A_DOUT_BRAM15(fabric_bram1_a_dout_i[15]),
        .Tile_X11Y4_A_ADDR_BRAM0(fabric_bram1_a_addr_o[0]),
        .Tile_X11Y4_A_ADDR_BRAM1(fabric_bram1_a_addr_o[1]),
        .Tile_X11Y4_A_ADDR_BRAM2(fabric_bram1_a_addr_o[2]),
        .Tile_X11Y4_A_ADDR_BRAM3(fabric_bram1_a_addr_o[3]),
        .Tile_X11Y4_A_ADDR_BRAM4(fabric_bram1_a_addr_o[4]),
        .Tile_X11Y4_A_ADDR_BRAM5(fabric_bram1_a_addr_o[5]),
        .Tile_X11Y4_A_ADDR_BRAM6(fabric_bram1_a_addr_o[6]),
        .Tile_X11Y4_A_ADDR_BRAM7(fabric_bram1_a_addr_o[7]),
        .Tile_X11Y4_A_ADDR_BRAM8(fabric_bram1_a_addr_o[8]),
        .Tile_X11Y4_A_ADDR_BRAM9(fabric_bram1_a_addr_o[9]),
        .Tile_X11Y4_A_BM_BRAM0(fabric_bram1_a_bm_o[0]),
        .Tile_X11Y4_A_BM_BRAM1(fabric_bram1_a_bm_o[1]),
        .Tile_X11Y4_A_BM_BRAM2(fabric_bram1_a_bm_o[2]),
        .Tile_X11Y4_A_BM_BRAM3(fabric_bram1_a_bm_o[3]),
        .Tile_X11Y4_A_BM_BRAM4(fabric_bram1_a_bm_o[4]),
        .Tile_X11Y4_A_BM_BRAM5(fabric_bram1_a_bm_o[5]),
        .Tile_X11Y4_A_BM_BRAM6(fabric_bram1_a_bm_o[6]),
        .Tile_X11Y4_A_BM_BRAM7(fabric_bram1_a_bm_o[7]),
        .Tile_X11Y4_A_BM_BRAM8(fabric_bram1_a_bm_o[8]),
        .Tile_X11Y4_A_BM_BRAM9(fabric_bram1_a_bm_o[9]),
        .Tile_X11Y4_A_BM_BRAM10(fabric_bram1_a_bm_o[10]),
        .Tile_X11Y4_A_BM_BRAM11(fabric_bram1_a_bm_o[11]),
        .Tile_X11Y4_A_BM_BRAM12(fabric_bram1_a_bm_o[12]),
        .Tile_X11Y4_A_BM_BRAM13(fabric_bram1_a_bm_o[13]),
        .Tile_X11Y4_A_BM_BRAM14(fabric_bram1_a_bm_o[14]),
        .Tile_X11Y4_A_BM_BRAM15(fabric_bram1_a_bm_o[15]),
        .Tile_X11Y4_A_DIN_BRAM0(fabric_bram1_a_din_o[0]),
        .Tile_X11Y4_A_DIN_BRAM1(fabric_bram1_a_din_o[1]),
        .Tile_X11Y4_A_DIN_BRAM2(fabric_bram1_a_din_o[2]),
        .Tile_X11Y4_A_DIN_BRAM3(fabric_bram1_a_din_o[3]),
        .Tile_X11Y4_A_DIN_BRAM4(fabric_bram1_a_din_o[4]),
        .Tile_X11Y4_A_DIN_BRAM5(fabric_bram1_a_din_o[5]),
        .Tile_X11Y4_A_DIN_BRAM6(fabric_bram1_a_din_o[6]),
        .Tile_X11Y4_A_DIN_BRAM7(fabric_bram1_a_din_o[7]),
        .Tile_X11Y4_A_DIN_BRAM8(fabric_bram1_a_din_o[8]),
        .Tile_X11Y4_A_DIN_BRAM9(fabric_bram1_a_din_o[9]),
        .Tile_X11Y4_A_DIN_BRAM10(fabric_bram1_a_din_o[10]),
        .Tile_X11Y4_A_DIN_BRAM11(fabric_bram1_a_din_o[11]),
        .Tile_X11Y4_A_DIN_BRAM12(fabric_bram1_a_din_o[12]),
        .Tile_X11Y4_A_DIN_BRAM13(fabric_bram1_a_din_o[13]),
        .Tile_X11Y4_A_DIN_BRAM14(fabric_bram1_a_din_o[14]),
        .Tile_X11Y4_A_DIN_BRAM15(fabric_bram1_a_din_o[15]),
        .Tile_X11Y4_A_WEN_BRAM(fabric_bram1_a_wen_o),
        .Tile_X11Y4_A_MEN_BRAM(fabric_bram1_a_men_o),
        .Tile_X11Y4_A_REN_BRAM(fabric_bram1_a_ren_o),
        .Tile_X11Y4_A_CLK_BRAM(fabric_bram1_a_clk_o),
        .Tile_X11Y4_A_TIE_HIGH_BRAM(fabric_bram1_a_tie_high_o),
        .Tile_X11Y4_A_TIE_LOW_BRAM(fabric_bram1_a_tie_low_o),

        // Port B
        .Tile_X11Y4_B_DOUT_BRAM0(fabric_bram1_b_dout_i[0]),
        .Tile_X11Y4_B_DOUT_BRAM1(fabric_bram1_b_dout_i[1]),
        .Tile_X11Y4_B_DOUT_BRAM2(fabric_bram1_b_dout_i[2]),
        .Tile_X11Y4_B_DOUT_BRAM3(fabric_bram1_b_dout_i[3]),
        .Tile_X11Y4_B_DOUT_BRAM4(fabric_bram1_b_dout_i[4]),
        .Tile_X11Y4_B_DOUT_BRAM5(fabric_bram1_b_dout_i[5]),
        .Tile_X11Y4_B_DOUT_BRAM6(fabric_bram1_b_dout_i[6]),
        .Tile_X11Y4_B_DOUT_BRAM7(fabric_bram1_b_dout_i[7]),
        .Tile_X11Y4_B_DOUT_BRAM8(fabric_bram1_b_dout_i[8]),
        .Tile_X11Y4_B_DOUT_BRAM9(fabric_bram1_b_dout_i[9]),
        .Tile_X11Y4_B_DOUT_BRAM10(fabric_bram1_b_dout_i[10]),
        .Tile_X11Y4_B_DOUT_BRAM11(fabric_bram1_b_dout_i[11]),
        .Tile_X11Y4_B_DOUT_BRAM12(fabric_bram1_b_dout_i[12]),
        .Tile_X11Y4_B_DOUT_BRAM13(fabric_bram1_b_dout_i[13]),
        .Tile_X11Y4_B_DOUT_BRAM14(fabric_bram1_b_dout_i[14]),
        .Tile_X11Y4_B_DOUT_BRAM15(fabric_bram1_b_dout_i[15]),
        .Tile_X11Y4_B_ADDR_BRAM0(fabric_bram1_b_addr_o[0]),
        .Tile_X11Y4_B_ADDR_BRAM1(fabric_bram1_b_addr_o[1]),
        .Tile_X11Y4_B_ADDR_BRAM2(fabric_bram1_b_addr_o[2]),
        .Tile_X11Y4_B_ADDR_BRAM3(fabric_bram1_b_addr_o[3]),
        .Tile_X11Y4_B_ADDR_BRAM4(fabric_bram1_b_addr_o[4]),
        .Tile_X11Y4_B_ADDR_BRAM5(fabric_bram1_b_addr_o[5]),
        .Tile_X11Y4_B_ADDR_BRAM6(fabric_bram1_b_addr_o[6]),
        .Tile_X11Y4_B_ADDR_BRAM7(fabric_bram1_b_addr_o[7]),
        .Tile_X11Y4_B_ADDR_BRAM8(fabric_bram1_b_addr_o[8]),
        .Tile_X11Y4_B_ADDR_BRAM9(fabric_bram1_b_addr_o[9]),
        .Tile_X11Y4_B_BM_BRAM0(fabric_bram1_b_bm_o[0]),
        .Tile_X11Y4_B_BM_BRAM1(fabric_bram1_b_bm_o[1]),
        .Tile_X11Y4_B_BM_BRAM2(fabric_bram1_b_bm_o[2]),
        .Tile_X11Y4_B_BM_BRAM3(fabric_bram1_b_bm_o[3]),
        .Tile_X11Y4_B_BM_BRAM4(fabric_bram1_b_bm_o[4]),
        .Tile_X11Y4_B_BM_BRAM5(fabric_bram1_b_bm_o[5]),
        .Tile_X11Y4_B_BM_BRAM6(fabric_bram1_b_bm_o[6]),
        .Tile_X11Y4_B_BM_BRAM7(fabric_bram1_b_bm_o[7]),
        .Tile_X11Y4_B_BM_BRAM8(fabric_bram1_b_bm_o[8]),
        .Tile_X11Y4_B_BM_BRAM9(fabric_bram1_b_bm_o[9]),
        .Tile_X11Y4_B_BM_BRAM10(fabric_bram1_b_bm_o[10]),
        .Tile_X11Y4_B_BM_BRAM11(fabric_bram1_b_bm_o[11]),
        .Tile_X11Y4_B_BM_BRAM12(fabric_bram1_b_bm_o[12]),
        .Tile_X11Y4_B_BM_BRAM13(fabric_bram1_b_bm_o[13]),
        .Tile_X11Y4_B_BM_BRAM14(fabric_bram1_b_bm_o[14]),
        .Tile_X11Y4_B_BM_BRAM15(fabric_bram1_b_bm_o[15]),
        .Tile_X11Y4_B_DIN_BRAM0(fabric_bram1_b_din_o[0]),
        .Tile_X11Y4_B_DIN_BRAM1(fabric_bram1_b_din_o[1]),
        .Tile_X11Y4_B_DIN_BRAM2(fabric_bram1_b_din_o[2]),
        .Tile_X11Y4_B_DIN_BRAM3(fabric_bram1_b_din_o[3]),
        .Tile_X11Y4_B_DIN_BRAM4(fabric_bram1_b_din_o[4]),
        .Tile_X11Y4_B_DIN_BRAM5(fabric_bram1_b_din_o[5]),
        .Tile_X11Y4_B_DIN_BRAM6(fabric_bram1_b_din_o[6]),
        .Tile_X11Y4_B_DIN_BRAM7(fabric_bram1_b_din_o[7]),
        .Tile_X11Y4_B_DIN_BRAM8(fabric_bram1_b_din_o[8]),
        .Tile_X11Y4_B_DIN_BRAM9(fabric_bram1_b_din_o[9]),
        .Tile_X11Y4_B_DIN_BRAM10(fabric_bram1_b_din_o[10]),
        .Tile_X11Y4_B_DIN_BRAM11(fabric_bram1_b_din_o[11]),
        .Tile_X11Y4_B_DIN_BRAM12(fabric_bram1_b_din_o[12]),
        .Tile_X11Y4_B_DIN_BRAM13(fabric_bram1_b_din_o[13]),
        .Tile_X11Y4_B_DIN_BRAM14(fabric_bram1_b_din_o[14]),
        .Tile_X11Y4_B_DIN_BRAM15(fabric_bram1_b_din_o[15]),
        .Tile_X11Y4_B_WEN_BRAM(fabric_bram1_b_wen_o),
        .Tile_X11Y4_B_MEN_BRAM(fabric_bram1_b_men_o),
        .Tile_X11Y4_B_REN_BRAM(fabric_bram1_b_ren_o),
        .Tile_X11Y4_B_CLK_BRAM(fabric_bram1_b_clk_o),
        .Tile_X11Y4_B_TIE_HIGH_BRAM(fabric_bram1_b_tie_high_o),
        .Tile_X11Y4_B_TIE_LOW_BRAM(fabric_bram1_b_tie_low_o),

        .Tile_X11Y4_CONFIGURED_top(configured_i),

        // BRAM 2
        // Port A
        .Tile_X11Y6_A_DOUT_BRAM0(fabric_bram2_a_dout_i[0]),
        .Tile_X11Y6_A_DOUT_BRAM1(fabric_bram2_a_dout_i[1]),
        .Tile_X11Y6_A_DOUT_BRAM2(fabric_bram2_a_dout_i[2]),
        .Tile_X11Y6_A_DOUT_BRAM3(fabric_bram2_a_dout_i[3]),
        .Tile_X11Y6_A_DOUT_BRAM4(fabric_bram2_a_dout_i[4]),
        .Tile_X11Y6_A_DOUT_BRAM5(fabric_bram2_a_dout_i[5]),
        .Tile_X11Y6_A_DOUT_BRAM6(fabric_bram2_a_dout_i[6]),
        .Tile_X11Y6_A_DOUT_BRAM7(fabric_bram2_a_dout_i[7]),
        .Tile_X11Y6_A_DOUT_BRAM8(fabric_bram2_a_dout_i[8]),
        .Tile_X11Y6_A_DOUT_BRAM9(fabric_bram2_a_dout_i[9]),
        .Tile_X11Y6_A_DOUT_BRAM10(fabric_bram2_a_dout_i[10]),
        .Tile_X11Y6_A_DOUT_BRAM11(fabric_bram2_a_dout_i[11]),
        .Tile_X11Y6_A_DOUT_BRAM12(fabric_bram2_a_dout_i[12]),
        .Tile_X11Y6_A_DOUT_BRAM13(fabric_bram2_a_dout_i[13]),
        .Tile_X11Y6_A_DOUT_BRAM14(fabric_bram2_a_dout_i[14]),
        .Tile_X11Y6_A_DOUT_BRAM15(fabric_bram2_a_dout_i[15]),
        .Tile_X11Y6_A_ADDR_BRAM0(fabric_bram2_a_addr_o[0]),
        .Tile_X11Y6_A_ADDR_BRAM1(fabric_bram2_a_addr_o[1]),
        .Tile_X11Y6_A_ADDR_BRAM2(fabric_bram2_a_addr_o[2]),
        .Tile_X11Y6_A_ADDR_BRAM3(fabric_bram2_a_addr_o[3]),
        .Tile_X11Y6_A_ADDR_BRAM4(fabric_bram2_a_addr_o[4]),
        .Tile_X11Y6_A_ADDR_BRAM5(fabric_bram2_a_addr_o[5]),
        .Tile_X11Y6_A_ADDR_BRAM6(fabric_bram2_a_addr_o[6]),
        .Tile_X11Y6_A_ADDR_BRAM7(fabric_bram2_a_addr_o[7]),
        .Tile_X11Y6_A_ADDR_BRAM8(fabric_bram2_a_addr_o[8]),
        .Tile_X11Y6_A_ADDR_BRAM9(fabric_bram2_a_addr_o[9]),
        .Tile_X11Y6_A_BM_BRAM0(fabric_bram2_a_bm_o[0]),
        .Tile_X11Y6_A_BM_BRAM1(fabric_bram2_a_bm_o[1]),
        .Tile_X11Y6_A_BM_BRAM2(fabric_bram2_a_bm_o[2]),
        .Tile_X11Y6_A_BM_BRAM3(fabric_bram2_a_bm_o[3]),
        .Tile_X11Y6_A_BM_BRAM4(fabric_bram2_a_bm_o[4]),
        .Tile_X11Y6_A_BM_BRAM5(fabric_bram2_a_bm_o[5]),
        .Tile_X11Y6_A_BM_BRAM6(fabric_bram2_a_bm_o[6]),
        .Tile_X11Y6_A_BM_BRAM7(fabric_bram2_a_bm_o[7]),
        .Tile_X11Y6_A_BM_BRAM8(fabric_bram2_a_bm_o[8]),
        .Tile_X11Y6_A_BM_BRAM9(fabric_bram2_a_bm_o[9]),
        .Tile_X11Y6_A_BM_BRAM10(fabric_bram2_a_bm_o[10]),
        .Tile_X11Y6_A_BM_BRAM11(fabric_bram2_a_bm_o[11]),
        .Tile_X11Y6_A_BM_BRAM12(fabric_bram2_a_bm_o[12]),
        .Tile_X11Y6_A_BM_BRAM13(fabric_bram2_a_bm_o[13]),
        .Tile_X11Y6_A_BM_BRAM14(fabric_bram2_a_bm_o[14]),
        .Tile_X11Y6_A_BM_BRAM15(fabric_bram2_a_bm_o[15]),
        .Tile_X11Y6_A_DIN_BRAM0(fabric_bram2_a_din_o[0]),
        .Tile_X11Y6_A_DIN_BRAM1(fabric_bram2_a_din_o[1]),
        .Tile_X11Y6_A_DIN_BRAM2(fabric_bram2_a_din_o[2]),
        .Tile_X11Y6_A_DIN_BRAM3(fabric_bram2_a_din_o[3]),
        .Tile_X11Y6_A_DIN_BRAM4(fabric_bram2_a_din_o[4]),
        .Tile_X11Y6_A_DIN_BRAM5(fabric_bram2_a_din_o[5]),
        .Tile_X11Y6_A_DIN_BRAM6(fabric_bram2_a_din_o[6]),
        .Tile_X11Y6_A_DIN_BRAM7(fabric_bram2_a_din_o[7]),
        .Tile_X11Y6_A_DIN_BRAM8(fabric_bram2_a_din_o[8]),
        .Tile_X11Y6_A_DIN_BRAM9(fabric_bram2_a_din_o[9]),
        .Tile_X11Y6_A_DIN_BRAM10(fabric_bram2_a_din_o[10]),
        .Tile_X11Y6_A_DIN_BRAM11(fabric_bram2_a_din_o[11]),
        .Tile_X11Y6_A_DIN_BRAM12(fabric_bram2_a_din_o[12]),
        .Tile_X11Y6_A_DIN_BRAM13(fabric_bram2_a_din_o[13]),
        .Tile_X11Y6_A_DIN_BRAM14(fabric_bram2_a_din_o[14]),
        .Tile_X11Y6_A_DIN_BRAM15(fabric_bram2_a_din_o[15]),
        .Tile_X11Y6_A_WEN_BRAM(fabric_bram2_a_wen_o),
        .Tile_X11Y6_A_MEN_BRAM(fabric_bram2_a_men_o),
        .Tile_X11Y6_A_REN_BRAM(fabric_bram2_a_ren_o),
        .Tile_X11Y6_A_CLK_BRAM(fabric_bram2_a_clk_o),
        .Tile_X11Y6_A_TIE_HIGH_BRAM(fabric_bram2_a_tie_high_o),
        .Tile_X11Y6_A_TIE_LOW_BRAM(fabric_bram2_a_tie_low_o),

        // Port B
        .Tile_X11Y6_B_DOUT_BRAM0(fabric_bram2_b_dout_i[0]),
        .Tile_X11Y6_B_DOUT_BRAM1(fabric_bram2_b_dout_i[1]),
        .Tile_X11Y6_B_DOUT_BRAM2(fabric_bram2_b_dout_i[2]),
        .Tile_X11Y6_B_DOUT_BRAM3(fabric_bram2_b_dout_i[3]),
        .Tile_X11Y6_B_DOUT_BRAM4(fabric_bram2_b_dout_i[4]),
        .Tile_X11Y6_B_DOUT_BRAM5(fabric_bram2_b_dout_i[5]),
        .Tile_X11Y6_B_DOUT_BRAM6(fabric_bram2_b_dout_i[6]),
        .Tile_X11Y6_B_DOUT_BRAM7(fabric_bram2_b_dout_i[7]),
        .Tile_X11Y6_B_DOUT_BRAM8(fabric_bram2_b_dout_i[8]),
        .Tile_X11Y6_B_DOUT_BRAM9(fabric_bram2_b_dout_i[9]),
        .Tile_X11Y6_B_DOUT_BRAM10(fabric_bram2_b_dout_i[10]),
        .Tile_X11Y6_B_DOUT_BRAM11(fabric_bram2_b_dout_i[11]),
        .Tile_X11Y6_B_DOUT_BRAM12(fabric_bram2_b_dout_i[12]),
        .Tile_X11Y6_B_DOUT_BRAM13(fabric_bram2_b_dout_i[13]),
        .Tile_X11Y6_B_DOUT_BRAM14(fabric_bram2_b_dout_i[14]),
        .Tile_X11Y6_B_DOUT_BRAM15(fabric_bram2_b_dout_i[15]),
        .Tile_X11Y6_B_ADDR_BRAM0(fabric_bram2_b_addr_o[0]),
        .Tile_X11Y6_B_ADDR_BRAM1(fabric_bram2_b_addr_o[1]),
        .Tile_X11Y6_B_ADDR_BRAM2(fabric_bram2_b_addr_o[2]),
        .Tile_X11Y6_B_ADDR_BRAM3(fabric_bram2_b_addr_o[3]),
        .Tile_X11Y6_B_ADDR_BRAM4(fabric_bram2_b_addr_o[4]),
        .Tile_X11Y6_B_ADDR_BRAM5(fabric_bram2_b_addr_o[5]),
        .Tile_X11Y6_B_ADDR_BRAM6(fabric_bram2_b_addr_o[6]),
        .Tile_X11Y6_B_ADDR_BRAM7(fabric_bram2_b_addr_o[7]),
        .Tile_X11Y6_B_ADDR_BRAM8(fabric_bram2_b_addr_o[8]),
        .Tile_X11Y6_B_ADDR_BRAM9(fabric_bram2_b_addr_o[9]),
        .Tile_X11Y6_B_BM_BRAM0(fabric_bram2_b_bm_o[0]),
        .Tile_X11Y6_B_BM_BRAM1(fabric_bram2_b_bm_o[1]),
        .Tile_X11Y6_B_BM_BRAM2(fabric_bram2_b_bm_o[2]),
        .Tile_X11Y6_B_BM_BRAM3(fabric_bram2_b_bm_o[3]),
        .Tile_X11Y6_B_BM_BRAM4(fabric_bram2_b_bm_o[4]),
        .Tile_X11Y6_B_BM_BRAM5(fabric_bram2_b_bm_o[5]),
        .Tile_X11Y6_B_BM_BRAM6(fabric_bram2_b_bm_o[6]),
        .Tile_X11Y6_B_BM_BRAM7(fabric_bram2_b_bm_o[7]),
        .Tile_X11Y6_B_BM_BRAM8(fabric_bram2_b_bm_o[8]),
        .Tile_X11Y6_B_BM_BRAM9(fabric_bram2_b_bm_o[9]),
        .Tile_X11Y6_B_BM_BRAM10(fabric_bram2_b_bm_o[10]),
        .Tile_X11Y6_B_BM_BRAM11(fabric_bram2_b_bm_o[11]),
        .Tile_X11Y6_B_BM_BRAM12(fabric_bram2_b_bm_o[12]),
        .Tile_X11Y6_B_BM_BRAM13(fabric_bram2_b_bm_o[13]),
        .Tile_X11Y6_B_BM_BRAM14(fabric_bram2_b_bm_o[14]),
        .Tile_X11Y6_B_BM_BRAM15(fabric_bram2_b_bm_o[15]),
        .Tile_X11Y6_B_DIN_BRAM0(fabric_bram2_b_din_o[0]),
        .Tile_X11Y6_B_DIN_BRAM1(fabric_bram2_b_din_o[1]),
        .Tile_X11Y6_B_DIN_BRAM2(fabric_bram2_b_din_o[2]),
        .Tile_X11Y6_B_DIN_BRAM3(fabric_bram2_b_din_o[3]),
        .Tile_X11Y6_B_DIN_BRAM4(fabric_bram2_b_din_o[4]),
        .Tile_X11Y6_B_DIN_BRAM5(fabric_bram2_b_din_o[5]),
        .Tile_X11Y6_B_DIN_BRAM6(fabric_bram2_b_din_o[6]),
        .Tile_X11Y6_B_DIN_BRAM7(fabric_bram2_b_din_o[7]),
        .Tile_X11Y6_B_DIN_BRAM8(fabric_bram2_b_din_o[8]),
        .Tile_X11Y6_B_DIN_BRAM9(fabric_bram2_b_din_o[9]),
        .Tile_X11Y6_B_DIN_BRAM10(fabric_bram2_b_din_o[10]),
        .Tile_X11Y6_B_DIN_BRAM11(fabric_bram2_b_din_o[11]),
        .Tile_X11Y6_B_DIN_BRAM12(fabric_bram2_b_din_o[12]),
        .Tile_X11Y6_B_DIN_BRAM13(fabric_bram2_b_din_o[13]),
        .Tile_X11Y6_B_DIN_BRAM14(fabric_bram2_b_din_o[14]),
        .Tile_X11Y6_B_DIN_BRAM15(fabric_bram2_b_din_o[15]),
        .Tile_X11Y6_B_WEN_BRAM(fabric_bram2_b_wen_o),
        .Tile_X11Y6_B_MEN_BRAM(fabric_bram2_b_men_o),
        .Tile_X11Y6_B_REN_BRAM(fabric_bram2_b_ren_o),
        .Tile_X11Y6_B_CLK_BRAM(fabric_bram2_b_clk_o),
        .Tile_X11Y6_B_TIE_HIGH_BRAM(fabric_bram2_b_tie_high_o),
        .Tile_X11Y6_B_TIE_LOW_BRAM(fabric_bram2_b_tie_low_o),

        .Tile_X11Y6_CONFIGURED_top(configured_i),

        // BRAM 3
        // Port A
        .Tile_X11Y8_A_DOUT_BRAM0(fabric_bram3_a_dout_i[0]),
        .Tile_X11Y8_A_DOUT_BRAM1(fabric_bram3_a_dout_i[1]),
        .Tile_X11Y8_A_DOUT_BRAM2(fabric_bram3_a_dout_i[2]),
        .Tile_X11Y8_A_DOUT_BRAM3(fabric_bram3_a_dout_i[3]),
        .Tile_X11Y8_A_DOUT_BRAM4(fabric_bram3_a_dout_i[4]),
        .Tile_X11Y8_A_DOUT_BRAM5(fabric_bram3_a_dout_i[5]),
        .Tile_X11Y8_A_DOUT_BRAM6(fabric_bram3_a_dout_i[6]),
        .Tile_X11Y8_A_DOUT_BRAM7(fabric_bram3_a_dout_i[7]),
        .Tile_X11Y8_A_DOUT_BRAM8(fabric_bram3_a_dout_i[8]),
        .Tile_X11Y8_A_DOUT_BRAM9(fabric_bram3_a_dout_i[9]),
        .Tile_X11Y8_A_DOUT_BRAM10(fabric_bram3_a_dout_i[10]),
        .Tile_X11Y8_A_DOUT_BRAM11(fabric_bram3_a_dout_i[11]),
        .Tile_X11Y8_A_DOUT_BRAM12(fabric_bram3_a_dout_i[12]),
        .Tile_X11Y8_A_DOUT_BRAM13(fabric_bram3_a_dout_i[13]),
        .Tile_X11Y8_A_DOUT_BRAM14(fabric_bram3_a_dout_i[14]),
        .Tile_X11Y8_A_DOUT_BRAM15(fabric_bram3_a_dout_i[15]),
        .Tile_X11Y8_A_ADDR_BRAM0(fabric_bram3_a_addr_o[0]),
        .Tile_X11Y8_A_ADDR_BRAM1(fabric_bram3_a_addr_o[1]),
        .Tile_X11Y8_A_ADDR_BRAM2(fabric_bram3_a_addr_o[2]),
        .Tile_X11Y8_A_ADDR_BRAM3(fabric_bram3_a_addr_o[3]),
        .Tile_X11Y8_A_ADDR_BRAM4(fabric_bram3_a_addr_o[4]),
        .Tile_X11Y8_A_ADDR_BRAM5(fabric_bram3_a_addr_o[5]),
        .Tile_X11Y8_A_ADDR_BRAM6(fabric_bram3_a_addr_o[6]),
        .Tile_X11Y8_A_ADDR_BRAM7(fabric_bram3_a_addr_o[7]),
        .Tile_X11Y8_A_ADDR_BRAM8(fabric_bram3_a_addr_o[8]),
        .Tile_X11Y8_A_ADDR_BRAM9(fabric_bram3_a_addr_o[9]),
        .Tile_X11Y8_A_BM_BRAM0(fabric_bram3_a_bm_o[0]),
        .Tile_X11Y8_A_BM_BRAM1(fabric_bram3_a_bm_o[1]),
        .Tile_X11Y8_A_BM_BRAM2(fabric_bram3_a_bm_o[2]),
        .Tile_X11Y8_A_BM_BRAM3(fabric_bram3_a_bm_o[3]),
        .Tile_X11Y8_A_BM_BRAM4(fabric_bram3_a_bm_o[4]),
        .Tile_X11Y8_A_BM_BRAM5(fabric_bram3_a_bm_o[5]),
        .Tile_X11Y8_A_BM_BRAM6(fabric_bram3_a_bm_o[6]),
        .Tile_X11Y8_A_BM_BRAM7(fabric_bram3_a_bm_o[7]),
        .Tile_X11Y8_A_BM_BRAM8(fabric_bram3_a_bm_o[8]),
        .Tile_X11Y8_A_BM_BRAM9(fabric_bram3_a_bm_o[9]),
        .Tile_X11Y8_A_BM_BRAM10(fabric_bram3_a_bm_o[10]),
        .Tile_X11Y8_A_BM_BRAM11(fabric_bram3_a_bm_o[11]),
        .Tile_X11Y8_A_BM_BRAM12(fabric_bram3_a_bm_o[12]),
        .Tile_X11Y8_A_BM_BRAM13(fabric_bram3_a_bm_o[13]),
        .Tile_X11Y8_A_BM_BRAM14(fabric_bram3_a_bm_o[14]),
        .Tile_X11Y8_A_BM_BRAM15(fabric_bram3_a_bm_o[15]),
        .Tile_X11Y8_A_DIN_BRAM0(fabric_bram3_a_din_o[0]),
        .Tile_X11Y8_A_DIN_BRAM1(fabric_bram3_a_din_o[1]),
        .Tile_X11Y8_A_DIN_BRAM2(fabric_bram3_a_din_o[2]),
        .Tile_X11Y8_A_DIN_BRAM3(fabric_bram3_a_din_o[3]),
        .Tile_X11Y8_A_DIN_BRAM4(fabric_bram3_a_din_o[4]),
        .Tile_X11Y8_A_DIN_BRAM5(fabric_bram3_a_din_o[5]),
        .Tile_X11Y8_A_DIN_BRAM6(fabric_bram3_a_din_o[6]),
        .Tile_X11Y8_A_DIN_BRAM7(fabric_bram3_a_din_o[7]),
        .Tile_X11Y8_A_DIN_BRAM8(fabric_bram3_a_din_o[8]),
        .Tile_X11Y8_A_DIN_BRAM9(fabric_bram3_a_din_o[9]),
        .Tile_X11Y8_A_DIN_BRAM10(fabric_bram3_a_din_o[10]),
        .Tile_X11Y8_A_DIN_BRAM11(fabric_bram3_a_din_o[11]),
        .Tile_X11Y8_A_DIN_BRAM12(fabric_bram3_a_din_o[12]),
        .Tile_X11Y8_A_DIN_BRAM13(fabric_bram3_a_din_o[13]),
        .Tile_X11Y8_A_DIN_BRAM14(fabric_bram3_a_din_o[14]),
        .Tile_X11Y8_A_DIN_BRAM15(fabric_bram3_a_din_o[15]),
        .Tile_X11Y8_A_WEN_BRAM(fabric_bram3_a_wen_o),
        .Tile_X11Y8_A_MEN_BRAM(fabric_bram3_a_men_o),
        .Tile_X11Y8_A_REN_BRAM(fabric_bram3_a_ren_o),
        .Tile_X11Y8_A_CLK_BRAM(fabric_bram3_a_clk_o),
        .Tile_X11Y8_A_TIE_HIGH_BRAM(fabric_bram3_a_tie_high_o),
        .Tile_X11Y8_A_TIE_LOW_BRAM(fabric_bram3_a_tie_low_o),

        // Port B
        .Tile_X11Y8_B_DOUT_BRAM0(fabric_bram3_b_dout_i[0]),
        .Tile_X11Y8_B_DOUT_BRAM1(fabric_bram3_b_dout_i[1]),
        .Tile_X11Y8_B_DOUT_BRAM2(fabric_bram3_b_dout_i[2]),
        .Tile_X11Y8_B_DOUT_BRAM3(fabric_bram3_b_dout_i[3]),
        .Tile_X11Y8_B_DOUT_BRAM4(fabric_bram3_b_dout_i[4]),
        .Tile_X11Y8_B_DOUT_BRAM5(fabric_bram3_b_dout_i[5]),
        .Tile_X11Y8_B_DOUT_BRAM6(fabric_bram3_b_dout_i[6]),
        .Tile_X11Y8_B_DOUT_BRAM7(fabric_bram3_b_dout_i[7]),
        .Tile_X11Y8_B_DOUT_BRAM8(fabric_bram3_b_dout_i[8]),
        .Tile_X11Y8_B_DOUT_BRAM9(fabric_bram3_b_dout_i[9]),
        .Tile_X11Y8_B_DOUT_BRAM10(fabric_bram3_b_dout_i[10]),
        .Tile_X11Y8_B_DOUT_BRAM11(fabric_bram3_b_dout_i[11]),
        .Tile_X11Y8_B_DOUT_BRAM12(fabric_bram3_b_dout_i[12]),
        .Tile_X11Y8_B_DOUT_BRAM13(fabric_bram3_b_dout_i[13]),
        .Tile_X11Y8_B_DOUT_BRAM14(fabric_bram3_b_dout_i[14]),
        .Tile_X11Y8_B_DOUT_BRAM15(fabric_bram3_b_dout_i[15]),
        .Tile_X11Y8_B_ADDR_BRAM0(fabric_bram3_b_addr_o[0]),
        .Tile_X11Y8_B_ADDR_BRAM1(fabric_bram3_b_addr_o[1]),
        .Tile_X11Y8_B_ADDR_BRAM2(fabric_bram3_b_addr_o[2]),
        .Tile_X11Y8_B_ADDR_BRAM3(fabric_bram3_b_addr_o[3]),
        .Tile_X11Y8_B_ADDR_BRAM4(fabric_bram3_b_addr_o[4]),
        .Tile_X11Y8_B_ADDR_BRAM5(fabric_bram3_b_addr_o[5]),
        .Tile_X11Y8_B_ADDR_BRAM6(fabric_bram3_b_addr_o[6]),
        .Tile_X11Y8_B_ADDR_BRAM7(fabric_bram3_b_addr_o[7]),
        .Tile_X11Y8_B_ADDR_BRAM8(fabric_bram3_b_addr_o[8]),
        .Tile_X11Y8_B_ADDR_BRAM9(fabric_bram3_b_addr_o[9]),
        .Tile_X11Y8_B_BM_BRAM0(fabric_bram3_b_bm_o[0]),
        .Tile_X11Y8_B_BM_BRAM1(fabric_bram3_b_bm_o[1]),
        .Tile_X11Y8_B_BM_BRAM2(fabric_bram3_b_bm_o[2]),
        .Tile_X11Y8_B_BM_BRAM3(fabric_bram3_b_bm_o[3]),
        .Tile_X11Y8_B_BM_BRAM4(fabric_bram3_b_bm_o[4]),
        .Tile_X11Y8_B_BM_BRAM5(fabric_bram3_b_bm_o[5]),
        .Tile_X11Y8_B_BM_BRAM6(fabric_bram3_b_bm_o[6]),
        .Tile_X11Y8_B_BM_BRAM7(fabric_bram3_b_bm_o[7]),
        .Tile_X11Y8_B_BM_BRAM8(fabric_bram3_b_bm_o[8]),
        .Tile_X11Y8_B_BM_BRAM9(fabric_bram3_b_bm_o[9]),
        .Tile_X11Y8_B_BM_BRAM10(fabric_bram3_b_bm_o[10]),
        .Tile_X11Y8_B_BM_BRAM11(fabric_bram3_b_bm_o[11]),
        .Tile_X11Y8_B_BM_BRAM12(fabric_bram3_b_bm_o[12]),
        .Tile_X11Y8_B_BM_BRAM13(fabric_bram3_b_bm_o[13]),
        .Tile_X11Y8_B_BM_BRAM14(fabric_bram3_b_bm_o[14]),
        .Tile_X11Y8_B_BM_BRAM15(fabric_bram3_b_bm_o[15]),
        .Tile_X11Y8_B_DIN_BRAM0(fabric_bram3_b_din_o[0]),
        .Tile_X11Y8_B_DIN_BRAM1(fabric_bram3_b_din_o[1]),
        .Tile_X11Y8_B_DIN_BRAM2(fabric_bram3_b_din_o[2]),
        .Tile_X11Y8_B_DIN_BRAM3(fabric_bram3_b_din_o[3]),
        .Tile_X11Y8_B_DIN_BRAM4(fabric_bram3_b_din_o[4]),
        .Tile_X11Y8_B_DIN_BRAM5(fabric_bram3_b_din_o[5]),
        .Tile_X11Y8_B_DIN_BRAM6(fabric_bram3_b_din_o[6]),
        .Tile_X11Y8_B_DIN_BRAM7(fabric_bram3_b_din_o[7]),
        .Tile_X11Y8_B_DIN_BRAM8(fabric_bram3_b_din_o[8]),
        .Tile_X11Y8_B_DIN_BRAM9(fabric_bram3_b_din_o[9]),
        .Tile_X11Y8_B_DIN_BRAM10(fabric_bram3_b_din_o[10]),
        .Tile_X11Y8_B_DIN_BRAM11(fabric_bram3_b_din_o[11]),
        .Tile_X11Y8_B_DIN_BRAM12(fabric_bram3_b_din_o[12]),
        .Tile_X11Y8_B_DIN_BRAM13(fabric_bram3_b_din_o[13]),
        .Tile_X11Y8_B_DIN_BRAM14(fabric_bram3_b_din_o[14]),
        .Tile_X11Y8_B_DIN_BRAM15(fabric_bram3_b_din_o[15]),
        .Tile_X11Y8_B_WEN_BRAM(fabric_bram3_b_wen_o),
        .Tile_X11Y8_B_MEN_BRAM(fabric_bram3_b_men_o),
        .Tile_X11Y8_B_REN_BRAM(fabric_bram3_b_ren_o),
        .Tile_X11Y8_B_CLK_BRAM(fabric_bram3_b_clk_o),
        .Tile_X11Y8_B_TIE_HIGH_BRAM(fabric_bram3_b_tie_high_o),
        .Tile_X11Y8_B_TIE_LOW_BRAM(fabric_bram3_b_tie_low_o),

        .Tile_X11Y8_CONFIGURED_top(configured_i)
    );

    // SRAM 0 instances

    RM_IHPSG13_1P_1024x32_c2_bm_bist sram0 (
        .A_CLK      (fabric_sram0_a_clk_o),
        .A_MEN      (fabric_sram0_a_men_o),
        .A_WEN      (fabric_sram0_a_wen_o),
        .A_REN      (fabric_sram0_a_ren_o),
        .A_ADDR     (fabric_sram0_a_addr_o),
        .A_DIN      (fabric_sram0_a_din_o),
        .A_DLY      (fabric_sram0_a_tie_high_o),
        .A_DOUT     (fabric_sram0_a_dout_i),
        .A_BM       (fabric_sram0_a_bm_o),

        .A_BIST_EN      (fabric_sram0_a_tie_low_o),
        .A_BIST_CLK     (fabric_sram0_a_tie_low_o),
        .A_BIST_MEN     (fabric_sram0_a_tie_low_o),
        .A_BIST_WEN     (fabric_sram0_a_tie_low_o),
        .A_BIST_REN     (fabric_sram0_a_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram0_a_tie_low_o}}),
        .A_BIST_DIN     ({32{fabric_sram0_a_tie_low_o}}),
        .A_BIST_BM      ({32{fabric_sram0_a_tie_low_o}})
    );

    // SRAM 1 instances

    RM_IHPSG13_1P_1024x32_c2_bm_bist sram1 (
        .A_CLK      (fabric_sram1_a_clk_o),
        .A_MEN      (fabric_sram1_a_men_o),
        .A_WEN      (fabric_sram1_a_wen_o),
        .A_REN      (fabric_sram1_a_ren_o),
        .A_ADDR     (fabric_sram1_a_addr_o),
        .A_DIN      (fabric_sram1_a_din_o),
        .A_DLY      (fabric_sram1_a_tie_high_o),
        .A_DOUT     (fabric_sram1_a_dout_i),
        .A_BM       (fabric_sram1_a_bm_o),

        .A_BIST_EN      (fabric_sram1_a_tie_low_o),
        .A_BIST_CLK     (fabric_sram1_a_tie_low_o),
        .A_BIST_MEN     (fabric_sram1_a_tie_low_o),
        .A_BIST_WEN     (fabric_sram1_a_tie_low_o),
        .A_BIST_REN     (fabric_sram1_a_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram1_a_tie_low_o}}),
        .A_BIST_DIN     ({32{fabric_sram1_a_tie_low_o}}),
        .A_BIST_BM      ({32{fabric_sram1_a_tie_low_o}})
    );

    // SRAM 2 instances

    RM_IHPSG13_1P_1024x32_c2_bm_bist sram2 (
        .A_CLK      (fabric_sram2_a_clk_o),
        .A_MEN      (fabric_sram2_a_men_o),
        .A_WEN      (fabric_sram2_a_wen_o),
        .A_REN      (fabric_sram2_a_ren_o),
        .A_ADDR     (fabric_sram2_a_addr_o),
        .A_DIN      (fabric_sram2_a_din_o),
        .A_DLY      (fabric_sram2_a_tie_high_o),
        .A_DOUT     (fabric_sram2_a_dout_i),
        .A_BM       (fabric_sram2_a_bm_o),

        .A_BIST_EN      (fabric_sram2_a_tie_low_o),
        .A_BIST_CLK     (fabric_sram2_a_tie_low_o),
        .A_BIST_MEN     (fabric_sram2_a_tie_low_o),
        .A_BIST_WEN     (fabric_sram2_a_tie_low_o),
        .A_BIST_REN     (fabric_sram2_a_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram2_a_tie_low_o}}),
        .A_BIST_DIN     ({32{fabric_sram2_a_tie_low_o}}),
        .A_BIST_BM      ({32{fabric_sram2_a_tie_low_o}})
    );

    // SRAM 3 instances

    RM_IHPSG13_1P_1024x32_c2_bm_bist sram3 (
        .A_CLK      (fabric_sram3_a_clk_o),
        .A_MEN      (fabric_sram3_a_men_o),
        .A_WEN      (fabric_sram3_a_wen_o),
        .A_REN      (fabric_sram3_a_ren_o),
        .A_ADDR     (fabric_sram3_a_addr_o),
        .A_DIN      (fabric_sram3_a_din_o),
        .A_DLY      (fabric_sram3_a_tie_high_o),
        .A_DOUT     (fabric_sram3_a_dout_i),
        .A_BM       (fabric_sram3_a_bm_o),

        .A_BIST_EN      (fabric_sram3_a_tie_low_o),
        .A_BIST_CLK     (fabric_sram3_a_tie_low_o),
        .A_BIST_MEN     (fabric_sram3_a_tie_low_o),
        .A_BIST_WEN     (fabric_sram3_a_tie_low_o),
        .A_BIST_REN     (fabric_sram3_a_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram3_a_tie_low_o}}),
        .A_BIST_DIN     ({32{fabric_sram3_a_tie_low_o}}),
        .A_BIST_BM      ({32{fabric_sram3_a_tie_low_o}})
    );

    // BRAM 0 instances

    RM_IHPSG13_2P_1024x16_c2_bm_bist bram0 (
        .A_CLK      (fabric_bram0_a_clk_o),
        .A_MEN      (fabric_bram0_a_men_o),
        .A_WEN      (fabric_bram0_a_wen_o),
        .A_REN      (fabric_bram0_a_ren_o),
        .A_ADDR     (fabric_bram0_a_addr_o),
        .A_DIN      (fabric_bram0_a_din_o),
        .A_DLY      (fabric_bram0_a_tie_high_o),
        .A_DOUT     (fabric_bram0_a_dout_i),
        .A_BM       (fabric_bram0_a_bm_o),

        .A_BIST_EN      (fabric_bram0_a_tie_low_o),
        .A_BIST_CLK     (fabric_bram0_a_tie_low_o),
        .A_BIST_MEN     (fabric_bram0_a_tie_low_o),
        .A_BIST_WEN     (fabric_bram0_a_tie_low_o),
        .A_BIST_REN     (fabric_bram0_a_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_bram0_a_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_bram0_a_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_bram0_a_tie_low_o}}),

        .B_CLK      (fabric_bram0_b_clk_o),
        .B_MEN      (fabric_bram0_b_men_o),
        .B_WEN      (fabric_bram0_b_wen_o),
        .B_REN      (fabric_bram0_b_ren_o),
        .B_ADDR     (fabric_bram0_b_addr_o),
        .B_DIN      (fabric_bram0_b_din_o),
        .B_DLY      (fabric_bram0_b_tie_high_o),
        .B_DOUT     (fabric_bram0_b_dout_i),
        .B_BM       (fabric_bram0_b_bm_o),

        .B_BIST_EN      (fabric_bram0_b_tie_low_o),
        .B_BIST_CLK     (fabric_bram0_b_tie_low_o),
        .B_BIST_MEN     (fabric_bram0_b_tie_low_o),
        .B_BIST_WEN     (fabric_bram0_b_tie_low_o),
        .B_BIST_REN     (fabric_bram0_b_tie_low_o),
        .B_BIST_ADDR    ({10{fabric_bram0_b_tie_low_o}}),
        .B_BIST_DIN     ({16{fabric_bram0_b_tie_low_o}}),
        .B_BIST_BM      ({16{fabric_bram0_b_tie_low_o}})
    );

    // BRAM 1 instances

    RM_IHPSG13_2P_1024x16_c2_bm_bist bram1 (
        .A_CLK      (fabric_bram1_a_clk_o),
        .A_MEN      (fabric_bram1_a_men_o),
        .A_WEN      (fabric_bram1_a_wen_o),
        .A_REN      (fabric_bram1_a_ren_o),
        .A_ADDR     (fabric_bram1_a_addr_o),
        .A_DIN      (fabric_bram1_a_din_o),
        .A_DLY      (fabric_bram1_a_tie_high_o),
        .A_DOUT     (fabric_bram1_a_dout_i),
        .A_BM       (fabric_bram1_a_bm_o),

        .A_BIST_EN      (fabric_bram1_a_tie_low_o),
        .A_BIST_CLK     (fabric_bram1_a_tie_low_o),
        .A_BIST_MEN     (fabric_bram1_a_tie_low_o),
        .A_BIST_WEN     (fabric_bram1_a_tie_low_o),
        .A_BIST_REN     (fabric_bram1_a_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_bram1_a_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_bram1_a_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_bram1_a_tie_low_o}}),

        .B_CLK      (fabric_bram1_b_clk_o),
        .B_MEN      (fabric_bram1_b_men_o),
        .B_WEN      (fabric_bram1_b_wen_o),
        .B_REN      (fabric_bram1_b_ren_o),
        .B_ADDR     (fabric_bram1_b_addr_o),
        .B_DIN      (fabric_bram1_b_din_o),
        .B_DLY      (fabric_bram1_b_tie_high_o),
        .B_DOUT     (fabric_bram1_b_dout_i),
        .B_BM       (fabric_bram1_b_bm_o),

        .B_BIST_EN      (fabric_bram1_b_tie_low_o),
        .B_BIST_CLK     (fabric_bram1_b_tie_low_o),
        .B_BIST_MEN     (fabric_bram1_b_tie_low_o),
        .B_BIST_WEN     (fabric_bram1_b_tie_low_o),
        .B_BIST_REN     (fabric_bram1_b_tie_low_o),
        .B_BIST_ADDR    ({10{fabric_bram1_b_tie_low_o}}),
        .B_BIST_DIN     ({16{fabric_bram1_b_tie_low_o}}),
        .B_BIST_BM      ({16{fabric_bram1_b_tie_low_o}})
    );

    // BRAM 2 instances

    RM_IHPSG13_2P_1024x16_c2_bm_bist bram2 (
        .A_CLK      (fabric_bram2_a_clk_o),
        .A_MEN      (fabric_bram2_a_men_o),
        .A_WEN      (fabric_bram2_a_wen_o),
        .A_REN      (fabric_bram2_a_ren_o),
        .A_ADDR     (fabric_bram2_a_addr_o),
        .A_DIN      (fabric_bram2_a_din_o),
        .A_DLY      (fabric_bram2_a_tie_high_o),
        .A_DOUT     (fabric_bram2_a_dout_i),
        .A_BM       (fabric_bram2_a_bm_o),

        .A_BIST_EN      (fabric_bram2_a_tie_low_o),
        .A_BIST_CLK     (fabric_bram2_a_tie_low_o),
        .A_BIST_MEN     (fabric_bram2_a_tie_low_o),
        .A_BIST_WEN     (fabric_bram2_a_tie_low_o),
        .A_BIST_REN     (fabric_bram2_a_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_bram2_a_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_bram2_a_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_bram2_a_tie_low_o}}),

        .B_CLK      (fabric_bram2_b_clk_o),
        .B_MEN      (fabric_bram2_b_men_o),
        .B_WEN      (fabric_bram2_b_wen_o),
        .B_REN      (fabric_bram2_b_ren_o),
        .B_ADDR     (fabric_bram2_b_addr_o),
        .B_DIN      (fabric_bram2_b_din_o),
        .B_DLY      (fabric_bram2_b_tie_high_o),
        .B_DOUT     (fabric_bram2_b_dout_i),
        .B_BM       (fabric_bram2_b_bm_o),

        .B_BIST_EN      (fabric_bram2_b_tie_low_o),
        .B_BIST_CLK     (fabric_bram2_b_tie_low_o),
        .B_BIST_MEN     (fabric_bram2_b_tie_low_o),
        .B_BIST_WEN     (fabric_bram2_b_tie_low_o),
        .B_BIST_REN     (fabric_bram2_b_tie_low_o),
        .B_BIST_ADDR    ({10{fabric_bram2_b_tie_low_o}}),
        .B_BIST_DIN     ({16{fabric_bram2_b_tie_low_o}}),
        .B_BIST_BM      ({16{fabric_bram2_b_tie_low_o}})
    );

    // BRAM 3 instances

    RM_IHPSG13_2P_1024x16_c2_bm_bist bram3 (
        .A_CLK      (fabric_bram3_a_clk_o),
        .A_MEN      (fabric_bram3_a_men_o),
        .A_WEN      (fabric_bram3_a_wen_o),
        .A_REN      (fabric_bram3_a_ren_o),
        .A_ADDR     (fabric_bram3_a_addr_o),
        .A_DIN      (fabric_bram3_a_din_o),
        .A_DLY      (fabric_bram3_a_tie_high_o),
        .A_DOUT     (fabric_bram3_a_dout_i),
        .A_BM       (fabric_bram3_a_bm_o),

        .A_BIST_EN      (fabric_bram3_a_tie_low_o),
        .A_BIST_CLK     (fabric_bram3_a_tie_low_o),
        .A_BIST_MEN     (fabric_bram3_a_tie_low_o),
        .A_BIST_WEN     (fabric_bram3_a_tie_low_o),
        .A_BIST_REN     (fabric_bram3_a_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_bram3_a_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_bram3_a_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_bram3_a_tie_low_o}}),

        .B_CLK      (fabric_bram3_b_clk_o),
        .B_MEN      (fabric_bram3_b_men_o),
        .B_WEN      (fabric_bram3_b_wen_o),
        .B_REN      (fabric_bram3_b_ren_o),
        .B_ADDR     (fabric_bram3_b_addr_o),
        .B_DIN      (fabric_bram3_b_din_o),
        .B_DLY      (fabric_bram3_b_tie_high_o),
        .B_DOUT     (fabric_bram3_b_dout_i),
        .B_BM       (fabric_bram3_b_bm_o),

        .B_BIST_EN      (fabric_bram3_b_tie_low_o),
        .B_BIST_CLK     (fabric_bram3_b_tie_low_o),
        .B_BIST_MEN     (fabric_bram3_b_tie_low_o),
        .B_BIST_WEN     (fabric_bram3_b_tie_low_o),
        .B_BIST_REN     (fabric_bram3_b_tie_low_o),
        .B_BIST_ADDR    ({10{fabric_bram3_b_tie_low_o}}),
        .B_BIST_DIN     ({16{fabric_bram3_b_tie_low_o}}),
        .B_BIST_BM      ({16{fabric_bram3_b_tie_low_o}})
    );


endmodule

`default_nettype wire
