magic
tech gf180mcuD
magscale 1 5
timestamp 1764971563
<< metal1 >>
rect 336 6677 15512 6694
rect 336 6651 2233 6677
rect 2259 6651 2285 6677
rect 2311 6651 2337 6677
rect 2363 6651 12233 6677
rect 12259 6651 12285 6677
rect 12311 6651 12337 6677
rect 12363 6651 15512 6677
rect 336 6634 15512 6651
rect 1079 6593 1105 6599
rect 1079 6561 1105 6567
rect 1863 6593 1889 6599
rect 1863 6561 1889 6567
rect 2983 6593 3009 6599
rect 2983 6561 3009 6567
rect 3767 6593 3793 6599
rect 3767 6561 3793 6567
rect 4887 6593 4913 6599
rect 4887 6561 4913 6567
rect 5671 6593 5697 6599
rect 5671 6561 5697 6567
rect 6567 6593 6593 6599
rect 6567 6561 6593 6567
rect 7015 6593 7041 6599
rect 7015 6561 7041 6567
rect 7855 6593 7881 6599
rect 7855 6561 7881 6567
rect 8135 6593 8161 6599
rect 8135 6561 8161 6567
rect 8247 6593 8273 6599
rect 8247 6561 8273 6567
rect 8751 6593 8777 6599
rect 8751 6561 8777 6567
rect 9255 6593 9281 6599
rect 9255 6561 9281 6567
rect 9479 6593 9505 6599
rect 9479 6561 9505 6567
rect 11271 6593 11297 6599
rect 11271 6561 11297 6567
rect 12223 6593 12249 6599
rect 12223 6561 12249 6567
rect 13007 6593 13033 6599
rect 13007 6561 13033 6567
rect 14127 6593 14153 6599
rect 14127 6561 14153 6567
rect 14911 6593 14937 6599
rect 14911 6561 14937 6567
rect 7575 6537 7601 6543
rect 3257 6511 3263 6537
rect 3289 6511 3295 6537
rect 7575 6505 7601 6511
rect 1353 6455 1359 6481
rect 1385 6455 1391 6481
rect 2137 6455 2143 6481
rect 2169 6455 2175 6481
rect 3929 6455 3935 6481
rect 3961 6455 3967 6481
rect 5161 6455 5167 6481
rect 5193 6455 5199 6481
rect 5945 6455 5951 6481
rect 5977 6455 5983 6481
rect 6729 6455 6735 6481
rect 6761 6455 6767 6481
rect 9081 6455 9087 6481
rect 9113 6455 9119 6481
rect 10817 6455 10823 6481
rect 10849 6455 10855 6481
rect 10985 6455 10991 6481
rect 11017 6455 11023 6481
rect 11937 6455 11943 6481
rect 11969 6455 11975 6481
rect 12721 6455 12727 6481
rect 12753 6455 12759 6481
rect 13953 6455 13959 6481
rect 13985 6455 13991 6481
rect 14625 6455 14631 6481
rect 14657 6455 14663 6481
rect 6287 6425 6313 6431
rect 6287 6393 6313 6399
rect 8863 6425 8889 6431
rect 13455 6425 13481 6431
rect 9697 6399 9703 6425
rect 9729 6399 9735 6425
rect 10481 6399 10487 6425
rect 10513 6399 10519 6425
rect 8863 6393 8889 6399
rect 13455 6393 13481 6399
rect 336 6285 15512 6302
rect 336 6259 1903 6285
rect 1929 6259 1955 6285
rect 1981 6259 2007 6285
rect 2033 6259 11903 6285
rect 11929 6259 11955 6285
rect 11981 6259 12007 6285
rect 12033 6259 15512 6285
rect 336 6242 15512 6259
rect 1919 6201 1945 6207
rect 1919 6169 1945 6175
rect 3655 6201 3681 6207
rect 3655 6169 3681 6175
rect 5055 6201 5081 6207
rect 5055 6169 5081 6175
rect 6007 6201 6033 6207
rect 6007 6169 6033 6175
rect 10431 6201 10457 6207
rect 10431 6169 10457 6175
rect 11383 6201 11409 6207
rect 11383 6169 11409 6175
rect 11999 6201 12025 6207
rect 11999 6169 12025 6175
rect 12951 6201 12977 6207
rect 12951 6169 12977 6175
rect 14519 6201 14545 6207
rect 14519 6169 14545 6175
rect 2591 6145 2617 6151
rect 9591 6145 9617 6151
rect 4153 6119 4159 6145
rect 4185 6119 4191 6145
rect 6785 6119 6791 6145
rect 6817 6119 6823 6145
rect 9249 6119 9255 6145
rect 9281 6119 9287 6145
rect 2591 6113 2617 6119
rect 9591 6113 9617 6119
rect 10039 6145 10065 6151
rect 10039 6113 10065 6119
rect 8135 6089 8161 6095
rect 2753 6063 2759 6089
rect 2785 6063 2791 6089
rect 7233 6063 7239 6089
rect 7265 6063 7271 6089
rect 8135 6057 8161 6063
rect 8583 6089 8609 6095
rect 8583 6057 8609 6063
rect 8751 6089 8777 6095
rect 9479 6089 9505 6095
rect 8969 6063 8975 6089
rect 9001 6063 9007 6089
rect 14345 6063 14351 6089
rect 14377 6063 14383 6089
rect 8751 6057 8777 6063
rect 9479 6057 9505 6063
rect 2983 6033 3009 6039
rect 6511 6033 6537 6039
rect 2193 6007 2199 6033
rect 2225 6007 2231 6033
rect 3145 6007 3151 6033
rect 3177 6007 3183 6033
rect 4545 6007 4551 6033
rect 4577 6007 4583 6033
rect 5329 6007 5335 6033
rect 5361 6007 5367 6033
rect 5497 6007 5503 6033
rect 5529 6007 5535 6033
rect 2983 6001 3009 6007
rect 6511 6001 6537 6007
rect 7407 6033 7433 6039
rect 7407 6001 7433 6007
rect 7855 6033 7881 6039
rect 7855 6001 7881 6007
rect 8303 6033 8329 6039
rect 13735 6033 13761 6039
rect 10929 6007 10935 6033
rect 10961 6007 10967 6033
rect 11097 6007 11103 6033
rect 11129 6007 11135 6033
rect 12497 6007 12503 6033
rect 12529 6007 12535 6033
rect 12665 6007 12671 6033
rect 12697 6007 12703 6033
rect 8303 6001 8329 6007
rect 13735 6001 13761 6007
rect 15303 6033 15329 6039
rect 15303 6001 15329 6007
rect 7687 5977 7713 5983
rect 7687 5945 7713 5951
rect 9759 5977 9785 5983
rect 9759 5945 9785 5951
rect 13455 5977 13481 5983
rect 13455 5945 13481 5951
rect 13959 5977 13985 5983
rect 13959 5945 13985 5951
rect 15023 5977 15049 5983
rect 15023 5945 15049 5951
rect 336 5893 15512 5910
rect 336 5867 2233 5893
rect 2259 5867 2285 5893
rect 2311 5867 2337 5893
rect 2363 5867 12233 5893
rect 12259 5867 12285 5893
rect 12311 5867 12337 5893
rect 12363 5867 15512 5893
rect 336 5850 15512 5867
rect 2311 5809 2337 5815
rect 2311 5777 2337 5783
rect 3095 5809 3121 5815
rect 3095 5777 3121 5783
rect 4775 5809 4801 5815
rect 4775 5777 4801 5783
rect 8079 5809 8105 5815
rect 8079 5777 8105 5783
rect 8751 5809 8777 5815
rect 8751 5777 8777 5783
rect 9143 5809 9169 5815
rect 9143 5777 9169 5783
rect 9535 5809 9561 5815
rect 9535 5777 9561 5783
rect 10711 5809 10737 5815
rect 10711 5777 10737 5783
rect 11103 5809 11129 5815
rect 11103 5777 11129 5783
rect 11607 5809 11633 5815
rect 11607 5777 11633 5783
rect 14127 5809 14153 5815
rect 14127 5777 14153 5783
rect 1807 5753 1833 5759
rect 1807 5721 1833 5727
rect 4495 5753 4521 5759
rect 5161 5727 5167 5753
rect 5193 5727 5199 5753
rect 7121 5727 7127 5753
rect 7153 5727 7159 5753
rect 4495 5721 4521 5727
rect 7631 5697 7657 5703
rect 1577 5671 1583 5697
rect 1609 5671 1615 5697
rect 2529 5671 2535 5697
rect 2561 5671 2567 5697
rect 3257 5671 3263 5697
rect 3289 5671 3295 5697
rect 4153 5671 4159 5697
rect 4185 5671 4191 5697
rect 4713 5671 4719 5697
rect 4745 5671 4751 5697
rect 5553 5671 5559 5697
rect 5585 5671 5591 5697
rect 5721 5671 5727 5697
rect 5753 5671 5759 5697
rect 7631 5665 7657 5671
rect 9423 5697 9449 5703
rect 9423 5665 9449 5671
rect 9759 5697 9785 5703
rect 9759 5665 9785 5671
rect 10207 5697 10233 5703
rect 11321 5671 11327 5697
rect 11353 5671 11359 5697
rect 12273 5671 12279 5697
rect 12305 5671 12311 5697
rect 13057 5671 13063 5697
rect 13089 5671 13095 5697
rect 13897 5671 13903 5697
rect 13929 5671 13935 5697
rect 14681 5671 14687 5697
rect 14713 5671 14719 5697
rect 10207 5665 10233 5671
rect 1415 5641 1441 5647
rect 1415 5609 1441 5615
rect 3879 5641 3905 5647
rect 6623 5641 6649 5647
rect 6057 5615 6063 5641
rect 6089 5615 6095 5641
rect 3879 5609 3905 5615
rect 6623 5609 6649 5615
rect 7463 5641 7489 5647
rect 7463 5609 7489 5615
rect 7911 5641 7937 5647
rect 7911 5609 7937 5615
rect 9647 5641 9673 5647
rect 9647 5609 9673 5615
rect 10039 5641 10065 5647
rect 10039 5609 10065 5615
rect 10487 5641 10513 5647
rect 12559 5641 12585 5647
rect 10929 5615 10935 5641
rect 10961 5615 10967 5641
rect 10487 5609 10513 5615
rect 12559 5609 12585 5615
rect 13567 5641 13593 5647
rect 13567 5609 13593 5615
rect 15191 5585 15217 5591
rect 15191 5553 15217 5559
rect 336 5501 15512 5518
rect 336 5475 1903 5501
rect 1929 5475 1955 5501
rect 1981 5475 2007 5501
rect 2033 5475 11903 5501
rect 11929 5475 11955 5501
rect 11981 5475 12007 5501
rect 12033 5475 15512 5501
rect 336 5458 15512 5475
rect 3487 5417 3513 5423
rect 3487 5385 3513 5391
rect 5055 5417 5081 5423
rect 5055 5385 5081 5391
rect 6511 5417 6537 5423
rect 6511 5385 6537 5391
rect 11831 5417 11857 5423
rect 11831 5385 11857 5391
rect 12615 5417 12641 5423
rect 12615 5385 12641 5391
rect 2591 5361 2617 5367
rect 1801 5335 1807 5361
rect 1833 5335 1839 5361
rect 2591 5329 2617 5335
rect 2983 5361 3009 5367
rect 8807 5361 8833 5367
rect 13847 5361 13873 5367
rect 4209 5335 4215 5361
rect 4241 5335 4247 5361
rect 5777 5335 5783 5361
rect 5809 5335 5815 5361
rect 8353 5335 8359 5361
rect 8385 5335 8391 5361
rect 9809 5335 9815 5361
rect 9841 5335 9847 5361
rect 10873 5335 10879 5361
rect 10905 5335 10911 5361
rect 11321 5335 11327 5361
rect 11353 5335 11359 5361
rect 13505 5335 13511 5361
rect 13537 5335 13543 5361
rect 2983 5329 3009 5335
rect 8807 5329 8833 5335
rect 13847 5329 13873 5335
rect 9087 5305 9113 5311
rect 2137 5279 2143 5305
rect 2169 5279 2175 5305
rect 2753 5279 2759 5305
rect 2785 5279 2791 5305
rect 3761 5279 3767 5305
rect 3793 5279 3799 5305
rect 4545 5279 4551 5305
rect 4577 5279 4583 5305
rect 5329 5279 5335 5305
rect 5361 5279 5367 5305
rect 7009 5279 7015 5305
rect 7041 5279 7047 5305
rect 7401 5279 7407 5305
rect 7433 5279 7439 5305
rect 9087 5273 9113 5279
rect 9535 5305 9561 5311
rect 10655 5305 10681 5311
rect 14239 5305 14265 5311
rect 9977 5279 9983 5305
rect 10009 5279 10015 5305
rect 11153 5279 11159 5305
rect 11185 5279 11191 5305
rect 11545 5279 11551 5305
rect 11577 5279 11583 5305
rect 13225 5279 13231 5305
rect 13257 5279 13263 5305
rect 14737 5279 14743 5305
rect 14769 5279 14775 5305
rect 9535 5273 9561 5279
rect 10655 5273 10681 5279
rect 14239 5273 14265 5279
rect 7183 5249 7209 5255
rect 6113 5223 6119 5249
rect 6145 5223 6151 5249
rect 7183 5217 7209 5223
rect 7967 5249 7993 5255
rect 7967 5217 7993 5223
rect 9255 5249 9281 5255
rect 14519 5249 14545 5255
rect 10481 5223 10487 5249
rect 10513 5223 10519 5249
rect 12329 5223 12335 5249
rect 12361 5223 12367 5249
rect 15073 5223 15079 5249
rect 15105 5223 15111 5249
rect 9255 5217 9281 5223
rect 14519 5217 14545 5223
rect 7687 5193 7713 5199
rect 7687 5161 7713 5167
rect 8135 5193 8161 5199
rect 8135 5161 8161 5167
rect 10319 5193 10345 5199
rect 10319 5161 10345 5167
rect 14015 5193 14041 5199
rect 14015 5161 14041 5167
rect 336 5109 15512 5126
rect 336 5083 2233 5109
rect 2259 5083 2285 5109
rect 2311 5083 2337 5109
rect 2363 5083 12233 5109
rect 12259 5083 12285 5109
rect 12311 5083 12337 5109
rect 12363 5083 15512 5109
rect 336 5066 15512 5083
rect 3095 5025 3121 5031
rect 3095 4993 3121 4999
rect 3879 5025 3905 5031
rect 3879 4993 3905 4999
rect 4607 5025 4633 5031
rect 4607 4993 4633 4999
rect 7183 5025 7209 5031
rect 7183 4993 7209 4999
rect 7351 5025 7377 5031
rect 7351 4993 7377 4999
rect 7631 5025 7657 5031
rect 7631 4993 7657 4999
rect 9255 5025 9281 5031
rect 9255 4993 9281 4999
rect 9703 5025 9729 5031
rect 9703 4993 9729 4999
rect 10151 5025 10177 5031
rect 10151 4993 10177 4999
rect 10319 5025 10345 5031
rect 10319 4993 10345 4999
rect 10431 5025 10457 5031
rect 10431 4993 10457 4999
rect 10543 5025 10569 5031
rect 10543 4993 10569 4999
rect 10991 5025 11017 5031
rect 10991 4993 11017 4999
rect 11551 5025 11577 5031
rect 11551 4993 11577 4999
rect 12559 5025 12585 5031
rect 12559 4993 12585 4999
rect 6455 4969 6481 4975
rect 4153 4943 4159 4969
rect 4185 4943 4191 4969
rect 4937 4943 4943 4969
rect 4969 4943 4975 4969
rect 14289 4943 14295 4969
rect 14321 4943 14327 4969
rect 14681 4943 14687 4969
rect 14713 4943 14719 4969
rect 6455 4937 6481 4943
rect 11383 4913 11409 4919
rect 2025 4887 2031 4913
rect 2057 4887 2063 4913
rect 3313 4887 3319 4913
rect 3345 4887 3351 4913
rect 5329 4887 5335 4913
rect 5361 4887 5367 4913
rect 6113 4887 6119 4913
rect 6145 4887 6151 4913
rect 6673 4887 6679 4913
rect 6705 4887 6711 4913
rect 12273 4887 12279 4913
rect 12305 4887 12311 4913
rect 13561 4887 13567 4913
rect 13593 4887 13599 4913
rect 13897 4887 13903 4913
rect 13929 4887 13935 4913
rect 11383 4881 11409 4887
rect 5615 4857 5641 4863
rect 2417 4831 2423 4857
rect 2449 4831 2455 4857
rect 5615 4825 5641 4831
rect 6903 4857 6929 4863
rect 6903 4825 6929 4831
rect 7463 4857 7489 4863
rect 7463 4825 7489 4831
rect 7967 4857 7993 4863
rect 11831 4857 11857 4863
rect 10761 4831 10767 4857
rect 10793 4831 10799 4857
rect 11153 4831 11159 4857
rect 11185 4831 11191 4857
rect 7967 4825 7993 4831
rect 11831 4825 11857 4831
rect 11943 4857 11969 4863
rect 11943 4825 11969 4831
rect 13175 4857 13201 4863
rect 13175 4825 13201 4831
rect 15191 4801 15217 4807
rect 15191 4769 15217 4775
rect 336 4717 15512 4734
rect 336 4691 1903 4717
rect 1929 4691 1955 4717
rect 1981 4691 2007 4717
rect 2033 4691 11903 4717
rect 11929 4691 11955 4717
rect 11981 4691 12007 4717
rect 12033 4691 15512 4717
rect 336 4674 15512 4691
rect 3711 4633 3737 4639
rect 3711 4601 3737 4607
rect 5223 4633 5249 4639
rect 5223 4601 5249 4607
rect 12671 4633 12697 4639
rect 12671 4601 12697 4607
rect 13455 4633 13481 4639
rect 13455 4601 13481 4607
rect 2423 4577 2449 4583
rect 6119 4577 6145 4583
rect 2921 4551 2927 4577
rect 2953 4551 2959 4577
rect 4321 4551 4327 4577
rect 4353 4551 4359 4577
rect 2423 4545 2449 4551
rect 6119 4545 6145 4551
rect 6903 4577 6929 4583
rect 6903 4545 6929 4551
rect 11271 4577 11297 4583
rect 11271 4545 11297 4551
rect 11775 4577 11801 4583
rect 14519 4577 14545 4583
rect 12161 4551 12167 4577
rect 12193 4551 12199 4577
rect 11775 4545 11801 4551
rect 14519 4545 14545 4551
rect 2143 4521 2169 4527
rect 6007 4521 6033 4527
rect 4769 4495 4775 4521
rect 4801 4495 4807 4521
rect 11993 4495 11999 4521
rect 12025 4495 12031 4521
rect 13057 4495 13063 4521
rect 13089 4495 13095 4521
rect 14289 4495 14295 4521
rect 14321 4495 14327 4521
rect 2143 4489 2169 4495
rect 6007 4489 6033 4495
rect 1863 4465 1889 4471
rect 5727 4465 5753 4471
rect 2585 4439 2591 4465
rect 2617 4439 2623 4465
rect 3985 4439 3991 4465
rect 4017 4439 4023 4465
rect 4937 4439 4943 4465
rect 4969 4439 4975 4465
rect 1863 4433 1889 4439
rect 5727 4433 5753 4439
rect 7855 4465 7881 4471
rect 7855 4433 7881 4439
rect 8471 4465 8497 4471
rect 13953 4439 13959 4465
rect 13985 4439 13991 4465
rect 14681 4439 14687 4465
rect 14713 4439 14719 4465
rect 15073 4439 15079 4465
rect 15105 4439 15111 4465
rect 8471 4433 8497 4439
rect 7407 4409 7433 4415
rect 7407 4377 7433 4383
rect 7575 4409 7601 4415
rect 7575 4377 7601 4383
rect 8079 4409 8105 4415
rect 8079 4377 8105 4383
rect 8191 4409 8217 4415
rect 8191 4377 8217 4383
rect 11327 4409 11353 4415
rect 11327 4377 11353 4383
rect 11495 4409 11521 4415
rect 11495 4377 11521 4383
rect 11943 4409 11969 4415
rect 11943 4377 11969 4383
rect 14239 4409 14265 4415
rect 14239 4377 14265 4383
rect 336 4325 15512 4342
rect 336 4299 2233 4325
rect 2259 4299 2285 4325
rect 2311 4299 2337 4325
rect 2363 4299 12233 4325
rect 12259 4299 12285 4325
rect 12311 4299 12337 4325
rect 12363 4299 15512 4325
rect 336 4282 15512 4299
rect 11831 4241 11857 4247
rect 11831 4209 11857 4215
rect 2311 4185 2337 4191
rect 4439 4185 4465 4191
rect 4153 4159 4159 4185
rect 4185 4159 4191 4185
rect 2311 4153 2337 4159
rect 4439 4153 4465 4159
rect 4719 4185 4745 4191
rect 4719 4153 4745 4159
rect 4887 4185 4913 4191
rect 4887 4153 4913 4159
rect 5279 4185 5305 4191
rect 5279 4153 5305 4159
rect 5503 4185 5529 4191
rect 5503 4153 5529 4159
rect 5951 4185 5977 4191
rect 5951 4153 5977 4159
rect 6231 4185 6257 4191
rect 6231 4153 6257 4159
rect 6399 4185 6425 4191
rect 12721 4159 12727 4185
rect 12753 4159 12759 4185
rect 6399 4153 6425 4159
rect 2591 4129 2617 4135
rect 5783 4129 5809 4135
rect 3369 4103 3375 4129
rect 3401 4103 3407 4129
rect 2591 4097 2617 4103
rect 5783 4097 5809 4103
rect 7799 4129 7825 4135
rect 12441 4103 12447 4129
rect 12473 4103 12479 4129
rect 13225 4103 13231 4129
rect 13257 4103 13263 4129
rect 14009 4103 14015 4129
rect 14041 4103 14047 4129
rect 14681 4103 14687 4129
rect 14713 4103 14719 4129
rect 7799 4097 7825 4103
rect 7631 4073 7657 4079
rect 2921 4047 2927 4073
rect 2953 4047 2959 4073
rect 3817 4047 3823 4073
rect 3849 4047 3855 4073
rect 5049 4047 5055 4073
rect 5081 4047 5087 4073
rect 7631 4041 7657 4047
rect 8079 4073 8105 4079
rect 8079 4041 8105 4047
rect 13623 4073 13649 4079
rect 13623 4041 13649 4047
rect 14407 4073 14433 4079
rect 14407 4041 14433 4047
rect 15191 4017 15217 4023
rect 15191 3985 15217 3991
rect 336 3933 15512 3950
rect 336 3907 1903 3933
rect 1929 3907 1955 3933
rect 1981 3907 2007 3933
rect 2033 3907 11903 3933
rect 11929 3907 11955 3933
rect 11981 3907 12007 3933
rect 12033 3907 15512 3933
rect 336 3890 15512 3907
rect 2759 3793 2785 3799
rect 2759 3761 2785 3767
rect 3431 3793 3457 3799
rect 5167 3793 5193 3799
rect 4097 3767 4103 3793
rect 4129 3767 4135 3793
rect 3431 3761 3457 3767
rect 5167 3761 5193 3767
rect 5615 3793 5641 3799
rect 5615 3761 5641 3767
rect 5671 3793 5697 3799
rect 5671 3761 5697 3767
rect 5951 3793 5977 3799
rect 5951 3761 5977 3767
rect 8079 3793 8105 3799
rect 12833 3767 12839 3793
rect 12865 3767 12871 3793
rect 13673 3767 13679 3793
rect 13705 3767 13711 3793
rect 15129 3767 15135 3793
rect 15161 3767 15167 3793
rect 8079 3761 8105 3767
rect 3711 3737 3737 3743
rect 3711 3705 3737 3711
rect 3823 3737 3849 3743
rect 3823 3705 3849 3711
rect 7799 3737 7825 3743
rect 13113 3711 13119 3737
rect 13145 3711 13151 3737
rect 14681 3711 14687 3737
rect 14713 3711 14719 3737
rect 7799 3705 7825 3711
rect 4327 3681 4353 3687
rect 4327 3649 4353 3655
rect 4439 3681 4465 3687
rect 4439 3649 4465 3655
rect 5447 3681 5473 3687
rect 5447 3649 5473 3655
rect 7631 3681 7657 3687
rect 13337 3655 13343 3681
rect 13369 3655 13375 3681
rect 7631 3649 7657 3655
rect 7239 3625 7265 3631
rect 7239 3593 7265 3599
rect 7351 3625 7377 3631
rect 7351 3593 7377 3599
rect 336 3541 15512 3558
rect 336 3515 2233 3541
rect 2259 3515 2285 3541
rect 2311 3515 2337 3541
rect 2363 3515 12233 3541
rect 12259 3515 12285 3541
rect 12311 3515 12337 3541
rect 12363 3515 15512 3541
rect 336 3498 15512 3515
rect 7687 3457 7713 3463
rect 7687 3425 7713 3431
rect 13113 3375 13119 3401
rect 13145 3375 13151 3401
rect 14681 3375 14687 3401
rect 14713 3375 14719 3401
rect 3879 3345 3905 3351
rect 3879 3313 3905 3319
rect 4159 3345 4185 3351
rect 4159 3313 4185 3319
rect 4439 3345 4465 3351
rect 4439 3313 4465 3319
rect 7183 3345 7209 3351
rect 7183 3313 7209 3319
rect 8359 3345 8385 3351
rect 13897 3319 13903 3345
rect 13929 3319 13935 3345
rect 8359 3313 8385 3319
rect 7015 3289 7041 3295
rect 7015 3257 7041 3263
rect 7463 3289 7489 3295
rect 7463 3257 7489 3263
rect 8079 3289 8105 3295
rect 8079 3257 8105 3263
rect 8639 3289 8665 3295
rect 8639 3257 8665 3263
rect 13623 3289 13649 3295
rect 13623 3257 13649 3263
rect 15191 3289 15217 3295
rect 15191 3257 15217 3263
rect 14407 3233 14433 3239
rect 14407 3201 14433 3207
rect 336 3149 15512 3166
rect 336 3123 1903 3149
rect 1929 3123 1955 3149
rect 1981 3123 2007 3149
rect 2033 3123 11903 3149
rect 11929 3123 11955 3149
rect 11981 3123 12007 3149
rect 12033 3123 15512 3149
rect 336 3106 15512 3123
rect 7519 3009 7545 3015
rect 15129 2983 15135 3009
rect 15161 2983 15167 3009
rect 7519 2977 7545 2983
rect 14737 2927 14743 2953
rect 14769 2927 14775 2953
rect 7071 2841 7097 2847
rect 7071 2809 7097 2815
rect 7239 2841 7265 2847
rect 7239 2809 7265 2815
rect 336 2757 15512 2774
rect 336 2731 2233 2757
rect 2259 2731 2285 2757
rect 2311 2731 2337 2757
rect 2363 2731 12233 2757
rect 12259 2731 12285 2757
rect 12311 2731 12337 2757
rect 12363 2731 15512 2757
rect 336 2714 15512 2731
rect 7239 2673 7265 2679
rect 7239 2641 7265 2647
rect 8863 2673 8889 2679
rect 8863 2641 8889 2647
rect 8079 2617 8105 2623
rect 8079 2585 8105 2591
rect 8695 2617 8721 2623
rect 8695 2585 8721 2591
rect 9143 2617 9169 2623
rect 13897 2591 13903 2617
rect 13929 2591 13935 2617
rect 15073 2591 15079 2617
rect 15105 2591 15111 2617
rect 9143 2585 9169 2591
rect 6623 2561 6649 2567
rect 6623 2529 6649 2535
rect 6791 2561 6817 2567
rect 6791 2529 6817 2535
rect 7519 2561 7545 2567
rect 7519 2529 7545 2535
rect 7631 2561 7657 2567
rect 7631 2529 7657 2535
rect 7799 2561 7825 2567
rect 7799 2529 7825 2535
rect 8415 2561 8441 2567
rect 14681 2535 14687 2561
rect 14713 2535 14719 2561
rect 8415 2529 8441 2535
rect 7071 2505 7097 2511
rect 7071 2473 7097 2479
rect 14407 2505 14433 2511
rect 14407 2473 14433 2479
rect 336 2365 15512 2382
rect 336 2339 1903 2365
rect 1929 2339 1955 2365
rect 1981 2339 2007 2365
rect 2033 2339 11903 2365
rect 11929 2339 11955 2365
rect 11981 2339 12007 2365
rect 12033 2339 15512 2365
rect 336 2322 15512 2339
rect 7127 2225 7153 2231
rect 8135 2225 8161 2231
rect 7513 2199 7519 2225
rect 7545 2199 7551 2225
rect 7127 2193 7153 2199
rect 8135 2193 8161 2199
rect 8751 2225 8777 2231
rect 15129 2199 15135 2225
rect 15161 2199 15167 2225
rect 8751 2193 8777 2199
rect 8303 2169 8329 2175
rect 14681 2143 14687 2169
rect 14713 2143 14719 2169
rect 8303 2137 8329 2143
rect 7015 2057 7041 2063
rect 7015 2025 7041 2031
rect 7295 2057 7321 2063
rect 7295 2025 7321 2031
rect 7687 2057 7713 2063
rect 7687 2025 7713 2031
rect 7855 2057 7881 2063
rect 7855 2025 7881 2031
rect 14575 2057 14601 2063
rect 14575 2025 14601 2031
rect 336 1973 15512 1990
rect 336 1947 2233 1973
rect 2259 1947 2285 1973
rect 2311 1947 2337 1973
rect 2363 1947 12233 1973
rect 12259 1947 12285 1973
rect 12311 1947 12337 1973
rect 12363 1947 15512 1973
rect 336 1930 15512 1947
rect 13567 1833 13593 1839
rect 13897 1807 13903 1833
rect 13929 1807 13935 1833
rect 14289 1807 14295 1833
rect 14321 1807 14327 1833
rect 13567 1801 13593 1807
rect 6959 1777 6985 1783
rect 6959 1745 6985 1751
rect 13287 1777 13313 1783
rect 13287 1745 13313 1751
rect 13679 1777 13705 1783
rect 14737 1751 14743 1777
rect 14769 1751 14775 1777
rect 13679 1745 13705 1751
rect 6791 1721 6817 1727
rect 6791 1689 6817 1695
rect 7239 1721 7265 1727
rect 7239 1689 7265 1695
rect 8023 1721 8049 1727
rect 8023 1689 8049 1695
rect 15191 1721 15217 1727
rect 15191 1689 15217 1695
rect 336 1581 15512 1598
rect 336 1555 1903 1581
rect 1929 1555 1955 1581
rect 1981 1555 2007 1581
rect 2033 1555 11903 1581
rect 11929 1555 11955 1581
rect 11981 1555 12007 1581
rect 12033 1555 15512 1581
rect 336 1538 15512 1555
rect 6847 1441 6873 1447
rect 6847 1409 6873 1415
rect 7295 1441 7321 1447
rect 8919 1441 8945 1447
rect 8353 1415 8359 1441
rect 8385 1415 8391 1441
rect 7295 1409 7321 1415
rect 8919 1409 8945 1415
rect 12055 1441 12081 1447
rect 12945 1415 12951 1441
rect 12977 1415 12983 1441
rect 14289 1415 14295 1441
rect 14321 1415 14327 1441
rect 15129 1415 15135 1441
rect 15161 1415 15167 1441
rect 12055 1409 12081 1415
rect 7015 1385 7041 1391
rect 7015 1353 7041 1359
rect 7519 1385 7545 1391
rect 7519 1353 7545 1359
rect 7687 1385 7713 1391
rect 7687 1353 7713 1359
rect 8639 1385 8665 1391
rect 14681 1359 14687 1385
rect 14713 1359 14719 1385
rect 8639 1353 8665 1359
rect 7967 1329 7993 1335
rect 13337 1303 13343 1329
rect 13369 1303 13375 1329
rect 13729 1303 13735 1329
rect 13761 1303 13767 1329
rect 7967 1297 7993 1303
rect 8135 1273 8161 1279
rect 8135 1241 8161 1247
rect 10711 1273 10737 1279
rect 10711 1241 10737 1247
rect 11663 1273 11689 1279
rect 11663 1241 11689 1247
rect 11775 1273 11801 1279
rect 11775 1241 11801 1247
rect 12615 1273 12641 1279
rect 12615 1241 12641 1247
rect 12727 1273 12753 1279
rect 12727 1241 12753 1247
rect 14519 1273 14545 1279
rect 14519 1241 14545 1247
rect 336 1189 15512 1206
rect 336 1163 2233 1189
rect 2259 1163 2285 1189
rect 2311 1163 2337 1189
rect 2363 1163 12233 1189
rect 12259 1163 12285 1189
rect 12311 1163 12337 1189
rect 12363 1163 15512 1189
rect 336 1146 15512 1163
rect 8527 1105 8553 1111
rect 8527 1073 8553 1079
rect 7407 1049 7433 1055
rect 7407 1017 7433 1023
rect 8079 1049 8105 1055
rect 8079 1017 8105 1023
rect 9591 1049 9617 1055
rect 9591 1017 9617 1023
rect 10655 1049 10681 1055
rect 10655 1017 10681 1023
rect 11103 1049 11129 1055
rect 11103 1017 11129 1023
rect 12839 1049 12865 1055
rect 13113 1023 13119 1049
rect 13145 1023 13151 1049
rect 13897 1023 13903 1049
rect 13929 1023 13935 1049
rect 15073 1023 15079 1049
rect 15105 1023 15111 1049
rect 12839 1017 12865 1023
rect 6959 993 6985 999
rect 6959 961 6985 967
rect 7127 993 7153 999
rect 7127 961 7153 967
rect 7799 993 7825 999
rect 7799 961 7825 967
rect 9311 993 9337 999
rect 9311 961 9337 967
rect 9815 993 9841 999
rect 9815 961 9841 967
rect 10207 993 10233 999
rect 10207 961 10233 967
rect 10375 993 10401 999
rect 10375 961 10401 967
rect 10823 993 10849 999
rect 10823 961 10849 967
rect 11327 993 11353 999
rect 11327 961 11353 967
rect 12559 993 12585 999
rect 14737 967 14743 993
rect 14769 967 14775 993
rect 12559 961 12585 967
rect 7631 937 7657 943
rect 6729 911 6735 937
rect 6761 911 6767 937
rect 7631 905 7657 911
rect 9143 937 9169 943
rect 12391 937 12417 943
rect 10033 911 10039 937
rect 10065 911 10071 937
rect 11545 911 11551 937
rect 11577 911 11583 937
rect 9143 905 9169 911
rect 12391 905 12417 911
rect 14407 937 14433 943
rect 14407 905 14433 911
rect 13623 881 13649 887
rect 13623 849 13649 855
rect 336 797 15512 814
rect 336 771 1903 797
rect 1929 771 1955 797
rect 1981 771 2007 797
rect 2033 771 11903 797
rect 11929 771 11955 797
rect 11981 771 12007 797
rect 12033 771 15512 797
rect 336 754 15512 771
rect 15191 713 15217 719
rect 15191 681 15217 687
rect 7071 657 7097 663
rect 8527 657 8553 663
rect 5553 631 5559 657
rect 5585 631 5591 657
rect 6337 631 6343 657
rect 6369 631 6375 657
rect 8353 631 8359 657
rect 8385 631 8391 657
rect 7071 625 7097 631
rect 8527 625 8553 631
rect 9199 657 9225 663
rect 9199 625 9225 631
rect 10823 657 10849 663
rect 11601 631 11607 657
rect 11633 631 11639 657
rect 14345 631 14351 657
rect 14377 631 14383 657
rect 10823 625 10849 631
rect 7855 601 7881 607
rect 6505 575 6511 601
rect 6537 575 6543 601
rect 12161 575 12167 601
rect 12193 575 12199 601
rect 13897 575 13903 601
rect 13929 575 13935 601
rect 14681 575 14687 601
rect 14713 575 14719 601
rect 7855 569 7881 575
rect 8135 545 8161 551
rect 10201 519 10207 545
rect 10233 519 10239 545
rect 12945 519 12951 545
rect 12977 519 12983 545
rect 13337 519 13343 545
rect 13369 519 13375 545
rect 8135 513 8161 519
rect 5783 489 5809 495
rect 5783 457 5809 463
rect 5895 489 5921 495
rect 5895 457 5921 463
rect 6679 489 6705 495
rect 6679 457 6705 463
rect 6959 489 6985 495
rect 6959 457 6985 463
rect 7463 489 7489 495
rect 7463 457 7489 463
rect 7575 489 7601 495
rect 7575 457 7601 463
rect 8807 489 8833 495
rect 8807 457 8833 463
rect 8919 489 8945 495
rect 8919 457 8945 463
rect 9647 489 9673 495
rect 9647 457 9673 463
rect 9815 489 9841 495
rect 9815 457 9841 463
rect 10039 489 10065 495
rect 10039 457 10065 463
rect 10431 489 10457 495
rect 10431 457 10457 463
rect 10543 489 10569 495
rect 10543 457 10569 463
rect 11103 489 11129 495
rect 11103 457 11129 463
rect 11159 489 11185 495
rect 11159 457 11185 463
rect 11383 489 11409 495
rect 11383 457 11409 463
rect 12447 489 12473 495
rect 12447 457 12473 463
rect 336 405 15512 422
rect 336 379 2233 405
rect 2259 379 2285 405
rect 2311 379 2337 405
rect 2363 379 12233 405
rect 12259 379 12285 405
rect 12311 379 12337 405
rect 12363 379 15512 405
rect 336 362 15512 379
<< via1 >>
rect 2233 6651 2259 6677
rect 2285 6651 2311 6677
rect 2337 6651 2363 6677
rect 12233 6651 12259 6677
rect 12285 6651 12311 6677
rect 12337 6651 12363 6677
rect 1079 6567 1105 6593
rect 1863 6567 1889 6593
rect 2983 6567 3009 6593
rect 3767 6567 3793 6593
rect 4887 6567 4913 6593
rect 5671 6567 5697 6593
rect 6567 6567 6593 6593
rect 7015 6567 7041 6593
rect 7855 6567 7881 6593
rect 8135 6567 8161 6593
rect 8247 6567 8273 6593
rect 8751 6567 8777 6593
rect 9255 6567 9281 6593
rect 9479 6567 9505 6593
rect 11271 6567 11297 6593
rect 12223 6567 12249 6593
rect 13007 6567 13033 6593
rect 14127 6567 14153 6593
rect 14911 6567 14937 6593
rect 3263 6511 3289 6537
rect 7575 6511 7601 6537
rect 1359 6455 1385 6481
rect 2143 6455 2169 6481
rect 3935 6455 3961 6481
rect 5167 6455 5193 6481
rect 5951 6455 5977 6481
rect 6735 6455 6761 6481
rect 9087 6455 9113 6481
rect 10823 6455 10849 6481
rect 10991 6455 11017 6481
rect 11943 6455 11969 6481
rect 12727 6455 12753 6481
rect 13959 6455 13985 6481
rect 14631 6455 14657 6481
rect 6287 6399 6313 6425
rect 8863 6399 8889 6425
rect 9703 6399 9729 6425
rect 10487 6399 10513 6425
rect 13455 6399 13481 6425
rect 1903 6259 1929 6285
rect 1955 6259 1981 6285
rect 2007 6259 2033 6285
rect 11903 6259 11929 6285
rect 11955 6259 11981 6285
rect 12007 6259 12033 6285
rect 1919 6175 1945 6201
rect 3655 6175 3681 6201
rect 5055 6175 5081 6201
rect 6007 6175 6033 6201
rect 10431 6175 10457 6201
rect 11383 6175 11409 6201
rect 11999 6175 12025 6201
rect 12951 6175 12977 6201
rect 14519 6175 14545 6201
rect 2591 6119 2617 6145
rect 4159 6119 4185 6145
rect 6791 6119 6817 6145
rect 9255 6119 9281 6145
rect 9591 6119 9617 6145
rect 10039 6119 10065 6145
rect 2759 6063 2785 6089
rect 7239 6063 7265 6089
rect 8135 6063 8161 6089
rect 8583 6063 8609 6089
rect 8751 6063 8777 6089
rect 8975 6063 9001 6089
rect 9479 6063 9505 6089
rect 14351 6063 14377 6089
rect 2199 6007 2225 6033
rect 2983 6007 3009 6033
rect 3151 6007 3177 6033
rect 4551 6007 4577 6033
rect 5335 6007 5361 6033
rect 5503 6007 5529 6033
rect 6511 6007 6537 6033
rect 7407 6007 7433 6033
rect 7855 6007 7881 6033
rect 8303 6007 8329 6033
rect 10935 6007 10961 6033
rect 11103 6007 11129 6033
rect 12503 6007 12529 6033
rect 12671 6007 12697 6033
rect 13735 6007 13761 6033
rect 15303 6007 15329 6033
rect 7687 5951 7713 5977
rect 9759 5951 9785 5977
rect 13455 5951 13481 5977
rect 13959 5951 13985 5977
rect 15023 5951 15049 5977
rect 2233 5867 2259 5893
rect 2285 5867 2311 5893
rect 2337 5867 2363 5893
rect 12233 5867 12259 5893
rect 12285 5867 12311 5893
rect 12337 5867 12363 5893
rect 2311 5783 2337 5809
rect 3095 5783 3121 5809
rect 4775 5783 4801 5809
rect 8079 5783 8105 5809
rect 8751 5783 8777 5809
rect 9143 5783 9169 5809
rect 9535 5783 9561 5809
rect 10711 5783 10737 5809
rect 11103 5783 11129 5809
rect 11607 5783 11633 5809
rect 14127 5783 14153 5809
rect 1807 5727 1833 5753
rect 4495 5727 4521 5753
rect 5167 5727 5193 5753
rect 7127 5727 7153 5753
rect 1583 5671 1609 5697
rect 2535 5671 2561 5697
rect 3263 5671 3289 5697
rect 4159 5671 4185 5697
rect 4719 5671 4745 5697
rect 5559 5671 5585 5697
rect 5727 5671 5753 5697
rect 7631 5671 7657 5697
rect 9423 5671 9449 5697
rect 9759 5671 9785 5697
rect 10207 5671 10233 5697
rect 11327 5671 11353 5697
rect 12279 5671 12305 5697
rect 13063 5671 13089 5697
rect 13903 5671 13929 5697
rect 14687 5671 14713 5697
rect 1415 5615 1441 5641
rect 3879 5615 3905 5641
rect 6063 5615 6089 5641
rect 6623 5615 6649 5641
rect 7463 5615 7489 5641
rect 7911 5615 7937 5641
rect 9647 5615 9673 5641
rect 10039 5615 10065 5641
rect 10487 5615 10513 5641
rect 10935 5615 10961 5641
rect 12559 5615 12585 5641
rect 13567 5615 13593 5641
rect 15191 5559 15217 5585
rect 1903 5475 1929 5501
rect 1955 5475 1981 5501
rect 2007 5475 2033 5501
rect 11903 5475 11929 5501
rect 11955 5475 11981 5501
rect 12007 5475 12033 5501
rect 3487 5391 3513 5417
rect 5055 5391 5081 5417
rect 6511 5391 6537 5417
rect 11831 5391 11857 5417
rect 12615 5391 12641 5417
rect 1807 5335 1833 5361
rect 2591 5335 2617 5361
rect 2983 5335 3009 5361
rect 4215 5335 4241 5361
rect 5783 5335 5809 5361
rect 8359 5335 8385 5361
rect 8807 5335 8833 5361
rect 9815 5335 9841 5361
rect 10879 5335 10905 5361
rect 11327 5335 11353 5361
rect 13511 5335 13537 5361
rect 13847 5335 13873 5361
rect 2143 5279 2169 5305
rect 2759 5279 2785 5305
rect 3767 5279 3793 5305
rect 4551 5279 4577 5305
rect 5335 5279 5361 5305
rect 7015 5279 7041 5305
rect 7407 5279 7433 5305
rect 9087 5279 9113 5305
rect 9535 5279 9561 5305
rect 9983 5279 10009 5305
rect 10655 5279 10681 5305
rect 11159 5279 11185 5305
rect 11551 5279 11577 5305
rect 13231 5279 13257 5305
rect 14239 5279 14265 5305
rect 14743 5279 14769 5305
rect 6119 5223 6145 5249
rect 7183 5223 7209 5249
rect 7967 5223 7993 5249
rect 9255 5223 9281 5249
rect 10487 5223 10513 5249
rect 12335 5223 12361 5249
rect 14519 5223 14545 5249
rect 15079 5223 15105 5249
rect 7687 5167 7713 5193
rect 8135 5167 8161 5193
rect 10319 5167 10345 5193
rect 14015 5167 14041 5193
rect 2233 5083 2259 5109
rect 2285 5083 2311 5109
rect 2337 5083 2363 5109
rect 12233 5083 12259 5109
rect 12285 5083 12311 5109
rect 12337 5083 12363 5109
rect 3095 4999 3121 5025
rect 3879 4999 3905 5025
rect 4607 4999 4633 5025
rect 7183 4999 7209 5025
rect 7351 4999 7377 5025
rect 7631 4999 7657 5025
rect 9255 4999 9281 5025
rect 9703 4999 9729 5025
rect 10151 4999 10177 5025
rect 10319 4999 10345 5025
rect 10431 4999 10457 5025
rect 10543 4999 10569 5025
rect 10991 4999 11017 5025
rect 11551 4999 11577 5025
rect 12559 4999 12585 5025
rect 4159 4943 4185 4969
rect 4943 4943 4969 4969
rect 6455 4943 6481 4969
rect 14295 4943 14321 4969
rect 14687 4943 14713 4969
rect 2031 4887 2057 4913
rect 3319 4887 3345 4913
rect 5335 4887 5361 4913
rect 6119 4887 6145 4913
rect 6679 4887 6705 4913
rect 11383 4887 11409 4913
rect 12279 4887 12305 4913
rect 13567 4887 13593 4913
rect 13903 4887 13929 4913
rect 2423 4831 2449 4857
rect 5615 4831 5641 4857
rect 6903 4831 6929 4857
rect 7463 4831 7489 4857
rect 7967 4831 7993 4857
rect 10767 4831 10793 4857
rect 11159 4831 11185 4857
rect 11831 4831 11857 4857
rect 11943 4831 11969 4857
rect 13175 4831 13201 4857
rect 15191 4775 15217 4801
rect 1903 4691 1929 4717
rect 1955 4691 1981 4717
rect 2007 4691 2033 4717
rect 11903 4691 11929 4717
rect 11955 4691 11981 4717
rect 12007 4691 12033 4717
rect 3711 4607 3737 4633
rect 5223 4607 5249 4633
rect 12671 4607 12697 4633
rect 13455 4607 13481 4633
rect 2423 4551 2449 4577
rect 2927 4551 2953 4577
rect 4327 4551 4353 4577
rect 6119 4551 6145 4577
rect 6903 4551 6929 4577
rect 11271 4551 11297 4577
rect 11775 4551 11801 4577
rect 12167 4551 12193 4577
rect 14519 4551 14545 4577
rect 2143 4495 2169 4521
rect 4775 4495 4801 4521
rect 6007 4495 6033 4521
rect 11999 4495 12025 4521
rect 13063 4495 13089 4521
rect 14295 4495 14321 4521
rect 1863 4439 1889 4465
rect 2591 4439 2617 4465
rect 3991 4439 4017 4465
rect 4943 4439 4969 4465
rect 5727 4439 5753 4465
rect 7855 4439 7881 4465
rect 8471 4439 8497 4465
rect 13959 4439 13985 4465
rect 14687 4439 14713 4465
rect 15079 4439 15105 4465
rect 7407 4383 7433 4409
rect 7575 4383 7601 4409
rect 8079 4383 8105 4409
rect 8191 4383 8217 4409
rect 11327 4383 11353 4409
rect 11495 4383 11521 4409
rect 11943 4383 11969 4409
rect 14239 4383 14265 4409
rect 2233 4299 2259 4325
rect 2285 4299 2311 4325
rect 2337 4299 2363 4325
rect 12233 4299 12259 4325
rect 12285 4299 12311 4325
rect 12337 4299 12363 4325
rect 11831 4215 11857 4241
rect 2311 4159 2337 4185
rect 4159 4159 4185 4185
rect 4439 4159 4465 4185
rect 4719 4159 4745 4185
rect 4887 4159 4913 4185
rect 5279 4159 5305 4185
rect 5503 4159 5529 4185
rect 5951 4159 5977 4185
rect 6231 4159 6257 4185
rect 6399 4159 6425 4185
rect 12727 4159 12753 4185
rect 2591 4103 2617 4129
rect 3375 4103 3401 4129
rect 5783 4103 5809 4129
rect 7799 4103 7825 4129
rect 12447 4103 12473 4129
rect 13231 4103 13257 4129
rect 14015 4103 14041 4129
rect 14687 4103 14713 4129
rect 2927 4047 2953 4073
rect 3823 4047 3849 4073
rect 5055 4047 5081 4073
rect 7631 4047 7657 4073
rect 8079 4047 8105 4073
rect 13623 4047 13649 4073
rect 14407 4047 14433 4073
rect 15191 3991 15217 4017
rect 1903 3907 1929 3933
rect 1955 3907 1981 3933
rect 2007 3907 2033 3933
rect 11903 3907 11929 3933
rect 11955 3907 11981 3933
rect 12007 3907 12033 3933
rect 2759 3767 2785 3793
rect 3431 3767 3457 3793
rect 4103 3767 4129 3793
rect 5167 3767 5193 3793
rect 5615 3767 5641 3793
rect 5671 3767 5697 3793
rect 5951 3767 5977 3793
rect 8079 3767 8105 3793
rect 12839 3767 12865 3793
rect 13679 3767 13705 3793
rect 15135 3767 15161 3793
rect 3711 3711 3737 3737
rect 3823 3711 3849 3737
rect 7799 3711 7825 3737
rect 13119 3711 13145 3737
rect 14687 3711 14713 3737
rect 4327 3655 4353 3681
rect 4439 3655 4465 3681
rect 5447 3655 5473 3681
rect 7631 3655 7657 3681
rect 13343 3655 13369 3681
rect 7239 3599 7265 3625
rect 7351 3599 7377 3625
rect 2233 3515 2259 3541
rect 2285 3515 2311 3541
rect 2337 3515 2363 3541
rect 12233 3515 12259 3541
rect 12285 3515 12311 3541
rect 12337 3515 12363 3541
rect 7687 3431 7713 3457
rect 13119 3375 13145 3401
rect 14687 3375 14713 3401
rect 3879 3319 3905 3345
rect 4159 3319 4185 3345
rect 4439 3319 4465 3345
rect 7183 3319 7209 3345
rect 8359 3319 8385 3345
rect 13903 3319 13929 3345
rect 7015 3263 7041 3289
rect 7463 3263 7489 3289
rect 8079 3263 8105 3289
rect 8639 3263 8665 3289
rect 13623 3263 13649 3289
rect 15191 3263 15217 3289
rect 14407 3207 14433 3233
rect 1903 3123 1929 3149
rect 1955 3123 1981 3149
rect 2007 3123 2033 3149
rect 11903 3123 11929 3149
rect 11955 3123 11981 3149
rect 12007 3123 12033 3149
rect 7519 2983 7545 3009
rect 15135 2983 15161 3009
rect 14743 2927 14769 2953
rect 7071 2815 7097 2841
rect 7239 2815 7265 2841
rect 2233 2731 2259 2757
rect 2285 2731 2311 2757
rect 2337 2731 2363 2757
rect 12233 2731 12259 2757
rect 12285 2731 12311 2757
rect 12337 2731 12363 2757
rect 7239 2647 7265 2673
rect 8863 2647 8889 2673
rect 8079 2591 8105 2617
rect 8695 2591 8721 2617
rect 9143 2591 9169 2617
rect 13903 2591 13929 2617
rect 15079 2591 15105 2617
rect 6623 2535 6649 2561
rect 6791 2535 6817 2561
rect 7519 2535 7545 2561
rect 7631 2535 7657 2561
rect 7799 2535 7825 2561
rect 8415 2535 8441 2561
rect 14687 2535 14713 2561
rect 7071 2479 7097 2505
rect 14407 2479 14433 2505
rect 1903 2339 1929 2365
rect 1955 2339 1981 2365
rect 2007 2339 2033 2365
rect 11903 2339 11929 2365
rect 11955 2339 11981 2365
rect 12007 2339 12033 2365
rect 7127 2199 7153 2225
rect 7519 2199 7545 2225
rect 8135 2199 8161 2225
rect 8751 2199 8777 2225
rect 15135 2199 15161 2225
rect 8303 2143 8329 2169
rect 14687 2143 14713 2169
rect 7015 2031 7041 2057
rect 7295 2031 7321 2057
rect 7687 2031 7713 2057
rect 7855 2031 7881 2057
rect 14575 2031 14601 2057
rect 2233 1947 2259 1973
rect 2285 1947 2311 1973
rect 2337 1947 2363 1973
rect 12233 1947 12259 1973
rect 12285 1947 12311 1973
rect 12337 1947 12363 1973
rect 13567 1807 13593 1833
rect 13903 1807 13929 1833
rect 14295 1807 14321 1833
rect 6959 1751 6985 1777
rect 13287 1751 13313 1777
rect 13679 1751 13705 1777
rect 14743 1751 14769 1777
rect 6791 1695 6817 1721
rect 7239 1695 7265 1721
rect 8023 1695 8049 1721
rect 15191 1695 15217 1721
rect 1903 1555 1929 1581
rect 1955 1555 1981 1581
rect 2007 1555 2033 1581
rect 11903 1555 11929 1581
rect 11955 1555 11981 1581
rect 12007 1555 12033 1581
rect 6847 1415 6873 1441
rect 7295 1415 7321 1441
rect 8359 1415 8385 1441
rect 8919 1415 8945 1441
rect 12055 1415 12081 1441
rect 12951 1415 12977 1441
rect 14295 1415 14321 1441
rect 15135 1415 15161 1441
rect 7015 1359 7041 1385
rect 7519 1359 7545 1385
rect 7687 1359 7713 1385
rect 8639 1359 8665 1385
rect 14687 1359 14713 1385
rect 7967 1303 7993 1329
rect 13343 1303 13369 1329
rect 13735 1303 13761 1329
rect 8135 1247 8161 1273
rect 10711 1247 10737 1273
rect 11663 1247 11689 1273
rect 11775 1247 11801 1273
rect 12615 1247 12641 1273
rect 12727 1247 12753 1273
rect 14519 1247 14545 1273
rect 2233 1163 2259 1189
rect 2285 1163 2311 1189
rect 2337 1163 2363 1189
rect 12233 1163 12259 1189
rect 12285 1163 12311 1189
rect 12337 1163 12363 1189
rect 8527 1079 8553 1105
rect 7407 1023 7433 1049
rect 8079 1023 8105 1049
rect 9591 1023 9617 1049
rect 10655 1023 10681 1049
rect 11103 1023 11129 1049
rect 12839 1023 12865 1049
rect 13119 1023 13145 1049
rect 13903 1023 13929 1049
rect 15079 1023 15105 1049
rect 6959 967 6985 993
rect 7127 967 7153 993
rect 7799 967 7825 993
rect 9311 967 9337 993
rect 9815 967 9841 993
rect 10207 967 10233 993
rect 10375 967 10401 993
rect 10823 967 10849 993
rect 11327 967 11353 993
rect 12559 967 12585 993
rect 14743 967 14769 993
rect 6735 911 6761 937
rect 7631 911 7657 937
rect 9143 911 9169 937
rect 10039 911 10065 937
rect 11551 911 11577 937
rect 12391 911 12417 937
rect 14407 911 14433 937
rect 13623 855 13649 881
rect 1903 771 1929 797
rect 1955 771 1981 797
rect 2007 771 2033 797
rect 11903 771 11929 797
rect 11955 771 11981 797
rect 12007 771 12033 797
rect 15191 687 15217 713
rect 5559 631 5585 657
rect 6343 631 6369 657
rect 7071 631 7097 657
rect 8359 631 8385 657
rect 8527 631 8553 657
rect 9199 631 9225 657
rect 10823 631 10849 657
rect 11607 631 11633 657
rect 14351 631 14377 657
rect 6511 575 6537 601
rect 7855 575 7881 601
rect 12167 575 12193 601
rect 13903 575 13929 601
rect 14687 575 14713 601
rect 8135 519 8161 545
rect 10207 519 10233 545
rect 12951 519 12977 545
rect 13343 519 13369 545
rect 5783 463 5809 489
rect 5895 463 5921 489
rect 6679 463 6705 489
rect 6959 463 6985 489
rect 7463 463 7489 489
rect 7575 463 7601 489
rect 8807 463 8833 489
rect 8919 463 8945 489
rect 9647 463 9673 489
rect 9815 463 9841 489
rect 10039 463 10065 489
rect 10431 463 10457 489
rect 10543 463 10569 489
rect 11103 463 11129 489
rect 11159 463 11185 489
rect 11383 463 11409 489
rect 12447 463 12473 489
rect 2233 379 2259 405
rect 2285 379 2311 405
rect 2337 379 2363 405
rect 12233 379 12259 405
rect 12285 379 12311 405
rect 12337 379 12363 405
<< metal2 >>
rect 2688 7056 2744 7112
rect 2800 7056 2856 7112
rect 2912 7056 2968 7112
rect 3024 7056 3080 7112
rect 3136 7056 3192 7112
rect 3248 7056 3304 7112
rect 3360 7056 3416 7112
rect 3472 7056 3528 7112
rect 3584 7056 3640 7112
rect 3696 7056 3752 7112
rect 3808 7056 3864 7112
rect 3920 7056 3976 7112
rect 4032 7056 4088 7112
rect 4144 7056 4200 7112
rect 4256 7056 4312 7112
rect 4368 7056 4424 7112
rect 4480 7056 4536 7112
rect 4592 7056 4648 7112
rect 4704 7056 4760 7112
rect 4816 7056 4872 7112
rect 4928 7056 4984 7112
rect 5040 7056 5096 7112
rect 5152 7056 5208 7112
rect 5264 7056 5320 7112
rect 5376 7056 5432 7112
rect 5488 7056 5544 7112
rect 5600 7056 5656 7112
rect 5712 7056 5768 7112
rect 5824 7056 5880 7112
rect 5936 7056 5992 7112
rect 6048 7056 6104 7112
rect 6160 7056 6216 7112
rect 6272 7056 6328 7112
rect 6384 7056 6440 7112
rect 6496 7056 6552 7112
rect 6608 7056 6664 7112
rect 6720 7056 6776 7112
rect 6832 7056 6888 7112
rect 6944 7056 7000 7112
rect 7056 7056 7112 7112
rect 7168 7056 7224 7112
rect 7280 7056 7336 7112
rect 7392 7056 7448 7112
rect 7504 7056 7560 7112
rect 7616 7056 7672 7112
rect 7728 7056 7784 7112
rect 7840 7056 7896 7112
rect 7952 7056 8008 7112
rect 8064 7056 8120 7112
rect 8176 7056 8232 7112
rect 8288 7056 8344 7112
rect 8400 7056 8456 7112
rect 8512 7056 8568 7112
rect 8624 7056 8680 7112
rect 8736 7056 8792 7112
rect 8848 7056 8904 7112
rect 8960 7056 9016 7112
rect 9072 7056 9128 7112
rect 9184 7056 9240 7112
rect 9296 7056 9352 7112
rect 9408 7056 9464 7112
rect 9520 7056 9576 7112
rect 9632 7056 9688 7112
rect 9744 7056 9800 7112
rect 9856 7056 9912 7112
rect 9968 7056 10024 7112
rect 10080 7056 10136 7112
rect 10192 7056 10248 7112
rect 10304 7056 10360 7112
rect 10416 7056 10472 7112
rect 10528 7056 10584 7112
rect 10640 7056 10696 7112
rect 10752 7056 10808 7112
rect 10864 7056 10920 7112
rect 10976 7056 11032 7112
rect 11088 7056 11144 7112
rect 11200 7056 11256 7112
rect 11312 7056 11368 7112
rect 11424 7056 11480 7112
rect 11536 7056 11592 7112
rect 11648 7056 11704 7112
rect 11760 7056 11816 7112
rect 11872 7056 11928 7112
rect 11984 7056 12040 7112
rect 12096 7056 12152 7112
rect 12208 7056 12264 7112
rect 12320 7056 12376 7112
rect 12432 7056 12488 7112
rect 12544 7056 12600 7112
rect 12656 7056 12712 7112
rect 12768 7056 12824 7112
rect 12880 7056 12936 7112
rect 12992 7056 13048 7112
rect 126 6986 154 6991
rect 70 6090 98 6095
rect 70 2450 98 6062
rect 126 3066 154 6958
rect 2086 6930 2114 6935
rect 1862 6874 1890 6879
rect 1078 6594 1106 6599
rect 1078 6547 1106 6566
rect 1862 6593 1890 6846
rect 1862 6567 1863 6593
rect 1889 6567 1890 6593
rect 1862 6561 1890 6567
rect 1358 6481 1386 6487
rect 1358 6455 1359 6481
rect 1385 6455 1386 6481
rect 1246 6314 1274 6319
rect 1078 5866 1106 5871
rect 686 5642 714 5647
rect 406 5194 434 5199
rect 406 4914 434 5166
rect 406 4881 434 4886
rect 686 3458 714 5614
rect 910 4746 938 4751
rect 910 4410 938 4718
rect 910 4377 938 4382
rect 686 3425 714 3430
rect 126 3033 154 3038
rect 126 2450 154 2455
rect 70 2422 126 2450
rect 126 2417 154 2422
rect 1078 1498 1106 5838
rect 1246 1890 1274 6286
rect 1358 5194 1386 6455
rect 1902 6286 2034 6291
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 1902 6253 2034 6258
rect 1918 6202 1946 6207
rect 1918 6155 1946 6174
rect 1806 5810 1834 5815
rect 1806 5753 1834 5782
rect 1806 5727 1807 5753
rect 1833 5727 1834 5753
rect 1806 5721 1834 5727
rect 1582 5697 1610 5703
rect 1582 5671 1583 5697
rect 1609 5671 1610 5697
rect 1414 5642 1442 5647
rect 1582 5642 1610 5671
rect 1414 5641 1610 5642
rect 1414 5615 1415 5641
rect 1441 5615 1610 5641
rect 1414 5614 1610 5615
rect 1414 5609 1442 5614
rect 1358 5161 1386 5166
rect 1582 4130 1610 5614
rect 1806 5642 1834 5647
rect 1806 5361 1834 5614
rect 1902 5502 2034 5507
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 1902 5469 2034 5474
rect 1806 5335 1807 5361
rect 1833 5335 1834 5361
rect 1806 5329 1834 5335
rect 2030 4913 2058 4919
rect 2030 4887 2031 4913
rect 2057 4887 2058 4913
rect 2030 4802 2058 4887
rect 2086 4914 2114 6902
rect 2232 6678 2364 6683
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2232 6645 2364 6650
rect 2142 6482 2170 6487
rect 2142 6481 2506 6482
rect 2142 6455 2143 6481
rect 2169 6455 2506 6481
rect 2142 6454 2506 6455
rect 2142 6449 2170 6454
rect 2198 6034 2226 6039
rect 2198 5987 2226 6006
rect 2232 5894 2364 5899
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2232 5861 2364 5866
rect 2310 5809 2338 5815
rect 2310 5783 2311 5809
rect 2337 5783 2338 5809
rect 2310 5754 2338 5783
rect 2310 5721 2338 5726
rect 2422 5698 2450 5703
rect 2142 5305 2170 5311
rect 2142 5279 2143 5305
rect 2169 5279 2170 5305
rect 2142 5026 2170 5279
rect 2232 5110 2364 5115
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2232 5077 2364 5082
rect 2142 4993 2170 4998
rect 2086 4886 2170 4914
rect 2030 4774 2114 4802
rect 1902 4718 2034 4723
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 1902 4685 2034 4690
rect 1862 4466 1890 4471
rect 1862 4419 1890 4438
rect 2086 4214 2114 4774
rect 2142 4578 2170 4886
rect 2422 4857 2450 5670
rect 2422 4831 2423 4857
rect 2449 4831 2450 4857
rect 2422 4825 2450 4831
rect 2422 4578 2450 4583
rect 2142 4577 2450 4578
rect 2142 4551 2423 4577
rect 2449 4551 2450 4577
rect 2142 4550 2450 4551
rect 2142 4521 2170 4550
rect 2422 4545 2450 4550
rect 2142 4495 2143 4521
rect 2169 4495 2170 4521
rect 2142 4489 2170 4495
rect 2232 4326 2364 4331
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2232 4293 2364 4298
rect 2086 4186 2338 4214
rect 2310 4185 2338 4186
rect 2310 4159 2311 4185
rect 2337 4159 2338 4185
rect 2310 4153 2338 4159
rect 1582 4097 1610 4102
rect 1902 3934 2034 3939
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 1902 3901 2034 3906
rect 2478 3906 2506 6454
rect 2590 6146 2618 6151
rect 2590 6099 2618 6118
rect 2534 5697 2562 5703
rect 2534 5671 2535 5697
rect 2561 5671 2562 5697
rect 2534 4858 2562 5671
rect 2702 5642 2730 7056
rect 2758 6146 2786 6151
rect 2758 6089 2786 6118
rect 2758 6063 2759 6089
rect 2785 6063 2786 6089
rect 2758 6057 2786 6063
rect 2702 5609 2730 5614
rect 2590 5362 2618 5367
rect 2590 5315 2618 5334
rect 2758 5362 2786 5367
rect 2758 5305 2786 5334
rect 2758 5279 2759 5305
rect 2785 5279 2786 5305
rect 2758 5273 2786 5279
rect 2534 4825 2562 4830
rect 2646 4914 2674 4919
rect 2590 4466 2618 4471
rect 2590 4419 2618 4438
rect 2590 4129 2618 4135
rect 2590 4103 2591 4129
rect 2617 4103 2618 4129
rect 2590 3962 2618 4103
rect 2590 3929 2618 3934
rect 2478 3873 2506 3878
rect 2534 3850 2562 3855
rect 2232 3542 2364 3547
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2232 3509 2364 3514
rect 1902 3150 2034 3155
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 1902 3117 2034 3122
rect 2232 2758 2364 2763
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2232 2725 2364 2730
rect 1414 2506 1442 2511
rect 1414 2170 1442 2478
rect 2534 2506 2562 3822
rect 2646 2842 2674 4886
rect 2814 4214 2842 7056
rect 2926 6202 2954 7056
rect 2982 6650 3010 6655
rect 2982 6593 3010 6622
rect 2982 6567 2983 6593
rect 3009 6567 3010 6593
rect 2982 6561 3010 6567
rect 2870 6174 2954 6202
rect 2870 5698 2898 6174
rect 3038 6146 3066 7056
rect 3150 6594 3178 7056
rect 3262 6706 3290 7056
rect 3150 6561 3178 6566
rect 3206 6678 3290 6706
rect 2870 5665 2898 5670
rect 2926 6118 3066 6146
rect 2926 4577 2954 6118
rect 2982 6034 3010 6039
rect 3150 6034 3178 6039
rect 2982 6033 3178 6034
rect 2982 6007 2983 6033
rect 3009 6007 3151 6033
rect 3177 6007 3178 6033
rect 2982 6006 3178 6007
rect 2982 6001 3010 6006
rect 3150 6001 3178 6006
rect 2982 5922 3010 5927
rect 2982 5361 3010 5894
rect 3094 5866 3122 5871
rect 3094 5809 3122 5838
rect 3094 5783 3095 5809
rect 3121 5783 3122 5809
rect 3094 5777 3122 5783
rect 3206 5754 3234 6678
rect 3262 6594 3290 6599
rect 3262 6537 3290 6566
rect 3262 6511 3263 6537
rect 3289 6511 3290 6537
rect 3262 6505 3290 6511
rect 3374 6202 3402 7056
rect 3374 6169 3402 6174
rect 3206 5721 3234 5726
rect 3262 5697 3290 5703
rect 3262 5671 3263 5697
rect 3289 5671 3290 5697
rect 2982 5335 2983 5361
rect 3009 5335 3010 5361
rect 2982 5329 3010 5335
rect 3094 5530 3122 5535
rect 3094 5025 3122 5502
rect 3094 4999 3095 5025
rect 3121 4999 3122 5025
rect 3094 4993 3122 4999
rect 2926 4551 2927 4577
rect 2953 4551 2954 4577
rect 2926 4545 2954 4551
rect 3262 4298 3290 5671
rect 3486 5530 3514 7056
rect 3486 5497 3514 5502
rect 3486 5418 3514 5423
rect 3486 5371 3514 5390
rect 3318 4914 3346 4919
rect 3318 4867 3346 4886
rect 3598 4802 3626 7056
rect 3654 6258 3682 6263
rect 3654 6201 3682 6230
rect 3654 6175 3655 6201
rect 3681 6175 3682 6201
rect 3654 6169 3682 6175
rect 3598 4769 3626 4774
rect 3710 4633 3738 7056
rect 3822 6874 3850 7056
rect 3822 6841 3850 6846
rect 3766 6818 3794 6823
rect 3766 6593 3794 6790
rect 3934 6594 3962 7056
rect 3766 6567 3767 6593
rect 3793 6567 3794 6593
rect 3766 6561 3794 6567
rect 3878 6566 3962 6594
rect 3766 6090 3794 6095
rect 3766 5305 3794 6062
rect 3878 5866 3906 6566
rect 3878 5833 3906 5838
rect 3934 6481 3962 6487
rect 3934 6455 3935 6481
rect 3961 6455 3962 6481
rect 3878 5642 3906 5647
rect 3878 5595 3906 5614
rect 3934 5362 3962 6455
rect 4046 5418 4074 7056
rect 4158 6818 4186 7056
rect 4046 5385 4074 5390
rect 4102 6790 4186 6818
rect 3766 5279 3767 5305
rect 3793 5279 3794 5305
rect 3766 5273 3794 5279
rect 3822 5334 3962 5362
rect 3710 4607 3711 4633
rect 3737 4607 3738 4633
rect 3710 4601 3738 4607
rect 3822 4522 3850 5334
rect 4102 5306 4130 6790
rect 4158 6706 4186 6711
rect 4158 6145 4186 6678
rect 4158 6119 4159 6145
rect 4185 6119 4186 6145
rect 4158 6113 4186 6119
rect 4214 6202 4242 6207
rect 4158 5698 4186 5703
rect 4158 5651 4186 5670
rect 3878 5278 4130 5306
rect 4158 5474 4186 5479
rect 3878 5025 3906 5278
rect 3878 4999 3879 5025
rect 3905 4999 3906 5025
rect 3878 4993 3906 4999
rect 4158 4969 4186 5446
rect 4214 5361 4242 6174
rect 4270 5754 4298 7056
rect 4382 6650 4410 7056
rect 4382 6617 4410 6622
rect 4494 6370 4522 7056
rect 4438 6342 4522 6370
rect 4270 5726 4354 5754
rect 4214 5335 4215 5361
rect 4241 5335 4242 5361
rect 4214 5329 4242 5335
rect 4158 4943 4159 4969
rect 4185 4943 4186 4969
rect 4158 4937 4186 4943
rect 3262 4265 3290 4270
rect 3598 4494 3850 4522
rect 3878 4802 3906 4807
rect 2814 4186 2954 4214
rect 2926 4073 2954 4186
rect 2926 4047 2927 4073
rect 2953 4047 2954 4073
rect 2926 4041 2954 4047
rect 3374 4129 3402 4135
rect 3374 4103 3375 4129
rect 3401 4103 3402 4129
rect 2758 3962 2786 3967
rect 2758 3793 2786 3934
rect 2758 3767 2759 3793
rect 2785 3767 2786 3793
rect 2758 3761 2786 3767
rect 3374 3794 3402 4103
rect 3486 4130 3514 4135
rect 3430 3794 3458 3799
rect 3374 3793 3458 3794
rect 3374 3767 3431 3793
rect 3457 3767 3458 3793
rect 3374 3766 3458 3767
rect 3430 3761 3458 3766
rect 2646 2809 2674 2814
rect 3374 3458 3402 3463
rect 2534 2473 2562 2478
rect 1902 2366 2034 2371
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 1902 2333 2034 2338
rect 1414 2137 1442 2142
rect 3374 2002 3402 3430
rect 2232 1974 2364 1979
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 3374 1969 3402 1974
rect 2232 1941 2364 1946
rect 1246 1857 1274 1862
rect 1902 1582 2034 1587
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 1902 1549 2034 1554
rect 1078 1465 1106 1470
rect 2232 1190 2364 1195
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2232 1157 2364 1162
rect 3150 994 3178 999
rect 1806 882 1834 887
rect 1134 98 1162 103
rect 1134 56 1162 70
rect 1806 56 1834 854
rect 1902 798 2034 803
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 1902 765 2034 770
rect 2232 406 2364 411
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2232 373 2364 378
rect 2478 98 2506 103
rect 2478 56 2506 70
rect 3150 56 3178 966
rect 3486 826 3514 4102
rect 3486 793 3514 798
rect 3598 434 3626 4494
rect 3878 4214 3906 4774
rect 4102 4746 4130 4751
rect 3822 4186 3906 4214
rect 3990 4465 4018 4471
rect 3990 4439 3991 4465
rect 4017 4439 4018 4465
rect 3822 4073 3850 4186
rect 3822 4047 3823 4073
rect 3849 4047 3850 4073
rect 3822 4041 3850 4047
rect 3990 4074 4018 4439
rect 3990 4041 4018 4046
rect 4102 3793 4130 4718
rect 4326 4577 4354 5726
rect 4438 5642 4466 6342
rect 4606 6202 4634 7056
rect 4718 6258 4746 7056
rect 4718 6225 4746 6230
rect 4774 6986 4802 6991
rect 4606 6169 4634 6174
rect 4494 6034 4522 6039
rect 4494 5753 4522 6006
rect 4550 6034 4578 6039
rect 4550 6033 4690 6034
rect 4550 6007 4551 6033
rect 4577 6007 4690 6033
rect 4550 6006 4690 6007
rect 4550 6001 4578 6006
rect 4494 5727 4495 5753
rect 4521 5727 4522 5753
rect 4494 5721 4522 5727
rect 4550 5922 4578 5927
rect 4438 5609 4466 5614
rect 4550 5305 4578 5894
rect 4662 5866 4690 6006
rect 4662 5833 4690 5838
rect 4774 5809 4802 6958
rect 4774 5783 4775 5809
rect 4801 5783 4802 5809
rect 4774 5777 4802 5783
rect 4718 5698 4746 5703
rect 4550 5279 4551 5305
rect 4577 5279 4578 5305
rect 4550 5273 4578 5279
rect 4662 5697 4746 5698
rect 4662 5671 4719 5697
rect 4745 5671 4746 5697
rect 4662 5670 4746 5671
rect 4326 4551 4327 4577
rect 4353 4551 4354 4577
rect 4326 4545 4354 4551
rect 4438 5026 4466 5031
rect 4158 4466 4186 4471
rect 4158 4185 4186 4438
rect 4158 4159 4159 4185
rect 4185 4159 4186 4185
rect 4158 4153 4186 4159
rect 4438 4185 4466 4998
rect 4606 5026 4634 5031
rect 4662 5026 4690 5670
rect 4718 5665 4746 5670
rect 4830 5306 4858 7056
rect 4886 6874 4914 6879
rect 4886 6593 4914 6846
rect 4886 6567 4887 6593
rect 4913 6567 4914 6593
rect 4886 6561 4914 6567
rect 4830 5273 4858 5278
rect 4606 5025 4690 5026
rect 4606 4999 4607 5025
rect 4633 4999 4690 5025
rect 4606 4998 4690 4999
rect 4606 4993 4634 4998
rect 4942 4969 4970 7056
rect 4942 4943 4943 4969
rect 4969 4943 4970 4969
rect 4942 4937 4970 4943
rect 4998 6986 5026 6991
rect 4998 4858 5026 6958
rect 5054 6818 5082 7056
rect 5054 6785 5082 6790
rect 5166 6706 5194 7056
rect 5166 6673 5194 6678
rect 5166 6481 5194 6487
rect 5166 6455 5167 6481
rect 5193 6455 5194 6481
rect 5166 6314 5194 6455
rect 5166 6281 5194 6286
rect 5054 6202 5082 6207
rect 5054 6155 5082 6174
rect 5166 6146 5194 6151
rect 5166 5753 5194 6118
rect 5166 5727 5167 5753
rect 5193 5727 5194 5753
rect 5166 5721 5194 5727
rect 5054 5418 5082 5423
rect 5278 5418 5306 7056
rect 5334 6034 5362 6039
rect 5334 5987 5362 6006
rect 5390 5866 5418 7056
rect 5502 6146 5530 7056
rect 5614 6202 5642 7056
rect 5670 6650 5698 6655
rect 5670 6593 5698 6622
rect 5670 6567 5671 6593
rect 5697 6567 5698 6593
rect 5670 6561 5698 6567
rect 5614 6169 5642 6174
rect 5502 6113 5530 6118
rect 5502 6033 5530 6039
rect 5502 6007 5503 6033
rect 5529 6007 5530 6033
rect 5502 5978 5530 6007
rect 5502 5945 5530 5950
rect 5726 5866 5754 7056
rect 5838 6874 5866 7056
rect 5838 6841 5866 6846
rect 5950 6706 5978 7056
rect 5950 6673 5978 6678
rect 5950 6481 5978 6487
rect 5950 6455 5951 6481
rect 5977 6455 5978 6481
rect 5950 6258 5978 6455
rect 5950 6225 5978 6230
rect 6006 6202 6034 6207
rect 6006 6155 6034 6174
rect 5838 5866 5866 5871
rect 5390 5838 5642 5866
rect 5726 5838 5810 5866
rect 5054 5417 5306 5418
rect 5054 5391 5055 5417
rect 5081 5391 5306 5417
rect 5054 5390 5306 5391
rect 5558 5697 5586 5703
rect 5558 5671 5559 5697
rect 5585 5671 5586 5697
rect 5054 5385 5082 5390
rect 5334 5362 5362 5367
rect 4886 4830 5026 4858
rect 5222 5306 5250 5311
rect 4774 4634 4802 4639
rect 4774 4521 4802 4606
rect 4774 4495 4775 4521
rect 4801 4495 4802 4521
rect 4774 4489 4802 4495
rect 4438 4159 4439 4185
rect 4465 4159 4466 4185
rect 4438 4153 4466 4159
rect 4718 4186 4746 4191
rect 4886 4186 4914 4830
rect 5222 4633 5250 5278
rect 5334 5305 5362 5334
rect 5334 5279 5335 5305
rect 5361 5279 5362 5305
rect 5334 5273 5362 5279
rect 5222 4607 5223 4633
rect 5249 4607 5250 4633
rect 5222 4601 5250 4607
rect 5334 4913 5362 4919
rect 5334 4887 5335 4913
rect 5361 4887 5362 4913
rect 5334 4578 5362 4887
rect 5334 4545 5362 4550
rect 4718 4185 4914 4186
rect 4718 4159 4719 4185
rect 4745 4159 4887 4185
rect 4913 4159 4914 4185
rect 4718 4158 4914 4159
rect 4718 4153 4746 4158
rect 4886 4153 4914 4158
rect 4942 4465 4970 4471
rect 4942 4439 4943 4465
rect 4969 4439 4970 4465
rect 4102 3767 4103 3793
rect 4129 3767 4130 3793
rect 4102 3761 4130 3767
rect 3710 3738 3738 3743
rect 3822 3738 3850 3743
rect 3710 3737 3822 3738
rect 3710 3711 3711 3737
rect 3737 3711 3822 3737
rect 3710 3710 3822 3711
rect 3710 3705 3738 3710
rect 3822 3691 3850 3710
rect 4326 3682 4354 3687
rect 4326 3635 4354 3654
rect 4438 3682 4466 3687
rect 4438 3635 4466 3654
rect 3878 3458 3906 3463
rect 3878 3345 3906 3430
rect 4942 3458 4970 4439
rect 5278 4354 5306 4359
rect 5278 4185 5306 4326
rect 5278 4159 5279 4185
rect 5305 4159 5306 4185
rect 5278 4153 5306 4159
rect 5502 4298 5530 4303
rect 5502 4185 5530 4270
rect 5502 4159 5503 4185
rect 5529 4159 5530 4185
rect 5502 4153 5530 4159
rect 5054 4074 5082 4079
rect 5054 4027 5082 4046
rect 5558 4018 5586 5671
rect 5614 4857 5642 5838
rect 5726 5697 5754 5703
rect 5726 5671 5727 5697
rect 5753 5671 5754 5697
rect 5614 4831 5615 4857
rect 5641 4831 5642 4857
rect 5614 4825 5642 4831
rect 5670 5642 5698 5647
rect 5558 3985 5586 3990
rect 5614 4354 5642 4359
rect 5166 3906 5194 3911
rect 5166 3793 5194 3878
rect 5166 3767 5167 3793
rect 5193 3767 5194 3793
rect 5166 3761 5194 3767
rect 5614 3793 5642 4326
rect 5614 3767 5615 3793
rect 5641 3767 5642 3793
rect 5614 3761 5642 3767
rect 5670 3793 5698 5614
rect 5726 4746 5754 5671
rect 5782 5361 5810 5838
rect 5782 5335 5783 5361
rect 5809 5335 5810 5361
rect 5782 5329 5810 5335
rect 5726 4713 5754 4718
rect 5726 4466 5754 4471
rect 5726 4419 5754 4438
rect 5838 4298 5866 5838
rect 6062 5641 6090 7056
rect 6174 6202 6202 7056
rect 6286 6650 6314 7056
rect 6286 6617 6314 6622
rect 6342 6706 6370 6711
rect 6174 6169 6202 6174
rect 6286 6425 6314 6431
rect 6286 6399 6287 6425
rect 6313 6399 6314 6425
rect 6286 5698 6314 6399
rect 6286 5665 6314 5670
rect 6062 5615 6063 5641
rect 6089 5615 6090 5641
rect 6062 5609 6090 5615
rect 6342 5586 6370 6678
rect 6398 5642 6426 7056
rect 6510 6146 6538 7056
rect 6510 6113 6538 6118
rect 6566 6818 6594 6823
rect 6566 6593 6594 6790
rect 6566 6567 6567 6593
rect 6593 6567 6594 6593
rect 6510 6034 6538 6039
rect 6566 6034 6594 6567
rect 6622 6594 6650 7056
rect 6734 6930 6762 7056
rect 6734 6897 6762 6902
rect 6622 6561 6650 6566
rect 6734 6481 6762 6487
rect 6734 6455 6735 6481
rect 6761 6455 6762 6481
rect 6510 6033 6594 6034
rect 6510 6007 6511 6033
rect 6537 6007 6594 6033
rect 6510 6006 6594 6007
rect 6678 6426 6706 6431
rect 6510 6001 6538 6006
rect 6622 5642 6650 5647
rect 6398 5641 6650 5642
rect 6398 5615 6623 5641
rect 6649 5615 6650 5641
rect 6398 5614 6650 5615
rect 6622 5609 6650 5614
rect 6342 5558 6538 5586
rect 6510 5417 6538 5558
rect 6510 5391 6511 5417
rect 6537 5391 6538 5417
rect 6510 5385 6538 5391
rect 6454 5306 6482 5311
rect 6118 5250 6146 5255
rect 6118 5203 6146 5222
rect 6174 5138 6202 5143
rect 5838 4265 5866 4270
rect 5950 4914 5978 4919
rect 5950 4185 5978 4886
rect 6118 4914 6146 4919
rect 6118 4867 6146 4886
rect 6118 4578 6146 4583
rect 6174 4578 6202 5110
rect 6454 4969 6482 5278
rect 6454 4943 6455 4969
rect 6481 4943 6482 4969
rect 6454 4937 6482 4943
rect 6678 4913 6706 6398
rect 6734 5306 6762 6455
rect 6790 6146 6818 6151
rect 6790 6099 6818 6118
rect 6734 5273 6762 5278
rect 6790 5754 6818 5759
rect 6678 4887 6679 4913
rect 6705 4887 6706 4913
rect 6678 4690 6706 4887
rect 6678 4657 6706 4662
rect 6006 4577 6202 4578
rect 6006 4551 6119 4577
rect 6145 4551 6202 4577
rect 6006 4550 6202 4551
rect 6006 4521 6034 4550
rect 6118 4545 6146 4550
rect 6006 4495 6007 4521
rect 6033 4495 6034 4521
rect 6006 4489 6034 4495
rect 6790 4354 6818 5726
rect 6790 4321 6818 4326
rect 5950 4159 5951 4185
rect 5977 4159 5978 4185
rect 5950 4153 5978 4159
rect 6230 4186 6258 4191
rect 6230 4139 6258 4158
rect 6398 4186 6426 4191
rect 6398 4139 6426 4158
rect 5782 4130 5810 4135
rect 5782 4083 5810 4102
rect 5670 3767 5671 3793
rect 5697 3767 5698 3793
rect 5446 3682 5474 3687
rect 5670 3682 5698 3767
rect 5950 4074 5978 4079
rect 5950 3793 5978 4046
rect 6846 3962 6874 7056
rect 6958 6090 6986 7056
rect 7070 6986 7098 7056
rect 7070 6953 7098 6958
rect 7014 6594 7042 6599
rect 7014 6547 7042 6566
rect 7126 6370 7154 6375
rect 6902 6062 6986 6090
rect 7014 6146 7042 6151
rect 6902 5586 6930 6062
rect 6902 5558 6986 5586
rect 6902 4858 6930 4863
rect 6902 4811 6930 4830
rect 6902 4690 6930 4695
rect 6902 4577 6930 4662
rect 6902 4551 6903 4577
rect 6929 4551 6930 4577
rect 6902 4545 6930 4551
rect 6846 3929 6874 3934
rect 5950 3767 5951 3793
rect 5977 3767 5978 3793
rect 5950 3761 5978 3767
rect 6902 3906 6930 3911
rect 5446 3681 5698 3682
rect 5446 3655 5447 3681
rect 5473 3655 5698 3681
rect 5446 3654 5698 3655
rect 5446 3649 5474 3654
rect 4942 3425 4970 3430
rect 3878 3319 3879 3345
rect 3905 3319 3906 3345
rect 3878 3313 3906 3319
rect 4158 3345 4186 3351
rect 4158 3319 4159 3345
rect 4185 3319 4186 3345
rect 4158 3234 4186 3319
rect 4158 3201 4186 3206
rect 4438 3346 4466 3351
rect 4438 3234 4466 3318
rect 4438 3201 4466 3206
rect 6622 2562 6650 2567
rect 6790 2562 6818 2567
rect 6622 2561 6818 2562
rect 6622 2535 6623 2561
rect 6649 2535 6791 2561
rect 6817 2535 6818 2561
rect 6622 2534 6818 2535
rect 6622 2058 6650 2534
rect 6790 2529 6818 2534
rect 6622 2025 6650 2030
rect 6902 1834 6930 3878
rect 6958 3738 6986 5558
rect 7014 5305 7042 6118
rect 7126 5753 7154 6342
rect 7126 5727 7127 5753
rect 7153 5727 7154 5753
rect 7126 5721 7154 5727
rect 7182 5586 7210 7056
rect 7238 6202 7266 6207
rect 7238 6089 7266 6174
rect 7238 6063 7239 6089
rect 7265 6063 7266 6089
rect 7238 6057 7266 6063
rect 7294 5642 7322 7056
rect 7294 5609 7322 5614
rect 7350 6706 7378 6711
rect 7014 5279 7015 5305
rect 7041 5279 7042 5305
rect 7014 5273 7042 5279
rect 7070 5558 7210 5586
rect 7070 4130 7098 5558
rect 7070 4097 7098 4102
rect 7126 5474 7154 5479
rect 6958 3705 6986 3710
rect 7126 3570 7154 5446
rect 7182 5249 7210 5255
rect 7182 5223 7183 5249
rect 7209 5223 7210 5249
rect 7182 5194 7210 5223
rect 7182 5161 7210 5166
rect 7182 5026 7210 5031
rect 7350 5026 7378 6678
rect 7406 6146 7434 7056
rect 7406 6118 7490 6146
rect 7406 6033 7434 6039
rect 7406 6007 7407 6033
rect 7433 6007 7434 6033
rect 7406 5922 7434 6007
rect 7406 5889 7434 5894
rect 7462 5754 7490 6118
rect 7462 5721 7490 5726
rect 7462 5641 7490 5647
rect 7462 5615 7463 5641
rect 7489 5615 7490 5641
rect 7462 5474 7490 5615
rect 7462 5441 7490 5446
rect 7406 5418 7434 5423
rect 7406 5305 7434 5390
rect 7406 5279 7407 5305
rect 7433 5279 7434 5305
rect 7406 5273 7434 5279
rect 7518 5138 7546 7056
rect 7574 6538 7602 6543
rect 7574 6491 7602 6510
rect 7630 5810 7658 7056
rect 7742 7042 7770 7056
rect 7742 7009 7770 7014
rect 7854 6706 7882 7056
rect 7854 6673 7882 6678
rect 7854 6594 7882 6599
rect 7854 6547 7882 6566
rect 7854 6033 7882 6039
rect 7854 6007 7855 6033
rect 7881 6007 7882 6033
rect 7686 5977 7714 5983
rect 7686 5951 7687 5977
rect 7713 5951 7714 5977
rect 7686 5922 7714 5951
rect 7686 5889 7714 5894
rect 7518 5105 7546 5110
rect 7574 5782 7658 5810
rect 7182 5025 7378 5026
rect 7182 4999 7183 5025
rect 7209 4999 7351 5025
rect 7377 4999 7378 5025
rect 7182 4998 7378 4999
rect 7182 4993 7210 4998
rect 7350 4993 7378 4998
rect 7462 4858 7490 4863
rect 7462 4522 7490 4830
rect 7574 4746 7602 5782
rect 7630 5697 7658 5703
rect 7630 5671 7631 5697
rect 7657 5671 7658 5697
rect 7630 5474 7658 5671
rect 7630 5441 7658 5446
rect 7686 5418 7714 5423
rect 7686 5362 7714 5390
rect 7630 5334 7714 5362
rect 7630 5025 7658 5334
rect 7630 4999 7631 5025
rect 7657 4999 7658 5025
rect 7630 4993 7658 4999
rect 7686 5193 7714 5199
rect 7686 5167 7687 5193
rect 7713 5167 7714 5193
rect 7686 4858 7714 5167
rect 7686 4825 7714 4830
rect 7574 4718 7658 4746
rect 7462 4489 7490 4494
rect 7406 4410 7434 4415
rect 7406 4363 7434 4382
rect 7574 4410 7602 4415
rect 7574 4363 7602 4382
rect 7630 4186 7658 4718
rect 7854 4634 7882 6007
rect 7910 5642 7938 5647
rect 7910 5595 7938 5614
rect 7966 5418 7994 7056
rect 8078 6874 8106 7056
rect 7966 5385 7994 5390
rect 8022 6846 8106 6874
rect 7966 5249 7994 5255
rect 7966 5223 7967 5249
rect 7993 5223 7994 5249
rect 7966 4970 7994 5223
rect 7966 4937 7994 4942
rect 7854 4601 7882 4606
rect 7966 4858 7994 4863
rect 7854 4465 7882 4471
rect 7854 4439 7855 4465
rect 7881 4439 7882 4465
rect 7854 4242 7882 4439
rect 7966 4298 7994 4830
rect 7966 4265 7994 4270
rect 7854 4209 7882 4214
rect 7630 4153 7658 4158
rect 7798 4129 7826 4135
rect 7798 4103 7799 4129
rect 7825 4103 7826 4129
rect 7630 4074 7658 4079
rect 7798 4074 7826 4103
rect 7574 4073 7826 4074
rect 7574 4047 7631 4073
rect 7657 4047 7826 4073
rect 7574 4046 7826 4047
rect 7126 3537 7154 3542
rect 7238 3626 7266 3631
rect 7350 3626 7378 3631
rect 7238 3625 7378 3626
rect 7238 3599 7239 3625
rect 7265 3599 7351 3625
rect 7377 3599 7378 3625
rect 7238 3598 7378 3599
rect 7238 3402 7266 3598
rect 7350 3593 7378 3598
rect 7574 3514 7602 4046
rect 7630 4041 7658 4046
rect 7686 3794 7714 3799
rect 7630 3681 7658 3687
rect 7630 3655 7631 3681
rect 7657 3655 7658 3681
rect 7630 3626 7658 3655
rect 7630 3593 7658 3598
rect 7574 3481 7602 3486
rect 7686 3457 7714 3766
rect 7798 3794 7826 3799
rect 7798 3737 7826 3766
rect 7798 3711 7799 3737
rect 7825 3711 7826 3737
rect 7798 3705 7826 3711
rect 7686 3431 7687 3457
rect 7713 3431 7714 3457
rect 7686 3425 7714 3431
rect 7238 3369 7266 3374
rect 7182 3345 7210 3351
rect 7182 3319 7183 3345
rect 7209 3319 7210 3345
rect 7014 3290 7042 3295
rect 7014 3243 7042 3262
rect 7182 3290 7210 3319
rect 7966 3346 7994 3351
rect 8022 3346 8050 6846
rect 8190 6818 8218 7056
rect 8078 6790 8218 6818
rect 8246 6930 8274 6935
rect 8078 6482 8106 6790
rect 8134 6594 8162 6599
rect 8246 6594 8274 6902
rect 8134 6547 8162 6566
rect 8190 6593 8274 6594
rect 8190 6567 8247 6593
rect 8273 6567 8274 6593
rect 8190 6566 8274 6567
rect 8078 6449 8106 6454
rect 8134 6090 8162 6095
rect 8190 6090 8218 6566
rect 8246 6561 8274 6566
rect 8302 6258 8330 7056
rect 8414 6818 8442 7056
rect 8414 6785 8442 6790
rect 8526 6594 8554 7056
rect 8638 6930 8666 7056
rect 8638 6897 8666 6902
rect 8750 6818 8778 7056
rect 8526 6561 8554 6566
rect 8582 6790 8778 6818
rect 8134 6089 8218 6090
rect 8134 6063 8135 6089
rect 8161 6063 8218 6089
rect 8134 6062 8218 6063
rect 8246 6230 8330 6258
rect 8134 6057 8162 6062
rect 8246 5978 8274 6230
rect 8582 6090 8610 6790
rect 8694 6706 8722 6711
rect 8694 6594 8722 6678
rect 8750 6594 8778 6599
rect 8694 6593 8778 6594
rect 8694 6567 8751 6593
rect 8777 6567 8778 6593
rect 8694 6566 8778 6567
rect 8750 6561 8778 6566
rect 8862 6538 8890 7056
rect 8862 6505 8890 6510
rect 8862 6425 8890 6431
rect 8862 6399 8863 6425
rect 8889 6399 8890 6425
rect 8806 6314 8834 6319
rect 8750 6090 8778 6095
rect 8582 6089 8722 6090
rect 8582 6063 8583 6089
rect 8609 6063 8722 6089
rect 8582 6062 8722 6063
rect 8582 6057 8610 6062
rect 8078 5950 8274 5978
rect 8302 6033 8330 6039
rect 8302 6007 8303 6033
rect 8329 6007 8330 6033
rect 8078 5922 8106 5950
rect 8078 5809 8106 5894
rect 8078 5783 8079 5809
rect 8105 5783 8106 5809
rect 8078 5777 8106 5783
rect 8302 5530 8330 6007
rect 8694 5810 8722 6062
rect 8750 6043 8778 6062
rect 8750 5810 8778 5815
rect 8694 5809 8778 5810
rect 8694 5783 8751 5809
rect 8777 5783 8778 5809
rect 8694 5782 8778 5783
rect 8750 5777 8778 5782
rect 8302 5497 8330 5502
rect 8358 5361 8386 5367
rect 8358 5335 8359 5361
rect 8385 5335 8386 5361
rect 8134 5193 8162 5199
rect 8134 5167 8135 5193
rect 8161 5167 8162 5193
rect 8134 4858 8162 5167
rect 8134 4825 8162 4830
rect 8302 4802 8330 4807
rect 8078 4410 8106 4415
rect 8190 4410 8218 4415
rect 8078 4409 8218 4410
rect 8078 4383 8079 4409
rect 8105 4383 8191 4409
rect 8217 4383 8218 4409
rect 8078 4382 8218 4383
rect 8078 4377 8106 4382
rect 8078 4074 8106 4079
rect 8078 4027 8106 4046
rect 8078 3794 8106 3799
rect 8078 3747 8106 3766
rect 7994 3318 8050 3346
rect 8078 3346 8106 3351
rect 7966 3313 7994 3318
rect 7182 3257 7210 3262
rect 7462 3290 7490 3295
rect 8078 3290 8106 3318
rect 7462 3243 7490 3262
rect 8022 3289 8106 3290
rect 8022 3263 8079 3289
rect 8105 3263 8106 3289
rect 8022 3262 8106 3263
rect 7518 3010 7546 3015
rect 7518 2963 7546 2982
rect 7182 2954 7210 2959
rect 7070 2842 7098 2847
rect 7070 2795 7098 2814
rect 7182 2674 7210 2926
rect 7462 2954 7490 2959
rect 7238 2842 7266 2847
rect 7238 2795 7266 2814
rect 7238 2674 7266 2679
rect 7182 2673 7266 2674
rect 7182 2647 7239 2673
rect 7265 2647 7266 2673
rect 7182 2646 7266 2647
rect 7070 2505 7098 2511
rect 7070 2479 7071 2505
rect 7097 2479 7098 2505
rect 7070 2226 7098 2479
rect 7070 2193 7098 2198
rect 7126 2226 7154 2231
rect 7182 2226 7210 2646
rect 7238 2641 7266 2646
rect 7126 2225 7210 2226
rect 7126 2199 7127 2225
rect 7153 2199 7210 2225
rect 7126 2198 7210 2199
rect 7126 2193 7154 2198
rect 6734 1806 6930 1834
rect 7014 2058 7042 2063
rect 7014 1834 7042 2030
rect 7294 2058 7322 2063
rect 7294 2011 7322 2030
rect 6734 937 6762 1806
rect 7014 1801 7042 1806
rect 6958 1778 6986 1783
rect 6790 1777 6986 1778
rect 6790 1751 6959 1777
rect 6985 1751 6986 1777
rect 6790 1750 6986 1751
rect 6790 1721 6818 1750
rect 6958 1745 6986 1750
rect 6790 1695 6791 1721
rect 6817 1695 6818 1721
rect 6790 1050 6818 1695
rect 7238 1722 7266 1727
rect 7238 1675 7266 1694
rect 6846 1666 6874 1671
rect 6846 1442 6874 1638
rect 7294 1666 7322 1671
rect 6846 1441 7042 1442
rect 6846 1415 6847 1441
rect 6873 1415 7042 1441
rect 6846 1414 7042 1415
rect 6846 1409 6874 1414
rect 7014 1385 7042 1414
rect 7294 1441 7322 1638
rect 7294 1415 7295 1441
rect 7321 1415 7322 1441
rect 7294 1409 7322 1415
rect 7014 1359 7015 1385
rect 7041 1359 7042 1385
rect 7014 1353 7042 1359
rect 6790 1017 6818 1022
rect 7406 1050 7434 1055
rect 7406 1003 7434 1022
rect 6958 994 6986 999
rect 6958 993 7098 994
rect 6958 967 6959 993
rect 6985 967 7098 993
rect 6958 966 7098 967
rect 6958 961 6986 966
rect 6734 911 6735 937
rect 6761 911 6762 937
rect 6734 905 6762 911
rect 3598 401 3626 406
rect 3822 882 3850 887
rect 3822 56 3850 854
rect 5166 826 5194 831
rect 4494 322 4522 327
rect 4494 56 4522 294
rect 5166 56 5194 798
rect 6958 826 6986 831
rect 6342 770 6370 775
rect 5558 658 5586 663
rect 5558 611 5586 630
rect 6342 657 6370 742
rect 6342 631 6343 657
rect 6369 631 6370 657
rect 6342 625 6370 631
rect 6510 601 6538 607
rect 6510 575 6511 601
rect 6537 575 6538 601
rect 5782 490 5810 495
rect 5894 490 5922 495
rect 5782 489 5922 490
rect 5782 463 5783 489
rect 5809 463 5895 489
rect 5921 463 5922 489
rect 5782 462 5922 463
rect 5782 457 5810 462
rect 5838 56 5866 462
rect 5894 457 5922 462
rect 6510 490 6538 575
rect 6678 490 6706 495
rect 6510 489 6706 490
rect 6510 463 6679 489
rect 6705 463 6706 489
rect 6510 462 6706 463
rect 6510 56 6538 462
rect 6678 457 6706 462
rect 6958 489 6986 798
rect 7070 658 7098 966
rect 7126 993 7154 999
rect 7126 967 7127 993
rect 7153 967 7154 993
rect 7126 826 7154 967
rect 7126 793 7154 798
rect 7462 658 7490 2926
rect 8022 2674 8050 3262
rect 8078 3257 8106 3262
rect 8022 2641 8050 2646
rect 8134 2954 8162 2959
rect 8078 2618 8106 2623
rect 8078 2571 8106 2590
rect 7518 2562 7546 2567
rect 7518 2515 7546 2534
rect 7630 2562 7658 2567
rect 7798 2562 7826 2567
rect 7630 2561 7826 2562
rect 7630 2535 7631 2561
rect 7657 2535 7799 2561
rect 7825 2535 7826 2561
rect 7630 2534 7826 2535
rect 7630 2282 7658 2534
rect 7798 2529 7826 2534
rect 7630 2249 7658 2254
rect 7518 2225 7546 2231
rect 7518 2199 7519 2225
rect 7545 2199 7546 2225
rect 7518 2114 7546 2199
rect 8134 2225 8162 2926
rect 8190 2506 8218 4382
rect 8190 2473 8218 2478
rect 8246 3738 8274 3743
rect 8134 2199 8135 2225
rect 8161 2199 8162 2225
rect 8134 2193 8162 2199
rect 7518 2081 7546 2086
rect 7686 2058 7714 2063
rect 7854 2058 7882 2063
rect 7686 2057 7882 2058
rect 7686 2031 7687 2057
rect 7713 2031 7855 2057
rect 7881 2031 7882 2057
rect 7686 2030 7882 2031
rect 7686 2002 7714 2030
rect 7854 2025 7882 2030
rect 7686 1969 7714 1974
rect 8022 1721 8050 1727
rect 8022 1695 8023 1721
rect 8049 1695 8050 1721
rect 7518 1386 7546 1391
rect 7518 1339 7546 1358
rect 7686 1386 7714 1391
rect 7686 1339 7714 1358
rect 7966 1329 7994 1335
rect 7966 1303 7967 1329
rect 7993 1303 7994 1329
rect 7966 1106 7994 1303
rect 8022 1274 8050 1695
rect 8022 1241 8050 1246
rect 8078 1442 8106 1447
rect 7966 1073 7994 1078
rect 8078 1049 8106 1414
rect 8134 1274 8162 1279
rect 8134 1227 8162 1246
rect 8078 1023 8079 1049
rect 8105 1023 8106 1049
rect 8078 1017 8106 1023
rect 7798 993 7826 999
rect 7798 967 7799 993
rect 7825 967 7826 993
rect 7630 938 7658 943
rect 7798 938 7826 967
rect 7630 937 7826 938
rect 7630 911 7631 937
rect 7657 911 7826 937
rect 7630 910 7826 911
rect 7630 714 7658 910
rect 8246 770 8274 3710
rect 8302 3010 8330 4774
rect 8358 4466 8386 5335
rect 8806 5361 8834 6286
rect 8862 6202 8890 6399
rect 8974 6426 9002 7056
rect 9086 6594 9114 7056
rect 9198 6706 9226 7056
rect 9198 6673 9226 6678
rect 9254 6594 9282 6599
rect 9086 6593 9282 6594
rect 9086 6567 9255 6593
rect 9281 6567 9282 6593
rect 9086 6566 9282 6567
rect 9086 6481 9114 6566
rect 9254 6561 9282 6566
rect 9086 6455 9087 6481
rect 9113 6455 9114 6481
rect 9086 6449 9114 6455
rect 9310 6482 9338 7056
rect 9422 6930 9450 7056
rect 9422 6902 9506 6930
rect 9478 6762 9506 6902
rect 9310 6449 9338 6454
rect 9422 6734 9506 6762
rect 8974 6393 9002 6398
rect 9422 6370 9450 6734
rect 9478 6650 9506 6655
rect 9478 6593 9506 6622
rect 9478 6567 9479 6593
rect 9505 6567 9506 6593
rect 9478 6561 9506 6567
rect 9310 6342 9450 6370
rect 8862 6169 8890 6174
rect 9198 6314 9226 6319
rect 8974 6090 9002 6095
rect 8974 6043 9002 6062
rect 9142 6090 9170 6095
rect 9142 5809 9170 6062
rect 9198 6034 9226 6286
rect 9254 6146 9282 6151
rect 9254 6099 9282 6118
rect 9198 6006 9282 6034
rect 9142 5783 9143 5809
rect 9169 5783 9170 5809
rect 9142 5777 9170 5783
rect 9086 5754 9114 5759
rect 8806 5335 8807 5361
rect 8833 5335 8834 5361
rect 8806 5329 8834 5335
rect 9030 5642 9058 5647
rect 8358 4433 8386 4438
rect 8414 5138 8442 5143
rect 8414 3794 8442 5110
rect 8470 4465 8498 4471
rect 8470 4439 8471 4465
rect 8497 4439 8498 4465
rect 8470 4130 8498 4439
rect 8470 4097 8498 4102
rect 9030 3906 9058 5614
rect 9086 5306 9114 5726
rect 9254 5474 9282 6006
rect 9310 5586 9338 6342
rect 9534 6314 9562 7056
rect 9646 6370 9674 7056
rect 9534 6281 9562 6286
rect 9590 6342 9674 6370
rect 9702 6425 9730 6431
rect 9702 6399 9703 6425
rect 9729 6399 9730 6425
rect 9702 6370 9730 6399
rect 9590 6146 9618 6342
rect 9702 6337 9730 6342
rect 9478 6145 9618 6146
rect 9478 6119 9591 6145
rect 9617 6119 9618 6145
rect 9478 6118 9618 6119
rect 9478 6089 9506 6118
rect 9590 6113 9618 6118
rect 9478 6063 9479 6089
rect 9505 6063 9506 6089
rect 9478 6057 9506 6063
rect 9758 6090 9786 7056
rect 9758 6062 9842 6090
rect 9366 5978 9394 5983
rect 9366 5698 9394 5950
rect 9758 5977 9786 5983
rect 9758 5951 9759 5977
rect 9785 5951 9786 5977
rect 9534 5922 9562 5927
rect 9534 5809 9562 5894
rect 9758 5922 9786 5951
rect 9758 5889 9786 5894
rect 9534 5783 9535 5809
rect 9561 5783 9562 5809
rect 9534 5777 9562 5783
rect 9814 5754 9842 6062
rect 9814 5721 9842 5726
rect 9422 5698 9450 5703
rect 9366 5697 9450 5698
rect 9366 5671 9423 5697
rect 9449 5671 9450 5697
rect 9366 5670 9450 5671
rect 9422 5665 9450 5670
rect 9758 5697 9786 5703
rect 9758 5671 9759 5697
rect 9785 5671 9786 5697
rect 9646 5642 9674 5647
rect 9758 5642 9786 5671
rect 9646 5641 9786 5642
rect 9646 5615 9647 5641
rect 9673 5615 9786 5641
rect 9646 5614 9786 5615
rect 9646 5586 9674 5614
rect 9310 5553 9338 5558
rect 9478 5558 9674 5586
rect 9366 5530 9394 5535
rect 9254 5446 9338 5474
rect 9086 5305 9226 5306
rect 9086 5279 9087 5305
rect 9113 5279 9226 5305
rect 9086 5278 9226 5279
rect 9086 5273 9114 5278
rect 9198 5138 9226 5278
rect 9254 5250 9282 5255
rect 9254 5203 9282 5222
rect 9198 5110 9282 5138
rect 9254 5025 9282 5110
rect 9254 4999 9255 5025
rect 9281 4999 9282 5025
rect 9254 4993 9282 4999
rect 9030 3873 9058 3878
rect 9310 3850 9338 5446
rect 9310 3817 9338 3822
rect 8414 3761 8442 3766
rect 8918 3682 8946 3687
rect 8358 3346 8386 3351
rect 8358 3299 8386 3318
rect 8302 2977 8330 2982
rect 8638 3289 8666 3295
rect 8638 3263 8639 3289
rect 8665 3263 8666 3289
rect 8414 2561 8442 2567
rect 8414 2535 8415 2561
rect 8441 2535 8442 2561
rect 8302 2170 8330 2175
rect 8414 2170 8442 2535
rect 8330 2142 8442 2170
rect 8638 2170 8666 3263
rect 8750 2730 8778 2735
rect 8694 2674 8722 2679
rect 8694 2617 8722 2646
rect 8694 2591 8695 2617
rect 8721 2591 8722 2617
rect 8694 2585 8722 2591
rect 8750 2225 8778 2702
rect 8862 2730 8890 2735
rect 8862 2673 8890 2702
rect 8862 2647 8863 2673
rect 8889 2647 8890 2673
rect 8862 2641 8890 2647
rect 8750 2199 8751 2225
rect 8777 2199 8778 2225
rect 8750 2193 8778 2199
rect 8302 2123 8330 2142
rect 8638 2137 8666 2142
rect 8638 1498 8666 1503
rect 8358 1441 8386 1447
rect 8358 1415 8359 1441
rect 8385 1415 8386 1441
rect 8358 1386 8386 1415
rect 8638 1386 8666 1470
rect 8918 1441 8946 3654
rect 9198 3458 9226 3463
rect 9142 2842 9170 2847
rect 9142 2617 9170 2814
rect 9142 2591 9143 2617
rect 9169 2591 9170 2617
rect 9142 2585 9170 2591
rect 8918 1415 8919 1441
rect 8945 1415 8946 1441
rect 8918 1409 8946 1415
rect 8358 1353 8386 1358
rect 8526 1385 8666 1386
rect 8526 1359 8639 1385
rect 8665 1359 8666 1385
rect 8526 1358 8666 1359
rect 8526 1105 8554 1358
rect 8638 1353 8666 1358
rect 8526 1079 8527 1105
rect 8553 1079 8554 1105
rect 8526 1073 8554 1079
rect 9142 938 9170 943
rect 9142 891 9170 910
rect 8246 737 8274 742
rect 7630 681 7658 686
rect 7070 657 7210 658
rect 7070 631 7071 657
rect 7097 631 7210 657
rect 7070 630 7210 631
rect 7070 625 7098 630
rect 6958 463 6959 489
rect 6985 463 6986 489
rect 6958 154 6986 463
rect 6958 121 6986 126
rect 7182 56 7210 630
rect 7462 625 7490 630
rect 8134 658 8162 663
rect 7854 602 7882 607
rect 7854 555 7882 574
rect 8134 546 8162 630
rect 8134 499 8162 518
rect 8358 657 8386 663
rect 8358 631 8359 657
rect 8385 631 8386 657
rect 8358 546 8386 631
rect 8526 658 8554 663
rect 8526 611 8554 630
rect 9198 657 9226 3430
rect 9310 993 9338 999
rect 9310 967 9311 993
rect 9337 967 9338 993
rect 9310 938 9338 967
rect 9310 905 9338 910
rect 9198 631 9199 657
rect 9225 631 9226 657
rect 9198 625 9226 631
rect 8358 513 8386 518
rect 7462 490 7490 495
rect 7574 490 7602 495
rect 7462 489 7602 490
rect 7462 463 7463 489
rect 7489 463 7575 489
rect 7601 463 7602 489
rect 7462 462 7602 463
rect 7462 266 7490 462
rect 7574 457 7602 462
rect 7854 490 7882 495
rect 7462 233 7490 238
rect 7854 56 7882 462
rect 8806 490 8834 495
rect 8806 443 8834 462
rect 8918 490 8946 495
rect 8918 443 8946 462
rect 8526 378 8554 383
rect 8526 56 8554 350
rect 9366 322 9394 5502
rect 9478 1890 9506 5558
rect 9870 5530 9898 7056
rect 9534 5502 9898 5530
rect 9926 6034 9954 6039
rect 9534 5305 9562 5502
rect 9534 5279 9535 5305
rect 9561 5279 9562 5305
rect 9534 5273 9562 5279
rect 9702 5025 9730 5502
rect 9926 5474 9954 6006
rect 9814 5446 9954 5474
rect 9814 5361 9842 5446
rect 9814 5335 9815 5361
rect 9841 5335 9842 5361
rect 9814 5329 9842 5335
rect 9982 5418 10010 7056
rect 10038 6258 10066 6263
rect 10038 6145 10066 6230
rect 10038 6119 10039 6145
rect 10065 6119 10066 6145
rect 10038 6113 10066 6119
rect 9982 5305 10010 5390
rect 9982 5279 9983 5305
rect 10009 5279 10010 5305
rect 9982 5273 10010 5279
rect 10038 5641 10066 5647
rect 10038 5615 10039 5641
rect 10065 5615 10066 5641
rect 9702 4999 9703 5025
rect 9729 4999 9730 5025
rect 9702 4993 9730 4999
rect 9926 5082 9954 5087
rect 9478 1857 9506 1862
rect 9590 4298 9618 4303
rect 9590 1049 9618 4270
rect 9926 3962 9954 5054
rect 10038 4634 10066 5615
rect 10094 5586 10122 7056
rect 10150 5978 10178 5983
rect 10150 5698 10178 5950
rect 10206 5810 10234 7056
rect 10262 6762 10290 6767
rect 10262 5978 10290 6734
rect 10262 5945 10290 5950
rect 10318 5866 10346 7056
rect 10430 6874 10458 7056
rect 10374 6846 10458 6874
rect 10374 5978 10402 6846
rect 10430 6762 10458 6767
rect 10430 6201 10458 6734
rect 10430 6175 10431 6201
rect 10457 6175 10458 6201
rect 10430 6169 10458 6175
rect 10486 6425 10514 6431
rect 10486 6399 10487 6425
rect 10513 6399 10514 6425
rect 10486 6090 10514 6399
rect 10542 6426 10570 7056
rect 10542 6393 10570 6398
rect 10486 6057 10514 6062
rect 10542 6034 10570 6039
rect 10374 5950 10514 5978
rect 10430 5866 10458 5871
rect 10318 5838 10430 5866
rect 10430 5833 10458 5838
rect 10206 5782 10402 5810
rect 10206 5698 10234 5703
rect 10150 5697 10234 5698
rect 10150 5671 10207 5697
rect 10233 5671 10234 5697
rect 10150 5670 10234 5671
rect 10206 5665 10234 5670
rect 10094 5553 10122 5558
rect 10150 5418 10178 5423
rect 10150 5025 10178 5390
rect 10374 5306 10402 5782
rect 10486 5754 10514 5950
rect 10430 5726 10514 5754
rect 10430 5698 10458 5726
rect 10430 5665 10458 5670
rect 10486 5642 10514 5647
rect 10486 5595 10514 5614
rect 10318 5194 10346 5199
rect 10150 4999 10151 5025
rect 10177 4999 10178 5025
rect 10150 4993 10178 4999
rect 10262 5193 10346 5194
rect 10262 5167 10319 5193
rect 10345 5167 10346 5193
rect 10262 5166 10346 5167
rect 10038 4601 10066 4606
rect 9926 3929 9954 3934
rect 9590 1023 9591 1049
rect 9617 1023 9618 1049
rect 9590 1017 9618 1023
rect 10038 3850 10066 3855
rect 9814 993 9842 999
rect 9814 967 9815 993
rect 9841 967 9842 993
rect 9814 602 9842 967
rect 10038 937 10066 3822
rect 10206 994 10234 999
rect 10206 947 10234 966
rect 10038 911 10039 937
rect 10065 911 10066 937
rect 10038 905 10066 911
rect 9702 574 9842 602
rect 9366 289 9394 294
rect 9646 490 9674 495
rect 9702 490 9730 574
rect 10206 546 10234 551
rect 10262 546 10290 5166
rect 10318 5161 10346 5166
rect 10318 5026 10346 5031
rect 10374 5026 10402 5278
rect 10318 5025 10402 5026
rect 10318 4999 10319 5025
rect 10345 4999 10402 5025
rect 10318 4998 10402 4999
rect 10430 5586 10458 5591
rect 10430 5026 10458 5558
rect 10486 5250 10514 5255
rect 10542 5250 10570 6006
rect 10654 5642 10682 7056
rect 10766 6034 10794 7056
rect 10878 6594 10906 7056
rect 10990 6650 11018 7056
rect 10990 6617 11018 6622
rect 10878 6561 10906 6566
rect 11102 6538 11130 7056
rect 11102 6505 11130 6510
rect 10766 6001 10794 6006
rect 10822 6481 10850 6487
rect 10822 6455 10823 6481
rect 10849 6455 10850 6481
rect 10710 5978 10738 5983
rect 10710 5809 10738 5950
rect 10710 5783 10711 5809
rect 10737 5783 10738 5809
rect 10710 5777 10738 5783
rect 10766 5922 10794 5927
rect 10654 5609 10682 5614
rect 10654 5306 10682 5311
rect 10654 5259 10682 5278
rect 10486 5249 10570 5250
rect 10486 5223 10487 5249
rect 10513 5223 10570 5249
rect 10486 5222 10570 5223
rect 10486 5217 10514 5222
rect 10542 5026 10570 5031
rect 10430 5025 10570 5026
rect 10430 4999 10431 5025
rect 10457 4999 10543 5025
rect 10569 4999 10570 5025
rect 10430 4998 10570 4999
rect 10318 4993 10346 4998
rect 10430 4993 10458 4998
rect 10542 4993 10570 4998
rect 10766 4970 10794 5894
rect 10822 5026 10850 6455
rect 10990 6481 11018 6487
rect 10990 6455 10991 6481
rect 11017 6455 11018 6481
rect 10878 6370 10906 6375
rect 10878 5922 10906 6342
rect 10878 5889 10906 5894
rect 10934 6033 10962 6039
rect 10934 6007 10935 6033
rect 10961 6007 10962 6033
rect 10934 5641 10962 6007
rect 10934 5615 10935 5641
rect 10961 5615 10962 5641
rect 10934 5609 10962 5615
rect 10990 5418 11018 6455
rect 11102 6034 11130 6039
rect 10934 5390 11018 5418
rect 11046 6033 11130 6034
rect 11046 6007 11103 6033
rect 11129 6007 11130 6033
rect 11046 6006 11130 6007
rect 10822 4993 10850 4998
rect 10878 5361 10906 5367
rect 10878 5335 10879 5361
rect 10905 5335 10906 5361
rect 10710 4942 10794 4970
rect 10654 4410 10682 4415
rect 10654 2450 10682 4382
rect 10654 2417 10682 2422
rect 10710 1694 10738 4942
rect 10878 4914 10906 5335
rect 10878 4881 10906 4886
rect 10766 4857 10794 4863
rect 10766 4831 10767 4857
rect 10793 4831 10794 4857
rect 10766 4018 10794 4831
rect 10934 4298 10962 5390
rect 10990 5306 11018 5311
rect 10990 5025 11018 5278
rect 10990 4999 10991 5025
rect 11017 4999 11018 5025
rect 10990 4993 11018 4999
rect 10934 4265 10962 4270
rect 10766 3985 10794 3990
rect 11046 3850 11074 6006
rect 11102 6001 11130 6006
rect 11102 5922 11130 5927
rect 11102 5809 11130 5894
rect 11102 5783 11103 5809
rect 11129 5783 11130 5809
rect 11102 5777 11130 5783
rect 11158 5866 11186 5871
rect 11158 5306 11186 5838
rect 11214 5810 11242 7056
rect 11270 6594 11298 6599
rect 11270 6547 11298 6566
rect 11326 6202 11354 7056
rect 11326 6169 11354 6174
rect 11382 6650 11410 6655
rect 11382 6201 11410 6622
rect 11382 6175 11383 6201
rect 11409 6175 11410 6201
rect 11382 6169 11410 6175
rect 11214 5777 11242 5782
rect 11326 5698 11354 5703
rect 11158 5273 11186 5278
rect 11214 5697 11354 5698
rect 11214 5671 11327 5697
rect 11353 5671 11354 5697
rect 11214 5670 11354 5671
rect 11046 3817 11074 3822
rect 11102 5250 11130 5255
rect 11102 3458 11130 5222
rect 11158 5194 11186 5199
rect 11158 4857 11186 5166
rect 11158 4831 11159 4857
rect 11185 4831 11186 4857
rect 11158 4825 11186 4831
rect 11102 3425 11130 3430
rect 10878 1834 10906 1839
rect 10710 1666 10794 1694
rect 10710 1274 10738 1279
rect 10710 1227 10738 1246
rect 10598 1162 10626 1167
rect 10374 994 10402 999
rect 10374 947 10402 966
rect 10206 545 10290 546
rect 10206 519 10207 545
rect 10233 519 10290 545
rect 10206 518 10290 519
rect 10206 513 10234 518
rect 9814 490 9842 495
rect 10038 490 10066 495
rect 9646 489 9730 490
rect 9646 463 9647 489
rect 9673 463 9730 489
rect 9646 462 9730 463
rect 9758 489 10066 490
rect 9758 463 9815 489
rect 9841 463 10039 489
rect 10065 463 10066 489
rect 9758 462 10066 463
rect 9198 266 9226 271
rect 9198 56 9226 238
rect 9646 98 9674 462
rect 9646 65 9674 70
rect 1120 0 1176 56
rect 1792 0 1848 56
rect 2464 0 2520 56
rect 3136 0 3192 56
rect 3808 0 3864 56
rect 4480 0 4536 56
rect 5152 0 5208 56
rect 5824 0 5880 56
rect 6496 0 6552 56
rect 7168 0 7224 56
rect 7840 0 7896 56
rect 8512 0 8568 56
rect 9184 0 9240 56
rect 9758 42 9786 462
rect 9814 457 9842 462
rect 10038 457 10066 462
rect 10430 490 10458 495
rect 10542 490 10570 495
rect 10430 489 10570 490
rect 10430 463 10431 489
rect 10457 463 10543 489
rect 10569 463 10570 489
rect 10430 462 10570 463
rect 9870 322 9898 327
rect 9870 56 9898 294
rect 10430 322 10458 462
rect 10542 457 10570 462
rect 10598 378 10626 1134
rect 10654 1050 10682 1055
rect 10766 1050 10794 1666
rect 10654 1049 10794 1050
rect 10654 1023 10655 1049
rect 10681 1023 10794 1049
rect 10654 1022 10794 1023
rect 10822 1274 10850 1279
rect 10654 1017 10682 1022
rect 10822 993 10850 1246
rect 10822 967 10823 993
rect 10849 967 10850 993
rect 10822 882 10850 967
rect 10822 849 10850 854
rect 10822 658 10850 663
rect 10878 658 10906 1806
rect 11214 1694 11242 5670
rect 11326 5665 11354 5670
rect 11438 5418 11466 7056
rect 11550 6930 11578 7056
rect 11550 6897 11578 6902
rect 11662 6482 11690 7056
rect 11662 6449 11690 6454
rect 11606 5810 11634 5815
rect 11606 5763 11634 5782
rect 11550 5754 11578 5759
rect 11438 5385 11466 5390
rect 11494 5698 11522 5703
rect 11326 5362 11354 5367
rect 11326 5315 11354 5334
rect 11494 5026 11522 5670
rect 11550 5305 11578 5726
rect 11774 5642 11802 7056
rect 11886 6370 11914 7056
rect 11998 6594 12026 7056
rect 11998 6561 12026 6566
rect 11774 5609 11802 5614
rect 11830 6342 11914 6370
rect 11942 6481 11970 6487
rect 11942 6455 11943 6481
rect 11969 6455 11970 6481
rect 11942 6370 11970 6455
rect 11830 5586 11858 6342
rect 11942 6337 11970 6342
rect 11902 6286 12034 6291
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 11902 6253 12034 6258
rect 11998 6202 12026 6207
rect 11998 6155 12026 6174
rect 11830 5553 11858 5558
rect 11902 5502 12034 5507
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 11902 5469 12034 5474
rect 12110 5474 12138 7056
rect 12222 6818 12250 7056
rect 12334 6874 12362 7056
rect 12334 6841 12362 6846
rect 12222 6785 12250 6790
rect 12232 6678 12364 6683
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12232 6645 12364 6650
rect 12222 6593 12250 6599
rect 12222 6567 12223 6593
rect 12249 6567 12250 6593
rect 12222 6538 12250 6567
rect 12222 6505 12250 6510
rect 12110 5441 12138 5446
rect 12166 6426 12194 6431
rect 11830 5418 11858 5423
rect 11830 5371 11858 5390
rect 11550 5279 11551 5305
rect 11577 5279 11578 5305
rect 11550 5273 11578 5279
rect 11774 5306 11802 5311
rect 11774 5082 11802 5278
rect 11774 5049 11802 5054
rect 11550 5026 11578 5031
rect 11270 5025 11578 5026
rect 11270 4999 11551 5025
rect 11577 4999 11578 5025
rect 11270 4998 11578 4999
rect 11270 4577 11298 4998
rect 11550 4993 11578 4998
rect 11718 5026 11746 5031
rect 11382 4913 11410 4919
rect 11382 4887 11383 4913
rect 11409 4887 11410 4913
rect 11382 4858 11410 4887
rect 11382 4825 11410 4830
rect 11606 4914 11634 4919
rect 11718 4914 11746 4998
rect 11718 4886 11802 4914
rect 11270 4551 11271 4577
rect 11297 4551 11298 4577
rect 11270 4545 11298 4551
rect 11326 4410 11354 4415
rect 11494 4410 11522 4415
rect 11354 4409 11522 4410
rect 11354 4383 11495 4409
rect 11521 4383 11522 4409
rect 11354 4382 11522 4383
rect 11326 4363 11354 4382
rect 11494 4377 11522 4382
rect 11550 4410 11578 4415
rect 11102 1666 11242 1694
rect 11102 1049 11130 1666
rect 11102 1023 11103 1049
rect 11129 1023 11130 1049
rect 11102 1017 11130 1023
rect 11326 993 11354 999
rect 11326 967 11327 993
rect 11353 967 11354 993
rect 10822 657 10906 658
rect 10822 631 10823 657
rect 10849 631 10906 657
rect 10822 630 10906 631
rect 11214 938 11242 943
rect 10822 625 10850 630
rect 10430 289 10458 294
rect 10542 350 10626 378
rect 11102 490 11130 495
rect 10542 56 10570 350
rect 11102 266 11130 462
rect 11158 489 11186 495
rect 11158 463 11159 489
rect 11185 463 11186 489
rect 11158 378 11186 463
rect 11158 345 11186 350
rect 11102 233 11130 238
rect 11214 56 11242 910
rect 11326 378 11354 967
rect 11550 937 11578 4382
rect 11550 911 11551 937
rect 11577 911 11578 937
rect 11550 905 11578 911
rect 11606 657 11634 4886
rect 11662 4858 11690 4863
rect 11662 4410 11690 4830
rect 11774 4577 11802 4886
rect 11774 4551 11775 4577
rect 11801 4551 11802 4577
rect 11774 4545 11802 4551
rect 11830 4857 11858 4863
rect 11830 4831 11831 4857
rect 11857 4831 11858 4857
rect 11662 4382 11802 4410
rect 11774 1386 11802 4382
rect 11830 4354 11858 4831
rect 11942 4858 11970 4863
rect 11942 4811 11970 4830
rect 11902 4718 12034 4723
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12166 4690 12194 6398
rect 12232 5894 12364 5899
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12232 5861 12364 5866
rect 12446 5754 12474 7056
rect 12558 6370 12586 7056
rect 12558 6337 12586 6342
rect 12670 6202 12698 7056
rect 12726 6481 12754 6487
rect 12726 6455 12727 6481
rect 12753 6455 12754 6481
rect 12726 6426 12754 6455
rect 12726 6393 12754 6398
rect 12670 6169 12698 6174
rect 12726 6314 12754 6319
rect 12502 6034 12530 6039
rect 12502 5987 12530 6006
rect 12670 6033 12698 6039
rect 12670 6007 12671 6033
rect 12697 6007 12698 6033
rect 12670 5866 12698 6007
rect 12670 5833 12698 5838
rect 12446 5726 12698 5754
rect 12278 5697 12306 5703
rect 12278 5671 12279 5697
rect 12305 5671 12306 5697
rect 12278 5306 12306 5671
rect 12558 5642 12586 5647
rect 12558 5595 12586 5614
rect 12614 5586 12642 5591
rect 12278 5273 12306 5278
rect 12558 5474 12586 5479
rect 12334 5250 12362 5255
rect 12334 5203 12362 5222
rect 12232 5110 12364 5115
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12232 5077 12364 5082
rect 12558 5025 12586 5446
rect 12614 5417 12642 5558
rect 12614 5391 12615 5417
rect 12641 5391 12642 5417
rect 12614 5385 12642 5391
rect 12558 4999 12559 5025
rect 12585 4999 12586 5025
rect 12558 4993 12586 4999
rect 12614 5026 12642 5031
rect 12278 4914 12306 4919
rect 12278 4867 12306 4886
rect 11902 4685 12034 4690
rect 12110 4662 12194 4690
rect 12110 4634 12138 4662
rect 11998 4606 12138 4634
rect 12446 4634 12474 4639
rect 11998 4521 12026 4606
rect 11998 4495 11999 4521
rect 12025 4495 12026 4521
rect 11998 4489 12026 4495
rect 12166 4577 12194 4583
rect 12166 4551 12167 4577
rect 12193 4551 12194 4577
rect 11942 4410 11970 4415
rect 11830 4321 11858 4326
rect 11886 4409 11970 4410
rect 11886 4383 11943 4409
rect 11969 4383 11970 4409
rect 11886 4382 11970 4383
rect 11830 4242 11858 4247
rect 11886 4242 11914 4382
rect 11942 4377 11970 4382
rect 11830 4241 11914 4242
rect 11830 4215 11831 4241
rect 11857 4215 11914 4241
rect 11830 4214 11914 4215
rect 11830 4209 11858 4214
rect 11902 3934 12034 3939
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 11902 3901 12034 3906
rect 12110 3794 12138 3799
rect 11902 3150 12034 3155
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 11902 3117 12034 3122
rect 11902 2366 12034 2371
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 11902 2333 12034 2338
rect 11902 1582 12034 1587
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 11902 1549 12034 1554
rect 12054 1442 12082 1447
rect 12110 1442 12138 3766
rect 12054 1441 12138 1442
rect 12054 1415 12055 1441
rect 12081 1415 12138 1441
rect 12054 1414 12138 1415
rect 12054 1409 12082 1414
rect 11774 1358 11858 1386
rect 11662 1274 11690 1279
rect 11774 1274 11802 1279
rect 11662 1273 11802 1274
rect 11662 1247 11663 1273
rect 11689 1247 11775 1273
rect 11801 1247 11802 1273
rect 11662 1246 11802 1247
rect 11662 1162 11690 1246
rect 11774 1241 11802 1246
rect 11662 1129 11690 1134
rect 11830 714 11858 1358
rect 11902 798 12034 803
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 11902 765 12034 770
rect 12166 714 12194 4551
rect 12232 4326 12364 4331
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12232 4293 12364 4298
rect 12446 4129 12474 4606
rect 12614 4410 12642 4998
rect 12670 4633 12698 5726
rect 12670 4607 12671 4633
rect 12697 4607 12698 4633
rect 12670 4601 12698 4607
rect 12614 4377 12642 4382
rect 12726 4185 12754 6286
rect 12782 5978 12810 7056
rect 12782 5945 12810 5950
rect 12838 6986 12866 6991
rect 12726 4159 12727 4185
rect 12753 4159 12754 4185
rect 12726 4153 12754 4159
rect 12446 4103 12447 4129
rect 12473 4103 12474 4129
rect 12446 4097 12474 4103
rect 12838 3793 12866 6958
rect 12894 6762 12922 7056
rect 13006 7042 13034 7056
rect 13006 7009 13034 7014
rect 13398 7042 13426 7047
rect 12894 6729 12922 6734
rect 12950 6930 12978 6935
rect 12950 6594 12978 6902
rect 13006 6594 13034 6599
rect 12950 6593 13034 6594
rect 12950 6567 13007 6593
rect 13033 6567 13034 6593
rect 12950 6566 13034 6567
rect 13006 6561 13034 6566
rect 12950 6482 12978 6487
rect 12950 6201 12978 6454
rect 12950 6175 12951 6201
rect 12977 6175 12978 6201
rect 12950 6169 12978 6175
rect 13006 6426 13034 6431
rect 12838 3767 12839 3793
rect 12865 3767 12866 3793
rect 12838 3761 12866 3767
rect 12894 5866 12922 5871
rect 12894 3738 12922 5838
rect 12894 3705 12922 3710
rect 12232 3542 12364 3547
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12232 3509 12364 3514
rect 12950 3514 12978 3519
rect 12232 2758 12364 2763
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12232 2725 12364 2730
rect 12232 1974 12364 1979
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12232 1941 12364 1946
rect 12950 1441 12978 3486
rect 13006 2898 13034 6398
rect 13174 5978 13202 5983
rect 13118 5922 13146 5927
rect 13062 5697 13090 5703
rect 13062 5671 13063 5697
rect 13089 5671 13090 5697
rect 13062 5026 13090 5671
rect 13062 4993 13090 4998
rect 13006 2865 13034 2870
rect 13062 4521 13090 4527
rect 13062 4495 13063 4521
rect 13089 4495 13090 4521
rect 12950 1415 12951 1441
rect 12977 1415 12978 1441
rect 12950 1409 12978 1415
rect 12614 1274 12642 1279
rect 12726 1274 12754 1279
rect 12614 1273 12754 1274
rect 12614 1247 12615 1273
rect 12641 1247 12727 1273
rect 12753 1247 12754 1273
rect 12614 1246 12754 1247
rect 12232 1190 12364 1195
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12232 1157 12364 1162
rect 12558 994 12586 999
rect 12558 947 12586 966
rect 12390 938 12418 943
rect 12390 891 12418 910
rect 12614 882 12642 1246
rect 12726 1241 12754 1246
rect 12838 1050 12866 1055
rect 13062 1050 13090 4495
rect 13118 3737 13146 5894
rect 13174 4857 13202 5950
rect 13398 5754 13426 7014
rect 13510 6874 13538 6879
rect 13454 6425 13482 6431
rect 13454 6399 13455 6425
rect 13481 6399 13482 6425
rect 13454 5977 13482 6399
rect 13454 5951 13455 5977
rect 13481 5951 13482 5977
rect 13454 5866 13482 5951
rect 13454 5833 13482 5838
rect 13398 5726 13482 5754
rect 13174 4831 13175 4857
rect 13201 4831 13202 4857
rect 13174 4825 13202 4831
rect 13230 5305 13258 5311
rect 13230 5279 13231 5305
rect 13257 5279 13258 5305
rect 13230 4242 13258 5279
rect 13454 4633 13482 5726
rect 13510 5361 13538 6846
rect 14126 6818 14154 6823
rect 13566 6594 13594 6599
rect 13566 5641 13594 6566
rect 14126 6593 14154 6790
rect 14126 6567 14127 6593
rect 14153 6567 14154 6593
rect 14126 6561 14154 6567
rect 14910 6762 14938 6767
rect 14910 6593 14938 6734
rect 14910 6567 14911 6593
rect 14937 6567 14938 6593
rect 14910 6561 14938 6567
rect 13790 6538 13818 6543
rect 13734 6034 13762 6039
rect 13734 5987 13762 6006
rect 13678 5866 13706 5871
rect 13566 5615 13567 5641
rect 13593 5615 13594 5641
rect 13566 5609 13594 5615
rect 13622 5642 13650 5647
rect 13510 5335 13511 5361
rect 13537 5335 13538 5361
rect 13510 5329 13538 5335
rect 13454 4607 13455 4633
rect 13481 4607 13482 4633
rect 13454 4601 13482 4607
rect 13566 4913 13594 4919
rect 13566 4887 13567 4913
rect 13593 4887 13594 4913
rect 13174 4214 13258 4242
rect 13174 3794 13202 4214
rect 13174 3761 13202 3766
rect 13230 4129 13258 4135
rect 13230 4103 13231 4129
rect 13257 4103 13258 4129
rect 13118 3711 13119 3737
rect 13145 3711 13146 3737
rect 13118 3705 13146 3711
rect 13118 3402 13146 3407
rect 13118 3355 13146 3374
rect 13230 2954 13258 4103
rect 13342 3682 13370 3687
rect 13342 3635 13370 3654
rect 13230 2921 13258 2926
rect 13566 1833 13594 4887
rect 13622 4073 13650 5614
rect 13622 4047 13623 4073
rect 13649 4047 13650 4073
rect 13622 4041 13650 4047
rect 13678 3793 13706 5838
rect 13790 4214 13818 6510
rect 13958 6482 13986 6487
rect 14630 6482 14658 6487
rect 13958 6481 14210 6482
rect 13958 6455 13959 6481
rect 13985 6455 14210 6481
rect 13958 6454 14210 6455
rect 13958 6449 13986 6454
rect 14126 6370 14154 6375
rect 13958 5978 13986 5983
rect 13846 5698 13874 5703
rect 13846 5361 13874 5670
rect 13846 5335 13847 5361
rect 13873 5335 13874 5361
rect 13846 5306 13874 5335
rect 13846 5273 13874 5278
rect 13902 5697 13930 5703
rect 13902 5671 13903 5697
rect 13929 5671 13930 5697
rect 13902 5194 13930 5671
rect 13902 5161 13930 5166
rect 13958 5082 13986 5950
rect 14126 5809 14154 6342
rect 14126 5783 14127 5809
rect 14153 5783 14154 5809
rect 14126 5777 14154 5783
rect 13678 3767 13679 3793
rect 13705 3767 13706 3793
rect 13678 3761 13706 3767
rect 13734 4186 13818 4214
rect 13846 5054 13986 5082
rect 14014 5193 14042 5199
rect 14014 5167 14015 5193
rect 14041 5167 14042 5193
rect 13734 3682 13762 4186
rect 13622 3654 13762 3682
rect 13622 3289 13650 3654
rect 13622 3263 13623 3289
rect 13649 3263 13650 3289
rect 13622 3257 13650 3263
rect 13846 3066 13874 5054
rect 13902 4913 13930 4919
rect 13902 4887 13903 4913
rect 13929 4887 13930 4913
rect 13902 4802 13930 4887
rect 13902 4769 13930 4774
rect 14014 4522 14042 5167
rect 14014 4489 14042 4494
rect 13958 4465 13986 4471
rect 13958 4439 13959 4465
rect 13985 4439 13986 4465
rect 13902 3345 13930 3351
rect 13902 3319 13903 3345
rect 13929 3319 13930 3345
rect 13902 3290 13930 3319
rect 13902 3257 13930 3262
rect 13846 3033 13874 3038
rect 13902 2674 13930 2679
rect 13902 2617 13930 2646
rect 13902 2591 13903 2617
rect 13929 2591 13930 2617
rect 13902 2585 13930 2591
rect 13566 1807 13567 1833
rect 13593 1807 13594 1833
rect 13566 1801 13594 1807
rect 13902 2114 13930 2119
rect 13902 1833 13930 2086
rect 13902 1807 13903 1833
rect 13929 1807 13930 1833
rect 13902 1801 13930 1807
rect 13286 1778 13314 1783
rect 13286 1694 13314 1750
rect 13678 1778 13706 1783
rect 13678 1731 13706 1750
rect 13230 1666 13314 1694
rect 13846 1722 13874 1727
rect 12838 1049 13090 1050
rect 12838 1023 12839 1049
rect 12865 1023 13090 1049
rect 12838 1022 13090 1023
rect 13118 1442 13146 1447
rect 13118 1049 13146 1414
rect 13118 1023 13119 1049
rect 13145 1023 13146 1049
rect 12838 1017 12866 1022
rect 13118 1017 13146 1023
rect 11830 686 11914 714
rect 11606 631 11607 657
rect 11633 631 11634 657
rect 11606 625 11634 631
rect 11382 490 11410 495
rect 11382 443 11410 462
rect 11326 345 11354 350
rect 11886 56 11914 686
rect 12110 686 12194 714
rect 12558 854 12642 882
rect 12110 434 12138 686
rect 12166 602 12194 607
rect 12166 555 12194 574
rect 12446 489 12474 495
rect 12446 463 12447 489
rect 12473 463 12474 489
rect 12110 401 12138 406
rect 12232 406 12364 411
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12232 373 12364 378
rect 12446 266 12474 463
rect 12446 233 12474 238
rect 12558 56 12586 854
rect 12950 546 12978 551
rect 12950 499 12978 518
rect 13230 56 13258 1666
rect 13342 1329 13370 1335
rect 13342 1303 13343 1329
rect 13369 1303 13370 1329
rect 13342 1050 13370 1303
rect 13342 1017 13370 1022
rect 13734 1329 13762 1335
rect 13734 1303 13735 1329
rect 13761 1303 13762 1329
rect 13622 881 13650 887
rect 13622 855 13623 881
rect 13649 855 13650 881
rect 13622 714 13650 855
rect 13622 681 13650 686
rect 13342 545 13370 551
rect 13342 519 13343 545
rect 13369 519 13370 545
rect 13342 490 13370 519
rect 13342 457 13370 462
rect 13734 98 13762 1303
rect 13846 602 13874 1694
rect 13958 1722 13986 4439
rect 14014 4129 14042 4135
rect 14014 4103 14015 4129
rect 14041 4103 14042 4129
rect 14014 2842 14042 4103
rect 14014 2809 14042 2814
rect 13958 1689 13986 1694
rect 14014 2226 14042 2231
rect 13902 1386 13930 1391
rect 13902 1049 13930 1358
rect 14014 1386 14042 2198
rect 14182 1834 14210 6454
rect 14574 6481 14658 6482
rect 14574 6455 14631 6481
rect 14657 6455 14658 6481
rect 14574 6454 14658 6455
rect 14518 6202 14546 6207
rect 14518 6155 14546 6174
rect 14350 6089 14378 6095
rect 14350 6063 14351 6089
rect 14377 6063 14378 6089
rect 14238 5306 14266 5311
rect 14238 5259 14266 5278
rect 14294 5194 14322 5199
rect 14294 4969 14322 5166
rect 14294 4943 14295 4969
rect 14321 4943 14322 4969
rect 14294 4937 14322 4943
rect 14294 4522 14322 4527
rect 14294 4475 14322 4494
rect 14182 1801 14210 1806
rect 14238 4409 14266 4415
rect 14238 4383 14239 4409
rect 14265 4383 14266 4409
rect 14014 1353 14042 1358
rect 13902 1023 13903 1049
rect 13929 1023 13930 1049
rect 13902 1017 13930 1023
rect 13902 602 13930 607
rect 13846 601 13930 602
rect 13846 575 13903 601
rect 13929 575 13930 601
rect 13846 574 13930 575
rect 13902 569 13930 574
rect 13734 65 13762 70
rect 13902 98 13930 103
rect 13902 56 13930 70
rect 14070 98 14098 103
rect 9758 9 9786 14
rect 9856 0 9912 56
rect 10528 0 10584 56
rect 11200 0 11256 56
rect 11872 0 11928 56
rect 12544 0 12600 56
rect 13216 0 13272 56
rect 13888 0 13944 56
rect 14070 42 14098 70
rect 14238 42 14266 4383
rect 14350 3514 14378 6063
rect 14406 5418 14434 5423
rect 14406 4073 14434 5390
rect 14518 5249 14546 5255
rect 14518 5223 14519 5249
rect 14545 5223 14546 5249
rect 14518 4858 14546 5223
rect 14518 4825 14546 4830
rect 14518 4578 14546 4583
rect 14574 4578 14602 6454
rect 14630 6449 14658 6454
rect 15302 6033 15330 6039
rect 15302 6007 15303 6033
rect 15329 6007 15330 6033
rect 15022 5978 15050 5983
rect 15022 5931 15050 5950
rect 15302 5922 15330 6007
rect 15302 5889 15330 5894
rect 14686 5697 14714 5703
rect 14686 5671 14687 5697
rect 14713 5671 14714 5697
rect 14686 5362 14714 5671
rect 14686 5329 14714 5334
rect 15190 5585 15218 5591
rect 15190 5559 15191 5585
rect 15217 5559 15218 5585
rect 14742 5305 14770 5311
rect 14742 5279 14743 5305
rect 14769 5279 14770 5305
rect 14686 4970 14714 4975
rect 14686 4923 14714 4942
rect 14518 4577 14602 4578
rect 14518 4551 14519 4577
rect 14545 4551 14602 4577
rect 14518 4550 14602 4551
rect 14518 4545 14546 4550
rect 14686 4466 14714 4471
rect 14686 4419 14714 4438
rect 14742 4242 14770 5279
rect 15078 5249 15106 5255
rect 15078 5223 15079 5249
rect 15105 5223 15106 5249
rect 15078 4746 15106 5223
rect 15190 4970 15218 5559
rect 15190 4937 15218 4942
rect 15078 4713 15106 4718
rect 15190 4801 15218 4807
rect 15190 4775 15191 4801
rect 15217 4775 15218 4801
rect 15190 4522 15218 4775
rect 15190 4489 15218 4494
rect 15078 4465 15106 4471
rect 15078 4439 15079 4465
rect 15105 4439 15106 4465
rect 15078 4298 15106 4439
rect 15078 4265 15106 4270
rect 14742 4209 14770 4214
rect 14686 4130 14714 4135
rect 14686 4083 14714 4102
rect 14406 4047 14407 4073
rect 14433 4047 14434 4073
rect 14406 4041 14434 4047
rect 14630 4074 14658 4079
rect 14350 3481 14378 3486
rect 14630 3402 14658 4046
rect 15134 4074 15162 4079
rect 14686 3850 14714 3855
rect 14686 3737 14714 3822
rect 15134 3793 15162 4046
rect 15190 4017 15218 4023
rect 15190 3991 15191 4017
rect 15217 3991 15218 4017
rect 15190 3850 15218 3991
rect 15190 3817 15218 3822
rect 15134 3767 15135 3793
rect 15161 3767 15162 3793
rect 15134 3761 15162 3767
rect 14686 3711 14687 3737
rect 14713 3711 14714 3737
rect 14686 3705 14714 3711
rect 14742 3626 14770 3631
rect 14686 3402 14714 3407
rect 14630 3401 14714 3402
rect 14630 3375 14687 3401
rect 14713 3375 14714 3401
rect 14630 3374 14714 3375
rect 14686 3369 14714 3374
rect 14406 3233 14434 3239
rect 14406 3207 14407 3233
rect 14433 3207 14434 3233
rect 14406 3178 14434 3207
rect 14406 3145 14434 3150
rect 14742 2953 14770 3598
rect 15190 3626 15218 3631
rect 15134 3402 15162 3407
rect 15134 3009 15162 3374
rect 15190 3289 15218 3598
rect 15190 3263 15191 3289
rect 15217 3263 15218 3289
rect 15190 3257 15218 3263
rect 15134 2983 15135 3009
rect 15161 2983 15162 3009
rect 15134 2977 15162 2983
rect 14742 2927 14743 2953
rect 14769 2927 14770 2953
rect 14742 2921 14770 2927
rect 15078 2954 15106 2959
rect 14742 2618 14770 2623
rect 14686 2562 14714 2567
rect 14686 2515 14714 2534
rect 14406 2506 14434 2511
rect 14406 2459 14434 2478
rect 14686 2170 14714 2175
rect 14686 2123 14714 2142
rect 14574 2057 14602 2063
rect 14574 2031 14575 2057
rect 14601 2031 14602 2057
rect 14294 1834 14322 1839
rect 14294 1787 14322 1806
rect 14294 1722 14322 1727
rect 14294 1441 14322 1694
rect 14294 1415 14295 1441
rect 14321 1415 14322 1441
rect 14294 1409 14322 1415
rect 14518 1274 14546 1279
rect 14574 1274 14602 2031
rect 14742 1777 14770 2590
rect 15078 2617 15106 2926
rect 15078 2591 15079 2617
rect 15105 2591 15106 2617
rect 15078 2585 15106 2591
rect 15134 2730 15162 2735
rect 15134 2225 15162 2702
rect 15134 2199 15135 2225
rect 15161 2199 15162 2225
rect 15134 2193 15162 2199
rect 15190 2282 15218 2287
rect 14742 1751 14743 1777
rect 14769 1751 14770 1777
rect 14742 1745 14770 1751
rect 15134 2058 15162 2063
rect 14742 1666 14770 1671
rect 14686 1386 14714 1391
rect 14686 1339 14714 1358
rect 14518 1273 14602 1274
rect 14518 1247 14519 1273
rect 14545 1247 14602 1273
rect 14518 1246 14602 1247
rect 14518 1241 14546 1246
rect 14406 1162 14434 1167
rect 14350 938 14378 943
rect 14350 657 14378 910
rect 14406 937 14434 1134
rect 14406 911 14407 937
rect 14433 911 14434 937
rect 14406 905 14434 911
rect 14350 631 14351 657
rect 14377 631 14378 657
rect 14350 625 14378 631
rect 14574 56 14602 1246
rect 14686 1106 14714 1111
rect 14686 601 14714 1078
rect 14742 993 14770 1638
rect 15078 1610 15106 1615
rect 15078 1049 15106 1582
rect 15134 1441 15162 2030
rect 15190 1721 15218 2254
rect 15190 1695 15191 1721
rect 15217 1695 15218 1721
rect 15190 1689 15218 1695
rect 15134 1415 15135 1441
rect 15161 1415 15162 1441
rect 15134 1409 15162 1415
rect 15078 1023 15079 1049
rect 15105 1023 15106 1049
rect 15078 1017 15106 1023
rect 15190 1386 15218 1391
rect 14742 967 14743 993
rect 14769 967 14770 993
rect 14742 961 14770 967
rect 15190 713 15218 1358
rect 15190 687 15191 713
rect 15217 687 15218 713
rect 15190 681 15218 687
rect 14686 575 14687 601
rect 14713 575 14714 601
rect 14686 569 14714 575
rect 14070 14 14266 42
rect 14560 0 14616 56
<< via2 >>
rect 126 6958 154 6986
rect 70 6062 98 6090
rect 2086 6902 2114 6930
rect 1862 6846 1890 6874
rect 1078 6593 1106 6594
rect 1078 6567 1079 6593
rect 1079 6567 1105 6593
rect 1105 6567 1106 6593
rect 1078 6566 1106 6567
rect 1246 6286 1274 6314
rect 1078 5838 1106 5866
rect 686 5614 714 5642
rect 406 5166 434 5194
rect 406 4886 434 4914
rect 910 4718 938 4746
rect 910 4382 938 4410
rect 686 3430 714 3458
rect 126 3038 154 3066
rect 126 2422 154 2450
rect 1902 6285 1930 6286
rect 1902 6259 1903 6285
rect 1903 6259 1929 6285
rect 1929 6259 1930 6285
rect 1902 6258 1930 6259
rect 1954 6285 1982 6286
rect 1954 6259 1955 6285
rect 1955 6259 1981 6285
rect 1981 6259 1982 6285
rect 1954 6258 1982 6259
rect 2006 6285 2034 6286
rect 2006 6259 2007 6285
rect 2007 6259 2033 6285
rect 2033 6259 2034 6285
rect 2006 6258 2034 6259
rect 1918 6201 1946 6202
rect 1918 6175 1919 6201
rect 1919 6175 1945 6201
rect 1945 6175 1946 6201
rect 1918 6174 1946 6175
rect 1806 5782 1834 5810
rect 1358 5166 1386 5194
rect 1806 5614 1834 5642
rect 1902 5501 1930 5502
rect 1902 5475 1903 5501
rect 1903 5475 1929 5501
rect 1929 5475 1930 5501
rect 1902 5474 1930 5475
rect 1954 5501 1982 5502
rect 1954 5475 1955 5501
rect 1955 5475 1981 5501
rect 1981 5475 1982 5501
rect 1954 5474 1982 5475
rect 2006 5501 2034 5502
rect 2006 5475 2007 5501
rect 2007 5475 2033 5501
rect 2033 5475 2034 5501
rect 2006 5474 2034 5475
rect 2232 6677 2260 6678
rect 2232 6651 2233 6677
rect 2233 6651 2259 6677
rect 2259 6651 2260 6677
rect 2232 6650 2260 6651
rect 2284 6677 2312 6678
rect 2284 6651 2285 6677
rect 2285 6651 2311 6677
rect 2311 6651 2312 6677
rect 2284 6650 2312 6651
rect 2336 6677 2364 6678
rect 2336 6651 2337 6677
rect 2337 6651 2363 6677
rect 2363 6651 2364 6677
rect 2336 6650 2364 6651
rect 2198 6033 2226 6034
rect 2198 6007 2199 6033
rect 2199 6007 2225 6033
rect 2225 6007 2226 6033
rect 2198 6006 2226 6007
rect 2232 5893 2260 5894
rect 2232 5867 2233 5893
rect 2233 5867 2259 5893
rect 2259 5867 2260 5893
rect 2232 5866 2260 5867
rect 2284 5893 2312 5894
rect 2284 5867 2285 5893
rect 2285 5867 2311 5893
rect 2311 5867 2312 5893
rect 2284 5866 2312 5867
rect 2336 5893 2364 5894
rect 2336 5867 2337 5893
rect 2337 5867 2363 5893
rect 2363 5867 2364 5893
rect 2336 5866 2364 5867
rect 2310 5726 2338 5754
rect 2422 5670 2450 5698
rect 2232 5109 2260 5110
rect 2232 5083 2233 5109
rect 2233 5083 2259 5109
rect 2259 5083 2260 5109
rect 2232 5082 2260 5083
rect 2284 5109 2312 5110
rect 2284 5083 2285 5109
rect 2285 5083 2311 5109
rect 2311 5083 2312 5109
rect 2284 5082 2312 5083
rect 2336 5109 2364 5110
rect 2336 5083 2337 5109
rect 2337 5083 2363 5109
rect 2363 5083 2364 5109
rect 2336 5082 2364 5083
rect 2142 4998 2170 5026
rect 1902 4717 1930 4718
rect 1902 4691 1903 4717
rect 1903 4691 1929 4717
rect 1929 4691 1930 4717
rect 1902 4690 1930 4691
rect 1954 4717 1982 4718
rect 1954 4691 1955 4717
rect 1955 4691 1981 4717
rect 1981 4691 1982 4717
rect 1954 4690 1982 4691
rect 2006 4717 2034 4718
rect 2006 4691 2007 4717
rect 2007 4691 2033 4717
rect 2033 4691 2034 4717
rect 2006 4690 2034 4691
rect 1862 4465 1890 4466
rect 1862 4439 1863 4465
rect 1863 4439 1889 4465
rect 1889 4439 1890 4465
rect 1862 4438 1890 4439
rect 2232 4325 2260 4326
rect 2232 4299 2233 4325
rect 2233 4299 2259 4325
rect 2259 4299 2260 4325
rect 2232 4298 2260 4299
rect 2284 4325 2312 4326
rect 2284 4299 2285 4325
rect 2285 4299 2311 4325
rect 2311 4299 2312 4325
rect 2284 4298 2312 4299
rect 2336 4325 2364 4326
rect 2336 4299 2337 4325
rect 2337 4299 2363 4325
rect 2363 4299 2364 4325
rect 2336 4298 2364 4299
rect 1582 4102 1610 4130
rect 1902 3933 1930 3934
rect 1902 3907 1903 3933
rect 1903 3907 1929 3933
rect 1929 3907 1930 3933
rect 1902 3906 1930 3907
rect 1954 3933 1982 3934
rect 1954 3907 1955 3933
rect 1955 3907 1981 3933
rect 1981 3907 1982 3933
rect 1954 3906 1982 3907
rect 2006 3933 2034 3934
rect 2006 3907 2007 3933
rect 2007 3907 2033 3933
rect 2033 3907 2034 3933
rect 2006 3906 2034 3907
rect 2590 6145 2618 6146
rect 2590 6119 2591 6145
rect 2591 6119 2617 6145
rect 2617 6119 2618 6145
rect 2590 6118 2618 6119
rect 2758 6118 2786 6146
rect 2702 5614 2730 5642
rect 2590 5361 2618 5362
rect 2590 5335 2591 5361
rect 2591 5335 2617 5361
rect 2617 5335 2618 5361
rect 2590 5334 2618 5335
rect 2758 5334 2786 5362
rect 2534 4830 2562 4858
rect 2646 4886 2674 4914
rect 2590 4465 2618 4466
rect 2590 4439 2591 4465
rect 2591 4439 2617 4465
rect 2617 4439 2618 4465
rect 2590 4438 2618 4439
rect 2590 3934 2618 3962
rect 2478 3878 2506 3906
rect 2534 3822 2562 3850
rect 2232 3541 2260 3542
rect 2232 3515 2233 3541
rect 2233 3515 2259 3541
rect 2259 3515 2260 3541
rect 2232 3514 2260 3515
rect 2284 3541 2312 3542
rect 2284 3515 2285 3541
rect 2285 3515 2311 3541
rect 2311 3515 2312 3541
rect 2284 3514 2312 3515
rect 2336 3541 2364 3542
rect 2336 3515 2337 3541
rect 2337 3515 2363 3541
rect 2363 3515 2364 3541
rect 2336 3514 2364 3515
rect 1902 3149 1930 3150
rect 1902 3123 1903 3149
rect 1903 3123 1929 3149
rect 1929 3123 1930 3149
rect 1902 3122 1930 3123
rect 1954 3149 1982 3150
rect 1954 3123 1955 3149
rect 1955 3123 1981 3149
rect 1981 3123 1982 3149
rect 1954 3122 1982 3123
rect 2006 3149 2034 3150
rect 2006 3123 2007 3149
rect 2007 3123 2033 3149
rect 2033 3123 2034 3149
rect 2006 3122 2034 3123
rect 2232 2757 2260 2758
rect 2232 2731 2233 2757
rect 2233 2731 2259 2757
rect 2259 2731 2260 2757
rect 2232 2730 2260 2731
rect 2284 2757 2312 2758
rect 2284 2731 2285 2757
rect 2285 2731 2311 2757
rect 2311 2731 2312 2757
rect 2284 2730 2312 2731
rect 2336 2757 2364 2758
rect 2336 2731 2337 2757
rect 2337 2731 2363 2757
rect 2363 2731 2364 2757
rect 2336 2730 2364 2731
rect 1414 2478 1442 2506
rect 2982 6622 3010 6650
rect 3150 6566 3178 6594
rect 2870 5670 2898 5698
rect 2982 5894 3010 5922
rect 3094 5838 3122 5866
rect 3262 6566 3290 6594
rect 3374 6174 3402 6202
rect 3206 5726 3234 5754
rect 3094 5502 3122 5530
rect 3486 5502 3514 5530
rect 3486 5417 3514 5418
rect 3486 5391 3487 5417
rect 3487 5391 3513 5417
rect 3513 5391 3514 5417
rect 3486 5390 3514 5391
rect 3318 4913 3346 4914
rect 3318 4887 3319 4913
rect 3319 4887 3345 4913
rect 3345 4887 3346 4913
rect 3318 4886 3346 4887
rect 3654 6230 3682 6258
rect 3598 4774 3626 4802
rect 3822 6846 3850 6874
rect 3766 6790 3794 6818
rect 3766 6062 3794 6090
rect 3878 5838 3906 5866
rect 3878 5641 3906 5642
rect 3878 5615 3879 5641
rect 3879 5615 3905 5641
rect 3905 5615 3906 5641
rect 3878 5614 3906 5615
rect 4046 5390 4074 5418
rect 4158 6678 4186 6706
rect 4214 6174 4242 6202
rect 4158 5697 4186 5698
rect 4158 5671 4159 5697
rect 4159 5671 4185 5697
rect 4185 5671 4186 5697
rect 4158 5670 4186 5671
rect 4158 5446 4186 5474
rect 4382 6622 4410 6650
rect 3262 4270 3290 4298
rect 3878 4774 3906 4802
rect 2758 3934 2786 3962
rect 3486 4102 3514 4130
rect 2646 2814 2674 2842
rect 3374 3430 3402 3458
rect 2534 2478 2562 2506
rect 1902 2365 1930 2366
rect 1902 2339 1903 2365
rect 1903 2339 1929 2365
rect 1929 2339 1930 2365
rect 1902 2338 1930 2339
rect 1954 2365 1982 2366
rect 1954 2339 1955 2365
rect 1955 2339 1981 2365
rect 1981 2339 1982 2365
rect 1954 2338 1982 2339
rect 2006 2365 2034 2366
rect 2006 2339 2007 2365
rect 2007 2339 2033 2365
rect 2033 2339 2034 2365
rect 2006 2338 2034 2339
rect 1414 2142 1442 2170
rect 2232 1973 2260 1974
rect 2232 1947 2233 1973
rect 2233 1947 2259 1973
rect 2259 1947 2260 1973
rect 2232 1946 2260 1947
rect 2284 1973 2312 1974
rect 2284 1947 2285 1973
rect 2285 1947 2311 1973
rect 2311 1947 2312 1973
rect 2284 1946 2312 1947
rect 2336 1973 2364 1974
rect 2336 1947 2337 1973
rect 2337 1947 2363 1973
rect 2363 1947 2364 1973
rect 3374 1974 3402 2002
rect 2336 1946 2364 1947
rect 1246 1862 1274 1890
rect 1902 1581 1930 1582
rect 1902 1555 1903 1581
rect 1903 1555 1929 1581
rect 1929 1555 1930 1581
rect 1902 1554 1930 1555
rect 1954 1581 1982 1582
rect 1954 1555 1955 1581
rect 1955 1555 1981 1581
rect 1981 1555 1982 1581
rect 1954 1554 1982 1555
rect 2006 1581 2034 1582
rect 2006 1555 2007 1581
rect 2007 1555 2033 1581
rect 2033 1555 2034 1581
rect 2006 1554 2034 1555
rect 1078 1470 1106 1498
rect 2232 1189 2260 1190
rect 2232 1163 2233 1189
rect 2233 1163 2259 1189
rect 2259 1163 2260 1189
rect 2232 1162 2260 1163
rect 2284 1189 2312 1190
rect 2284 1163 2285 1189
rect 2285 1163 2311 1189
rect 2311 1163 2312 1189
rect 2284 1162 2312 1163
rect 2336 1189 2364 1190
rect 2336 1163 2337 1189
rect 2337 1163 2363 1189
rect 2363 1163 2364 1189
rect 2336 1162 2364 1163
rect 3150 966 3178 994
rect 1806 854 1834 882
rect 1134 70 1162 98
rect 1902 797 1930 798
rect 1902 771 1903 797
rect 1903 771 1929 797
rect 1929 771 1930 797
rect 1902 770 1930 771
rect 1954 797 1982 798
rect 1954 771 1955 797
rect 1955 771 1981 797
rect 1981 771 1982 797
rect 1954 770 1982 771
rect 2006 797 2034 798
rect 2006 771 2007 797
rect 2007 771 2033 797
rect 2033 771 2034 797
rect 2006 770 2034 771
rect 2232 405 2260 406
rect 2232 379 2233 405
rect 2233 379 2259 405
rect 2259 379 2260 405
rect 2232 378 2260 379
rect 2284 405 2312 406
rect 2284 379 2285 405
rect 2285 379 2311 405
rect 2311 379 2312 405
rect 2284 378 2312 379
rect 2336 405 2364 406
rect 2336 379 2337 405
rect 2337 379 2363 405
rect 2363 379 2364 405
rect 2336 378 2364 379
rect 2478 70 2506 98
rect 3486 798 3514 826
rect 4102 4718 4130 4746
rect 3990 4046 4018 4074
rect 4718 6230 4746 6258
rect 4774 6958 4802 6986
rect 4606 6174 4634 6202
rect 4494 6006 4522 6034
rect 4550 5894 4578 5922
rect 4438 5614 4466 5642
rect 4662 5838 4690 5866
rect 4438 4998 4466 5026
rect 4158 4438 4186 4466
rect 4886 6846 4914 6874
rect 4830 5278 4858 5306
rect 4998 6958 5026 6986
rect 5054 6790 5082 6818
rect 5166 6678 5194 6706
rect 5166 6286 5194 6314
rect 5054 6201 5082 6202
rect 5054 6175 5055 6201
rect 5055 6175 5081 6201
rect 5081 6175 5082 6201
rect 5054 6174 5082 6175
rect 5166 6118 5194 6146
rect 5334 6033 5362 6034
rect 5334 6007 5335 6033
rect 5335 6007 5361 6033
rect 5361 6007 5362 6033
rect 5334 6006 5362 6007
rect 5670 6622 5698 6650
rect 5614 6174 5642 6202
rect 5502 6118 5530 6146
rect 5502 5950 5530 5978
rect 5838 6846 5866 6874
rect 5950 6678 5978 6706
rect 5950 6230 5978 6258
rect 6006 6201 6034 6202
rect 6006 6175 6007 6201
rect 6007 6175 6033 6201
rect 6033 6175 6034 6201
rect 6006 6174 6034 6175
rect 5334 5334 5362 5362
rect 5222 5278 5250 5306
rect 4774 4606 4802 4634
rect 5334 4550 5362 4578
rect 3822 3737 3850 3738
rect 3822 3711 3823 3737
rect 3823 3711 3849 3737
rect 3849 3711 3850 3737
rect 3822 3710 3850 3711
rect 4326 3681 4354 3682
rect 4326 3655 4327 3681
rect 4327 3655 4353 3681
rect 4353 3655 4354 3681
rect 4326 3654 4354 3655
rect 4438 3681 4466 3682
rect 4438 3655 4439 3681
rect 4439 3655 4465 3681
rect 4465 3655 4466 3681
rect 4438 3654 4466 3655
rect 3878 3430 3906 3458
rect 5278 4326 5306 4354
rect 5502 4270 5530 4298
rect 5054 4073 5082 4074
rect 5054 4047 5055 4073
rect 5055 4047 5081 4073
rect 5081 4047 5082 4073
rect 5054 4046 5082 4047
rect 5670 5614 5698 5642
rect 5558 3990 5586 4018
rect 5614 4326 5642 4354
rect 5166 3878 5194 3906
rect 5838 5838 5866 5866
rect 5726 4718 5754 4746
rect 5726 4465 5754 4466
rect 5726 4439 5727 4465
rect 5727 4439 5753 4465
rect 5753 4439 5754 4465
rect 5726 4438 5754 4439
rect 6286 6622 6314 6650
rect 6342 6678 6370 6706
rect 6174 6174 6202 6202
rect 6286 5670 6314 5698
rect 6510 6118 6538 6146
rect 6566 6790 6594 6818
rect 6734 6902 6762 6930
rect 6622 6566 6650 6594
rect 6678 6398 6706 6426
rect 6454 5278 6482 5306
rect 6118 5249 6146 5250
rect 6118 5223 6119 5249
rect 6119 5223 6145 5249
rect 6145 5223 6146 5249
rect 6118 5222 6146 5223
rect 6174 5110 6202 5138
rect 5838 4270 5866 4298
rect 5950 4886 5978 4914
rect 6118 4913 6146 4914
rect 6118 4887 6119 4913
rect 6119 4887 6145 4913
rect 6145 4887 6146 4913
rect 6118 4886 6146 4887
rect 6790 6145 6818 6146
rect 6790 6119 6791 6145
rect 6791 6119 6817 6145
rect 6817 6119 6818 6145
rect 6790 6118 6818 6119
rect 6734 5278 6762 5306
rect 6790 5726 6818 5754
rect 6678 4662 6706 4690
rect 6790 4326 6818 4354
rect 6230 4185 6258 4186
rect 6230 4159 6231 4185
rect 6231 4159 6257 4185
rect 6257 4159 6258 4185
rect 6230 4158 6258 4159
rect 6398 4185 6426 4186
rect 6398 4159 6399 4185
rect 6399 4159 6425 4185
rect 6425 4159 6426 4185
rect 6398 4158 6426 4159
rect 5782 4129 5810 4130
rect 5782 4103 5783 4129
rect 5783 4103 5809 4129
rect 5809 4103 5810 4129
rect 5782 4102 5810 4103
rect 5950 4046 5978 4074
rect 7070 6958 7098 6986
rect 7014 6593 7042 6594
rect 7014 6567 7015 6593
rect 7015 6567 7041 6593
rect 7041 6567 7042 6593
rect 7014 6566 7042 6567
rect 7126 6342 7154 6370
rect 7014 6118 7042 6146
rect 6902 4857 6930 4858
rect 6902 4831 6903 4857
rect 6903 4831 6929 4857
rect 6929 4831 6930 4857
rect 6902 4830 6930 4831
rect 6902 4662 6930 4690
rect 6846 3934 6874 3962
rect 6902 3878 6930 3906
rect 4942 3430 4970 3458
rect 4158 3206 4186 3234
rect 4438 3345 4466 3346
rect 4438 3319 4439 3345
rect 4439 3319 4465 3345
rect 4465 3319 4466 3345
rect 4438 3318 4466 3319
rect 4438 3206 4466 3234
rect 6622 2030 6650 2058
rect 7238 6174 7266 6202
rect 7294 5614 7322 5642
rect 7350 6678 7378 6706
rect 7070 4102 7098 4130
rect 7126 5446 7154 5474
rect 6958 3710 6986 3738
rect 7182 5166 7210 5194
rect 7406 5894 7434 5922
rect 7462 5726 7490 5754
rect 7462 5446 7490 5474
rect 7406 5390 7434 5418
rect 7574 6537 7602 6538
rect 7574 6511 7575 6537
rect 7575 6511 7601 6537
rect 7601 6511 7602 6537
rect 7574 6510 7602 6511
rect 7742 7014 7770 7042
rect 7854 6678 7882 6706
rect 7854 6593 7882 6594
rect 7854 6567 7855 6593
rect 7855 6567 7881 6593
rect 7881 6567 7882 6593
rect 7854 6566 7882 6567
rect 7686 5894 7714 5922
rect 7518 5110 7546 5138
rect 7462 4857 7490 4858
rect 7462 4831 7463 4857
rect 7463 4831 7489 4857
rect 7489 4831 7490 4857
rect 7462 4830 7490 4831
rect 7630 5446 7658 5474
rect 7686 5390 7714 5418
rect 7686 4830 7714 4858
rect 7462 4494 7490 4522
rect 7406 4409 7434 4410
rect 7406 4383 7407 4409
rect 7407 4383 7433 4409
rect 7433 4383 7434 4409
rect 7406 4382 7434 4383
rect 7574 4409 7602 4410
rect 7574 4383 7575 4409
rect 7575 4383 7601 4409
rect 7601 4383 7602 4409
rect 7574 4382 7602 4383
rect 7910 5641 7938 5642
rect 7910 5615 7911 5641
rect 7911 5615 7937 5641
rect 7937 5615 7938 5641
rect 7910 5614 7938 5615
rect 7966 5390 7994 5418
rect 7966 4942 7994 4970
rect 7854 4606 7882 4634
rect 7966 4857 7994 4858
rect 7966 4831 7967 4857
rect 7967 4831 7993 4857
rect 7993 4831 7994 4857
rect 7966 4830 7994 4831
rect 7966 4270 7994 4298
rect 7854 4214 7882 4242
rect 7630 4158 7658 4186
rect 7126 3542 7154 3570
rect 7686 3766 7714 3794
rect 7630 3598 7658 3626
rect 7574 3486 7602 3514
rect 7798 3766 7826 3794
rect 7238 3374 7266 3402
rect 7014 3289 7042 3290
rect 7014 3263 7015 3289
rect 7015 3263 7041 3289
rect 7041 3263 7042 3289
rect 7014 3262 7042 3263
rect 8246 6902 8274 6930
rect 8134 6593 8162 6594
rect 8134 6567 8135 6593
rect 8135 6567 8161 6593
rect 8161 6567 8162 6593
rect 8134 6566 8162 6567
rect 8078 6454 8106 6482
rect 8414 6790 8442 6818
rect 8638 6902 8666 6930
rect 8526 6566 8554 6594
rect 8694 6678 8722 6706
rect 8862 6510 8890 6538
rect 8806 6286 8834 6314
rect 8078 5894 8106 5922
rect 8750 6089 8778 6090
rect 8750 6063 8751 6089
rect 8751 6063 8777 6089
rect 8777 6063 8778 6089
rect 8750 6062 8778 6063
rect 8302 5502 8330 5530
rect 8134 4830 8162 4858
rect 8302 4774 8330 4802
rect 8078 4073 8106 4074
rect 8078 4047 8079 4073
rect 8079 4047 8105 4073
rect 8105 4047 8106 4073
rect 8078 4046 8106 4047
rect 8078 3793 8106 3794
rect 8078 3767 8079 3793
rect 8079 3767 8105 3793
rect 8105 3767 8106 3793
rect 8078 3766 8106 3767
rect 7966 3318 7994 3346
rect 8078 3318 8106 3346
rect 7182 3262 7210 3290
rect 7462 3289 7490 3290
rect 7462 3263 7463 3289
rect 7463 3263 7489 3289
rect 7489 3263 7490 3289
rect 7462 3262 7490 3263
rect 7518 3009 7546 3010
rect 7518 2983 7519 3009
rect 7519 2983 7545 3009
rect 7545 2983 7546 3009
rect 7518 2982 7546 2983
rect 7182 2926 7210 2954
rect 7070 2841 7098 2842
rect 7070 2815 7071 2841
rect 7071 2815 7097 2841
rect 7097 2815 7098 2841
rect 7070 2814 7098 2815
rect 7462 2926 7490 2954
rect 7238 2841 7266 2842
rect 7238 2815 7239 2841
rect 7239 2815 7265 2841
rect 7265 2815 7266 2841
rect 7238 2814 7266 2815
rect 7070 2198 7098 2226
rect 7014 2057 7042 2058
rect 7014 2031 7015 2057
rect 7015 2031 7041 2057
rect 7041 2031 7042 2057
rect 7014 2030 7042 2031
rect 7294 2057 7322 2058
rect 7294 2031 7295 2057
rect 7295 2031 7321 2057
rect 7321 2031 7322 2057
rect 7294 2030 7322 2031
rect 7014 1806 7042 1834
rect 7238 1721 7266 1722
rect 7238 1695 7239 1721
rect 7239 1695 7265 1721
rect 7265 1695 7266 1721
rect 7238 1694 7266 1695
rect 6846 1638 6874 1666
rect 7294 1638 7322 1666
rect 6790 1022 6818 1050
rect 7406 1049 7434 1050
rect 7406 1023 7407 1049
rect 7407 1023 7433 1049
rect 7433 1023 7434 1049
rect 7406 1022 7434 1023
rect 3598 406 3626 434
rect 3822 854 3850 882
rect 5166 798 5194 826
rect 4494 294 4522 322
rect 6958 798 6986 826
rect 6342 742 6370 770
rect 5558 657 5586 658
rect 5558 631 5559 657
rect 5559 631 5585 657
rect 5585 631 5586 657
rect 5558 630 5586 631
rect 7126 798 7154 826
rect 8022 2646 8050 2674
rect 8134 2926 8162 2954
rect 8078 2617 8106 2618
rect 8078 2591 8079 2617
rect 8079 2591 8105 2617
rect 8105 2591 8106 2617
rect 8078 2590 8106 2591
rect 7518 2561 7546 2562
rect 7518 2535 7519 2561
rect 7519 2535 7545 2561
rect 7545 2535 7546 2561
rect 7518 2534 7546 2535
rect 7630 2254 7658 2282
rect 8190 2478 8218 2506
rect 8246 3710 8274 3738
rect 7518 2086 7546 2114
rect 7686 1974 7714 2002
rect 7518 1385 7546 1386
rect 7518 1359 7519 1385
rect 7519 1359 7545 1385
rect 7545 1359 7546 1385
rect 7518 1358 7546 1359
rect 7686 1385 7714 1386
rect 7686 1359 7687 1385
rect 7687 1359 7713 1385
rect 7713 1359 7714 1385
rect 7686 1358 7714 1359
rect 8022 1246 8050 1274
rect 8078 1414 8106 1442
rect 7966 1078 7994 1106
rect 8134 1273 8162 1274
rect 8134 1247 8135 1273
rect 8135 1247 8161 1273
rect 8161 1247 8162 1273
rect 8134 1246 8162 1247
rect 9198 6678 9226 6706
rect 9310 6454 9338 6482
rect 8974 6398 9002 6426
rect 9478 6622 9506 6650
rect 8862 6174 8890 6202
rect 9198 6286 9226 6314
rect 8974 6089 9002 6090
rect 8974 6063 8975 6089
rect 8975 6063 9001 6089
rect 9001 6063 9002 6089
rect 8974 6062 9002 6063
rect 9142 6062 9170 6090
rect 9254 6145 9282 6146
rect 9254 6119 9255 6145
rect 9255 6119 9281 6145
rect 9281 6119 9282 6145
rect 9254 6118 9282 6119
rect 9086 5726 9114 5754
rect 9030 5614 9058 5642
rect 8358 4438 8386 4466
rect 8414 5110 8442 5138
rect 8470 4102 8498 4130
rect 9534 6286 9562 6314
rect 9702 6342 9730 6370
rect 9366 5950 9394 5978
rect 9534 5894 9562 5922
rect 9758 5894 9786 5922
rect 9814 5726 9842 5754
rect 9310 5558 9338 5586
rect 9366 5502 9394 5530
rect 9254 5249 9282 5250
rect 9254 5223 9255 5249
rect 9255 5223 9281 5249
rect 9281 5223 9282 5249
rect 9254 5222 9282 5223
rect 9030 3878 9058 3906
rect 9310 3822 9338 3850
rect 8414 3766 8442 3794
rect 8918 3654 8946 3682
rect 8358 3345 8386 3346
rect 8358 3319 8359 3345
rect 8359 3319 8385 3345
rect 8385 3319 8386 3345
rect 8358 3318 8386 3319
rect 8302 2982 8330 3010
rect 8302 2169 8330 2170
rect 8302 2143 8303 2169
rect 8303 2143 8329 2169
rect 8329 2143 8330 2169
rect 8302 2142 8330 2143
rect 8750 2702 8778 2730
rect 8694 2646 8722 2674
rect 8862 2702 8890 2730
rect 8638 2142 8666 2170
rect 8638 1470 8666 1498
rect 9198 3430 9226 3458
rect 9142 2814 9170 2842
rect 8358 1358 8386 1386
rect 9142 937 9170 938
rect 9142 911 9143 937
rect 9143 911 9169 937
rect 9169 911 9170 937
rect 9142 910 9170 911
rect 8246 742 8274 770
rect 7630 686 7658 714
rect 6958 126 6986 154
rect 7462 630 7490 658
rect 8134 630 8162 658
rect 7854 601 7882 602
rect 7854 575 7855 601
rect 7855 575 7881 601
rect 7881 575 7882 601
rect 7854 574 7882 575
rect 8134 545 8162 546
rect 8134 519 8135 545
rect 8135 519 8161 545
rect 8161 519 8162 545
rect 8134 518 8162 519
rect 8526 657 8554 658
rect 8526 631 8527 657
rect 8527 631 8553 657
rect 8553 631 8554 657
rect 8526 630 8554 631
rect 9310 910 9338 938
rect 8358 518 8386 546
rect 7854 462 7882 490
rect 7462 238 7490 266
rect 8806 489 8834 490
rect 8806 463 8807 489
rect 8807 463 8833 489
rect 8833 463 8834 489
rect 8806 462 8834 463
rect 8918 489 8946 490
rect 8918 463 8919 489
rect 8919 463 8945 489
rect 8945 463 8946 489
rect 8918 462 8946 463
rect 8526 350 8554 378
rect 9926 6006 9954 6034
rect 10038 6230 10066 6258
rect 9982 5390 10010 5418
rect 9926 5054 9954 5082
rect 9478 1862 9506 1890
rect 9590 4270 9618 4298
rect 10150 5950 10178 5978
rect 10262 6734 10290 6762
rect 10262 5950 10290 5978
rect 10430 6734 10458 6762
rect 10542 6398 10570 6426
rect 10486 6062 10514 6090
rect 10542 6006 10570 6034
rect 10430 5838 10458 5866
rect 10094 5558 10122 5586
rect 10150 5390 10178 5418
rect 10430 5670 10458 5698
rect 10486 5641 10514 5642
rect 10486 5615 10487 5641
rect 10487 5615 10513 5641
rect 10513 5615 10514 5641
rect 10486 5614 10514 5615
rect 10374 5278 10402 5306
rect 10038 4606 10066 4634
rect 9926 3934 9954 3962
rect 10038 3822 10066 3850
rect 10206 993 10234 994
rect 10206 967 10207 993
rect 10207 967 10233 993
rect 10233 967 10234 993
rect 10206 966 10234 967
rect 9366 294 9394 322
rect 10430 5558 10458 5586
rect 10990 6622 11018 6650
rect 10878 6566 10906 6594
rect 11102 6510 11130 6538
rect 10766 6006 10794 6034
rect 10710 5950 10738 5978
rect 10766 5894 10794 5922
rect 10654 5614 10682 5642
rect 10654 5305 10682 5306
rect 10654 5279 10655 5305
rect 10655 5279 10681 5305
rect 10681 5279 10682 5305
rect 10654 5278 10682 5279
rect 10878 6342 10906 6370
rect 10878 5894 10906 5922
rect 10822 4998 10850 5026
rect 10654 4382 10682 4410
rect 10654 2422 10682 2450
rect 10878 4886 10906 4914
rect 10990 5278 11018 5306
rect 10934 4270 10962 4298
rect 10766 3990 10794 4018
rect 11102 5894 11130 5922
rect 11158 5838 11186 5866
rect 11270 6593 11298 6594
rect 11270 6567 11271 6593
rect 11271 6567 11297 6593
rect 11297 6567 11298 6593
rect 11270 6566 11298 6567
rect 11326 6174 11354 6202
rect 11382 6622 11410 6650
rect 11214 5782 11242 5810
rect 11158 5305 11186 5306
rect 11158 5279 11159 5305
rect 11159 5279 11185 5305
rect 11185 5279 11186 5305
rect 11158 5278 11186 5279
rect 11046 3822 11074 3850
rect 11102 5222 11130 5250
rect 11158 5166 11186 5194
rect 11102 3430 11130 3458
rect 10878 1806 10906 1834
rect 10710 1273 10738 1274
rect 10710 1247 10711 1273
rect 10711 1247 10737 1273
rect 10737 1247 10738 1273
rect 10710 1246 10738 1247
rect 10598 1134 10626 1162
rect 10374 993 10402 994
rect 10374 967 10375 993
rect 10375 967 10401 993
rect 10401 967 10402 993
rect 10374 966 10402 967
rect 9198 238 9226 266
rect 9646 70 9674 98
rect 9870 294 9898 322
rect 10822 1246 10850 1274
rect 10822 854 10850 882
rect 11550 6902 11578 6930
rect 11662 6454 11690 6482
rect 11606 5809 11634 5810
rect 11606 5783 11607 5809
rect 11607 5783 11633 5809
rect 11633 5783 11634 5809
rect 11606 5782 11634 5783
rect 11550 5726 11578 5754
rect 11438 5390 11466 5418
rect 11494 5670 11522 5698
rect 11326 5361 11354 5362
rect 11326 5335 11327 5361
rect 11327 5335 11353 5361
rect 11353 5335 11354 5361
rect 11326 5334 11354 5335
rect 11998 6566 12026 6594
rect 11774 5614 11802 5642
rect 11942 6342 11970 6370
rect 11902 6285 11930 6286
rect 11902 6259 11903 6285
rect 11903 6259 11929 6285
rect 11929 6259 11930 6285
rect 11902 6258 11930 6259
rect 11954 6285 11982 6286
rect 11954 6259 11955 6285
rect 11955 6259 11981 6285
rect 11981 6259 11982 6285
rect 11954 6258 11982 6259
rect 12006 6285 12034 6286
rect 12006 6259 12007 6285
rect 12007 6259 12033 6285
rect 12033 6259 12034 6285
rect 12006 6258 12034 6259
rect 11998 6201 12026 6202
rect 11998 6175 11999 6201
rect 11999 6175 12025 6201
rect 12025 6175 12026 6201
rect 11998 6174 12026 6175
rect 11830 5558 11858 5586
rect 11902 5501 11930 5502
rect 11902 5475 11903 5501
rect 11903 5475 11929 5501
rect 11929 5475 11930 5501
rect 11902 5474 11930 5475
rect 11954 5501 11982 5502
rect 11954 5475 11955 5501
rect 11955 5475 11981 5501
rect 11981 5475 11982 5501
rect 11954 5474 11982 5475
rect 12006 5501 12034 5502
rect 12006 5475 12007 5501
rect 12007 5475 12033 5501
rect 12033 5475 12034 5501
rect 12006 5474 12034 5475
rect 12334 6846 12362 6874
rect 12222 6790 12250 6818
rect 12232 6677 12260 6678
rect 12232 6651 12233 6677
rect 12233 6651 12259 6677
rect 12259 6651 12260 6677
rect 12232 6650 12260 6651
rect 12284 6677 12312 6678
rect 12284 6651 12285 6677
rect 12285 6651 12311 6677
rect 12311 6651 12312 6677
rect 12284 6650 12312 6651
rect 12336 6677 12364 6678
rect 12336 6651 12337 6677
rect 12337 6651 12363 6677
rect 12363 6651 12364 6677
rect 12336 6650 12364 6651
rect 12222 6510 12250 6538
rect 12110 5446 12138 5474
rect 12166 6398 12194 6426
rect 11830 5417 11858 5418
rect 11830 5391 11831 5417
rect 11831 5391 11857 5417
rect 11857 5391 11858 5417
rect 11830 5390 11858 5391
rect 11774 5278 11802 5306
rect 11774 5054 11802 5082
rect 11718 4998 11746 5026
rect 11382 4830 11410 4858
rect 11606 4886 11634 4914
rect 11326 4409 11354 4410
rect 11326 4383 11327 4409
rect 11327 4383 11353 4409
rect 11353 4383 11354 4409
rect 11326 4382 11354 4383
rect 11550 4382 11578 4410
rect 11214 910 11242 938
rect 10430 294 10458 322
rect 11102 489 11130 490
rect 11102 463 11103 489
rect 11103 463 11129 489
rect 11129 463 11130 489
rect 11102 462 11130 463
rect 11158 350 11186 378
rect 11102 238 11130 266
rect 11662 4830 11690 4858
rect 11942 4857 11970 4858
rect 11942 4831 11943 4857
rect 11943 4831 11969 4857
rect 11969 4831 11970 4857
rect 11942 4830 11970 4831
rect 11902 4717 11930 4718
rect 11902 4691 11903 4717
rect 11903 4691 11929 4717
rect 11929 4691 11930 4717
rect 11902 4690 11930 4691
rect 11954 4717 11982 4718
rect 11954 4691 11955 4717
rect 11955 4691 11981 4717
rect 11981 4691 11982 4717
rect 11954 4690 11982 4691
rect 12006 4717 12034 4718
rect 12006 4691 12007 4717
rect 12007 4691 12033 4717
rect 12033 4691 12034 4717
rect 12006 4690 12034 4691
rect 12232 5893 12260 5894
rect 12232 5867 12233 5893
rect 12233 5867 12259 5893
rect 12259 5867 12260 5893
rect 12232 5866 12260 5867
rect 12284 5893 12312 5894
rect 12284 5867 12285 5893
rect 12285 5867 12311 5893
rect 12311 5867 12312 5893
rect 12284 5866 12312 5867
rect 12336 5893 12364 5894
rect 12336 5867 12337 5893
rect 12337 5867 12363 5893
rect 12363 5867 12364 5893
rect 12336 5866 12364 5867
rect 12558 6342 12586 6370
rect 12726 6398 12754 6426
rect 12670 6174 12698 6202
rect 12726 6286 12754 6314
rect 12502 6033 12530 6034
rect 12502 6007 12503 6033
rect 12503 6007 12529 6033
rect 12529 6007 12530 6033
rect 12502 6006 12530 6007
rect 12670 5838 12698 5866
rect 12558 5641 12586 5642
rect 12558 5615 12559 5641
rect 12559 5615 12585 5641
rect 12585 5615 12586 5641
rect 12558 5614 12586 5615
rect 12614 5558 12642 5586
rect 12278 5278 12306 5306
rect 12558 5446 12586 5474
rect 12334 5249 12362 5250
rect 12334 5223 12335 5249
rect 12335 5223 12361 5249
rect 12361 5223 12362 5249
rect 12334 5222 12362 5223
rect 12232 5109 12260 5110
rect 12232 5083 12233 5109
rect 12233 5083 12259 5109
rect 12259 5083 12260 5109
rect 12232 5082 12260 5083
rect 12284 5109 12312 5110
rect 12284 5083 12285 5109
rect 12285 5083 12311 5109
rect 12311 5083 12312 5109
rect 12284 5082 12312 5083
rect 12336 5109 12364 5110
rect 12336 5083 12337 5109
rect 12337 5083 12363 5109
rect 12363 5083 12364 5109
rect 12336 5082 12364 5083
rect 12614 4998 12642 5026
rect 12278 4913 12306 4914
rect 12278 4887 12279 4913
rect 12279 4887 12305 4913
rect 12305 4887 12306 4913
rect 12278 4886 12306 4887
rect 12446 4606 12474 4634
rect 11830 4326 11858 4354
rect 11902 3933 11930 3934
rect 11902 3907 11903 3933
rect 11903 3907 11929 3933
rect 11929 3907 11930 3933
rect 11902 3906 11930 3907
rect 11954 3933 11982 3934
rect 11954 3907 11955 3933
rect 11955 3907 11981 3933
rect 11981 3907 11982 3933
rect 11954 3906 11982 3907
rect 12006 3933 12034 3934
rect 12006 3907 12007 3933
rect 12007 3907 12033 3933
rect 12033 3907 12034 3933
rect 12006 3906 12034 3907
rect 12110 3766 12138 3794
rect 11902 3149 11930 3150
rect 11902 3123 11903 3149
rect 11903 3123 11929 3149
rect 11929 3123 11930 3149
rect 11902 3122 11930 3123
rect 11954 3149 11982 3150
rect 11954 3123 11955 3149
rect 11955 3123 11981 3149
rect 11981 3123 11982 3149
rect 11954 3122 11982 3123
rect 12006 3149 12034 3150
rect 12006 3123 12007 3149
rect 12007 3123 12033 3149
rect 12033 3123 12034 3149
rect 12006 3122 12034 3123
rect 11902 2365 11930 2366
rect 11902 2339 11903 2365
rect 11903 2339 11929 2365
rect 11929 2339 11930 2365
rect 11902 2338 11930 2339
rect 11954 2365 11982 2366
rect 11954 2339 11955 2365
rect 11955 2339 11981 2365
rect 11981 2339 11982 2365
rect 11954 2338 11982 2339
rect 12006 2365 12034 2366
rect 12006 2339 12007 2365
rect 12007 2339 12033 2365
rect 12033 2339 12034 2365
rect 12006 2338 12034 2339
rect 11902 1581 11930 1582
rect 11902 1555 11903 1581
rect 11903 1555 11929 1581
rect 11929 1555 11930 1581
rect 11902 1554 11930 1555
rect 11954 1581 11982 1582
rect 11954 1555 11955 1581
rect 11955 1555 11981 1581
rect 11981 1555 11982 1581
rect 11954 1554 11982 1555
rect 12006 1581 12034 1582
rect 12006 1555 12007 1581
rect 12007 1555 12033 1581
rect 12033 1555 12034 1581
rect 12006 1554 12034 1555
rect 11662 1134 11690 1162
rect 11902 797 11930 798
rect 11902 771 11903 797
rect 11903 771 11929 797
rect 11929 771 11930 797
rect 11902 770 11930 771
rect 11954 797 11982 798
rect 11954 771 11955 797
rect 11955 771 11981 797
rect 11981 771 11982 797
rect 11954 770 11982 771
rect 12006 797 12034 798
rect 12006 771 12007 797
rect 12007 771 12033 797
rect 12033 771 12034 797
rect 12006 770 12034 771
rect 12232 4325 12260 4326
rect 12232 4299 12233 4325
rect 12233 4299 12259 4325
rect 12259 4299 12260 4325
rect 12232 4298 12260 4299
rect 12284 4325 12312 4326
rect 12284 4299 12285 4325
rect 12285 4299 12311 4325
rect 12311 4299 12312 4325
rect 12284 4298 12312 4299
rect 12336 4325 12364 4326
rect 12336 4299 12337 4325
rect 12337 4299 12363 4325
rect 12363 4299 12364 4325
rect 12336 4298 12364 4299
rect 12614 4382 12642 4410
rect 12782 5950 12810 5978
rect 12838 6958 12866 6986
rect 13006 7014 13034 7042
rect 13398 7014 13426 7042
rect 12894 6734 12922 6762
rect 12950 6902 12978 6930
rect 12950 6454 12978 6482
rect 13006 6398 13034 6426
rect 12894 5838 12922 5866
rect 12894 3710 12922 3738
rect 12232 3541 12260 3542
rect 12232 3515 12233 3541
rect 12233 3515 12259 3541
rect 12259 3515 12260 3541
rect 12232 3514 12260 3515
rect 12284 3541 12312 3542
rect 12284 3515 12285 3541
rect 12285 3515 12311 3541
rect 12311 3515 12312 3541
rect 12284 3514 12312 3515
rect 12336 3541 12364 3542
rect 12336 3515 12337 3541
rect 12337 3515 12363 3541
rect 12363 3515 12364 3541
rect 12336 3514 12364 3515
rect 12950 3486 12978 3514
rect 12232 2757 12260 2758
rect 12232 2731 12233 2757
rect 12233 2731 12259 2757
rect 12259 2731 12260 2757
rect 12232 2730 12260 2731
rect 12284 2757 12312 2758
rect 12284 2731 12285 2757
rect 12285 2731 12311 2757
rect 12311 2731 12312 2757
rect 12284 2730 12312 2731
rect 12336 2757 12364 2758
rect 12336 2731 12337 2757
rect 12337 2731 12363 2757
rect 12363 2731 12364 2757
rect 12336 2730 12364 2731
rect 12232 1973 12260 1974
rect 12232 1947 12233 1973
rect 12233 1947 12259 1973
rect 12259 1947 12260 1973
rect 12232 1946 12260 1947
rect 12284 1973 12312 1974
rect 12284 1947 12285 1973
rect 12285 1947 12311 1973
rect 12311 1947 12312 1973
rect 12284 1946 12312 1947
rect 12336 1973 12364 1974
rect 12336 1947 12337 1973
rect 12337 1947 12363 1973
rect 12363 1947 12364 1973
rect 12336 1946 12364 1947
rect 13174 5950 13202 5978
rect 13118 5894 13146 5922
rect 13062 4998 13090 5026
rect 13006 2870 13034 2898
rect 12232 1189 12260 1190
rect 12232 1163 12233 1189
rect 12233 1163 12259 1189
rect 12259 1163 12260 1189
rect 12232 1162 12260 1163
rect 12284 1189 12312 1190
rect 12284 1163 12285 1189
rect 12285 1163 12311 1189
rect 12311 1163 12312 1189
rect 12284 1162 12312 1163
rect 12336 1189 12364 1190
rect 12336 1163 12337 1189
rect 12337 1163 12363 1189
rect 12363 1163 12364 1189
rect 12336 1162 12364 1163
rect 12558 993 12586 994
rect 12558 967 12559 993
rect 12559 967 12585 993
rect 12585 967 12586 993
rect 12558 966 12586 967
rect 12390 937 12418 938
rect 12390 911 12391 937
rect 12391 911 12417 937
rect 12417 911 12418 937
rect 12390 910 12418 911
rect 13510 6846 13538 6874
rect 13454 5838 13482 5866
rect 14126 6790 14154 6818
rect 13566 6566 13594 6594
rect 14910 6734 14938 6762
rect 13790 6510 13818 6538
rect 13734 6033 13762 6034
rect 13734 6007 13735 6033
rect 13735 6007 13761 6033
rect 13761 6007 13762 6033
rect 13734 6006 13762 6007
rect 13678 5838 13706 5866
rect 13622 5614 13650 5642
rect 13174 3766 13202 3794
rect 13118 3401 13146 3402
rect 13118 3375 13119 3401
rect 13119 3375 13145 3401
rect 13145 3375 13146 3401
rect 13118 3374 13146 3375
rect 13342 3681 13370 3682
rect 13342 3655 13343 3681
rect 13343 3655 13369 3681
rect 13369 3655 13370 3681
rect 13342 3654 13370 3655
rect 13230 2926 13258 2954
rect 14126 6342 14154 6370
rect 13958 5977 13986 5978
rect 13958 5951 13959 5977
rect 13959 5951 13985 5977
rect 13985 5951 13986 5977
rect 13958 5950 13986 5951
rect 13846 5670 13874 5698
rect 13846 5278 13874 5306
rect 13902 5166 13930 5194
rect 13902 4774 13930 4802
rect 14014 4494 14042 4522
rect 13902 3262 13930 3290
rect 13846 3038 13874 3066
rect 13902 2646 13930 2674
rect 13902 2086 13930 2114
rect 13286 1777 13314 1778
rect 13286 1751 13287 1777
rect 13287 1751 13313 1777
rect 13313 1751 13314 1777
rect 13286 1750 13314 1751
rect 13678 1777 13706 1778
rect 13678 1751 13679 1777
rect 13679 1751 13705 1777
rect 13705 1751 13706 1777
rect 13678 1750 13706 1751
rect 13846 1694 13874 1722
rect 13118 1414 13146 1442
rect 11382 489 11410 490
rect 11382 463 11383 489
rect 11383 463 11409 489
rect 11409 463 11410 489
rect 11382 462 11410 463
rect 11326 350 11354 378
rect 12166 601 12194 602
rect 12166 575 12167 601
rect 12167 575 12193 601
rect 12193 575 12194 601
rect 12166 574 12194 575
rect 12110 406 12138 434
rect 12232 405 12260 406
rect 12232 379 12233 405
rect 12233 379 12259 405
rect 12259 379 12260 405
rect 12232 378 12260 379
rect 12284 405 12312 406
rect 12284 379 12285 405
rect 12285 379 12311 405
rect 12311 379 12312 405
rect 12284 378 12312 379
rect 12336 405 12364 406
rect 12336 379 12337 405
rect 12337 379 12363 405
rect 12363 379 12364 405
rect 12336 378 12364 379
rect 12446 238 12474 266
rect 12950 545 12978 546
rect 12950 519 12951 545
rect 12951 519 12977 545
rect 12977 519 12978 545
rect 12950 518 12978 519
rect 13342 1022 13370 1050
rect 13622 686 13650 714
rect 13342 462 13370 490
rect 14014 2814 14042 2842
rect 13958 1694 13986 1722
rect 14014 2198 14042 2226
rect 13902 1358 13930 1386
rect 14518 6201 14546 6202
rect 14518 6175 14519 6201
rect 14519 6175 14545 6201
rect 14545 6175 14546 6201
rect 14518 6174 14546 6175
rect 14238 5305 14266 5306
rect 14238 5279 14239 5305
rect 14239 5279 14265 5305
rect 14265 5279 14266 5305
rect 14238 5278 14266 5279
rect 14294 5166 14322 5194
rect 14294 4521 14322 4522
rect 14294 4495 14295 4521
rect 14295 4495 14321 4521
rect 14321 4495 14322 4521
rect 14294 4494 14322 4495
rect 14182 1806 14210 1834
rect 14014 1358 14042 1386
rect 13734 70 13762 98
rect 13902 70 13930 98
rect 14070 70 14098 98
rect 9758 14 9786 42
rect 14406 5390 14434 5418
rect 14518 4830 14546 4858
rect 15022 5977 15050 5978
rect 15022 5951 15023 5977
rect 15023 5951 15049 5977
rect 15049 5951 15050 5977
rect 15022 5950 15050 5951
rect 15302 5894 15330 5922
rect 14686 5334 14714 5362
rect 14686 4969 14714 4970
rect 14686 4943 14687 4969
rect 14687 4943 14713 4969
rect 14713 4943 14714 4969
rect 14686 4942 14714 4943
rect 14686 4465 14714 4466
rect 14686 4439 14687 4465
rect 14687 4439 14713 4465
rect 14713 4439 14714 4465
rect 14686 4438 14714 4439
rect 15190 4942 15218 4970
rect 15078 4718 15106 4746
rect 15190 4494 15218 4522
rect 15078 4270 15106 4298
rect 14742 4214 14770 4242
rect 14686 4129 14714 4130
rect 14686 4103 14687 4129
rect 14687 4103 14713 4129
rect 14713 4103 14714 4129
rect 14686 4102 14714 4103
rect 14630 4046 14658 4074
rect 14350 3486 14378 3514
rect 15134 4046 15162 4074
rect 14686 3822 14714 3850
rect 15190 3822 15218 3850
rect 14742 3598 14770 3626
rect 14406 3150 14434 3178
rect 15190 3598 15218 3626
rect 15134 3374 15162 3402
rect 15078 2926 15106 2954
rect 14742 2590 14770 2618
rect 14686 2561 14714 2562
rect 14686 2535 14687 2561
rect 14687 2535 14713 2561
rect 14713 2535 14714 2561
rect 14686 2534 14714 2535
rect 14406 2505 14434 2506
rect 14406 2479 14407 2505
rect 14407 2479 14433 2505
rect 14433 2479 14434 2505
rect 14406 2478 14434 2479
rect 14686 2169 14714 2170
rect 14686 2143 14687 2169
rect 14687 2143 14713 2169
rect 14713 2143 14714 2169
rect 14686 2142 14714 2143
rect 14294 1833 14322 1834
rect 14294 1807 14295 1833
rect 14295 1807 14321 1833
rect 14321 1807 14322 1833
rect 14294 1806 14322 1807
rect 14294 1694 14322 1722
rect 15134 2702 15162 2730
rect 15190 2254 15218 2282
rect 15134 2030 15162 2058
rect 14742 1638 14770 1666
rect 14686 1385 14714 1386
rect 14686 1359 14687 1385
rect 14687 1359 14713 1385
rect 14713 1359 14714 1385
rect 14686 1358 14714 1359
rect 14406 1134 14434 1162
rect 14350 910 14378 938
rect 14686 1078 14714 1106
rect 15078 1582 15106 1610
rect 15190 1358 15218 1386
<< metal3 >>
rect 4774 7014 7742 7042
rect 7770 7014 7775 7042
rect 13001 7014 13006 7042
rect 13034 7014 13398 7042
rect 13426 7014 13431 7042
rect 0 6986 56 7000
rect 4774 6986 4802 7014
rect 15792 6986 15848 7000
rect 0 6958 126 6986
rect 154 6958 159 6986
rect 4769 6958 4774 6986
rect 4802 6958 4807 6986
rect 4993 6958 4998 6986
rect 5026 6958 7070 6986
rect 7098 6958 7103 6986
rect 12833 6958 12838 6986
rect 12866 6958 15848 6986
rect 0 6944 56 6958
rect 15792 6944 15848 6958
rect 2081 6902 2086 6930
rect 2114 6902 6734 6930
rect 6762 6902 6767 6930
rect 8241 6902 8246 6930
rect 8274 6902 8638 6930
rect 8666 6902 8671 6930
rect 11545 6902 11550 6930
rect 11578 6902 12950 6930
rect 12978 6902 12983 6930
rect 1857 6846 1862 6874
rect 1890 6846 3822 6874
rect 3850 6846 3855 6874
rect 4881 6846 4886 6874
rect 4914 6846 5838 6874
rect 5866 6846 5871 6874
rect 12329 6846 12334 6874
rect 12362 6846 13510 6874
rect 13538 6846 13543 6874
rect 3761 6790 3766 6818
rect 3794 6790 5054 6818
rect 5082 6790 5087 6818
rect 6561 6790 6566 6818
rect 6594 6790 8414 6818
rect 8442 6790 8447 6818
rect 12217 6790 12222 6818
rect 12250 6790 14126 6818
rect 14154 6790 14159 6818
rect 0 6762 56 6776
rect 15792 6762 15848 6776
rect 0 6734 10262 6762
rect 10290 6734 10295 6762
rect 10425 6734 10430 6762
rect 10458 6734 12474 6762
rect 12889 6734 12894 6762
rect 12922 6734 14910 6762
rect 14938 6734 14943 6762
rect 15022 6734 15848 6762
rect 0 6720 56 6734
rect 12446 6706 12474 6734
rect 15022 6706 15050 6734
rect 15792 6720 15848 6734
rect 4153 6678 4158 6706
rect 4186 6678 5166 6706
rect 5194 6678 5199 6706
rect 5945 6678 5950 6706
rect 5978 6678 6342 6706
rect 6370 6678 6375 6706
rect 7345 6678 7350 6706
rect 7378 6678 7854 6706
rect 7882 6678 7887 6706
rect 8689 6678 8694 6706
rect 8722 6678 9198 6706
rect 9226 6678 9506 6706
rect 12446 6678 15050 6706
rect 2227 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2369 6678
rect 9478 6650 9506 6678
rect 12227 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12369 6678
rect 2977 6622 2982 6650
rect 3010 6622 4382 6650
rect 4410 6622 4415 6650
rect 5665 6622 5670 6650
rect 5698 6622 6286 6650
rect 6314 6622 6319 6650
rect 9473 6622 9478 6650
rect 9506 6622 9511 6650
rect 10985 6622 10990 6650
rect 11018 6622 11382 6650
rect 11410 6622 11415 6650
rect 1073 6566 1078 6594
rect 1106 6566 3150 6594
rect 3178 6566 3183 6594
rect 3257 6566 3262 6594
rect 3290 6566 5922 6594
rect 6617 6566 6622 6594
rect 6650 6566 7014 6594
rect 7042 6566 7047 6594
rect 7849 6566 7854 6594
rect 7882 6566 8134 6594
rect 8162 6566 8526 6594
rect 8554 6566 8559 6594
rect 10873 6566 10878 6594
rect 10906 6566 11270 6594
rect 11298 6566 11303 6594
rect 11993 6566 11998 6594
rect 12026 6566 13566 6594
rect 13594 6566 13599 6594
rect 0 6538 56 6552
rect 5894 6538 5922 6566
rect 15792 6538 15848 6552
rect 0 6510 5782 6538
rect 5810 6510 5815 6538
rect 5894 6510 7574 6538
rect 7602 6510 7607 6538
rect 8843 6510 8862 6538
rect 8890 6510 8895 6538
rect 11097 6510 11102 6538
rect 11130 6510 12222 6538
rect 12250 6510 12255 6538
rect 13785 6510 13790 6538
rect 13818 6510 15848 6538
rect 0 6496 56 6510
rect 15792 6496 15848 6510
rect 4942 6454 8078 6482
rect 8106 6454 8111 6482
rect 9305 6454 9310 6482
rect 9338 6454 9758 6482
rect 9786 6454 9791 6482
rect 11657 6454 11662 6482
rect 11690 6454 12950 6482
rect 12978 6454 12983 6482
rect 0 6314 56 6328
rect 0 6286 1246 6314
rect 1274 6286 1279 6314
rect 0 6272 56 6286
rect 1897 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2039 6286
rect 3649 6230 3654 6258
rect 3682 6230 4718 6258
rect 4746 6230 4751 6258
rect 1913 6174 1918 6202
rect 1946 6174 3374 6202
rect 3402 6174 3407 6202
rect 4209 6174 4214 6202
rect 4242 6174 4606 6202
rect 4634 6174 4639 6202
rect 4942 6146 4970 6454
rect 6673 6398 6678 6426
rect 6706 6398 8974 6426
rect 9002 6398 9007 6426
rect 10537 6398 10542 6426
rect 10570 6398 12166 6426
rect 12194 6398 12199 6426
rect 12721 6398 12726 6426
rect 12754 6398 13006 6426
rect 13034 6398 13039 6426
rect 7121 6342 7126 6370
rect 7154 6342 9702 6370
rect 9730 6342 9735 6370
rect 10873 6342 10878 6370
rect 10906 6342 11942 6370
rect 11970 6342 11975 6370
rect 12553 6342 12558 6370
rect 12586 6342 14126 6370
rect 14154 6342 14159 6370
rect 15792 6314 15848 6328
rect 5161 6286 5166 6314
rect 5194 6286 8806 6314
rect 8834 6286 8839 6314
rect 9193 6286 9198 6314
rect 9226 6286 9534 6314
rect 9562 6286 9567 6314
rect 12721 6286 12726 6314
rect 12754 6286 15848 6314
rect 11897 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12039 6286
rect 15792 6272 15848 6286
rect 5945 6230 5950 6258
rect 5978 6230 10038 6258
rect 10066 6230 10071 6258
rect 5049 6174 5054 6202
rect 5082 6174 5614 6202
rect 5642 6174 5647 6202
rect 6001 6174 6006 6202
rect 6034 6174 6174 6202
rect 6202 6174 6207 6202
rect 7233 6174 7238 6202
rect 7266 6174 8862 6202
rect 8890 6174 8895 6202
rect 11321 6174 11326 6202
rect 11354 6174 11998 6202
rect 12026 6174 12031 6202
rect 12665 6174 12670 6202
rect 12698 6174 14518 6202
rect 14546 6174 14551 6202
rect 2585 6118 2590 6146
rect 2618 6118 2758 6146
rect 2786 6118 4970 6146
rect 5161 6118 5166 6146
rect 5194 6118 5502 6146
rect 5530 6118 5535 6146
rect 6505 6118 6510 6146
rect 6538 6118 6790 6146
rect 6818 6118 6823 6146
rect 7009 6118 7014 6146
rect 7042 6118 9254 6146
rect 9282 6118 9287 6146
rect 0 6090 56 6104
rect 15792 6090 15848 6104
rect 0 6062 70 6090
rect 98 6062 103 6090
rect 3761 6062 3766 6090
rect 3794 6062 8750 6090
rect 8778 6062 8783 6090
rect 8857 6062 8862 6090
rect 8890 6062 8974 6090
rect 9002 6062 9142 6090
rect 9170 6062 9175 6090
rect 10481 6062 10486 6090
rect 10514 6062 15848 6090
rect 0 6048 56 6062
rect 15792 6048 15848 6062
rect 2193 6006 2198 6034
rect 2226 6006 4494 6034
rect 4522 6006 4527 6034
rect 5329 6006 5334 6034
rect 5362 6006 9926 6034
rect 9954 6006 9959 6034
rect 10537 6006 10542 6034
rect 10570 6006 10766 6034
rect 10794 6006 10799 6034
rect 12497 6006 12502 6034
rect 12530 6006 13734 6034
rect 13762 6006 13767 6034
rect 2982 5950 5502 5978
rect 5530 5950 5535 5978
rect 5777 5950 5782 5978
rect 5810 5950 9366 5978
rect 9394 5950 10150 5978
rect 10178 5950 10183 5978
rect 10257 5950 10262 5978
rect 10290 5950 10710 5978
rect 10738 5950 11130 5978
rect 12777 5950 12782 5978
rect 12810 5950 13174 5978
rect 13202 5950 13207 5978
rect 13953 5950 13958 5978
rect 13986 5950 15022 5978
rect 15050 5950 15055 5978
rect 2982 5922 3010 5950
rect 11102 5922 11130 5950
rect 2977 5894 2982 5922
rect 3010 5894 3015 5922
rect 4545 5894 4550 5922
rect 4578 5894 7406 5922
rect 7434 5894 7439 5922
rect 7681 5894 7686 5922
rect 7714 5894 8078 5922
rect 8106 5894 8111 5922
rect 9529 5894 9534 5922
rect 9562 5894 9758 5922
rect 9786 5894 9791 5922
rect 10761 5894 10766 5922
rect 10794 5894 10878 5922
rect 10906 5894 10911 5922
rect 11097 5894 11102 5922
rect 11130 5894 11135 5922
rect 13113 5894 13118 5922
rect 13146 5894 15302 5922
rect 15330 5894 15335 5922
rect 0 5866 56 5880
rect 2227 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2369 5894
rect 12227 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12369 5894
rect 15792 5866 15848 5880
rect 0 5838 1078 5866
rect 1106 5838 1111 5866
rect 3089 5838 3094 5866
rect 3122 5838 3878 5866
rect 3906 5838 3911 5866
rect 4657 5838 4662 5866
rect 4690 5838 5838 5866
rect 5866 5838 5871 5866
rect 10425 5838 10430 5866
rect 10458 5838 11158 5866
rect 11186 5838 11191 5866
rect 12665 5838 12670 5866
rect 12698 5838 12894 5866
rect 12922 5838 12927 5866
rect 13449 5838 13454 5866
rect 13482 5838 13487 5866
rect 13673 5838 13678 5866
rect 13706 5838 15848 5866
rect 0 5824 56 5838
rect 1801 5782 1806 5810
rect 1834 5782 9954 5810
rect 11209 5782 11214 5810
rect 11242 5782 11606 5810
rect 11634 5782 11639 5810
rect 9926 5754 9954 5782
rect 13454 5754 13482 5838
rect 15792 5824 15848 5838
rect 2305 5726 2310 5754
rect 2338 5726 3206 5754
rect 3234 5726 3239 5754
rect 6785 5726 6790 5754
rect 6818 5726 7462 5754
rect 7490 5726 7495 5754
rect 9081 5726 9086 5754
rect 9114 5726 9814 5754
rect 9842 5726 9847 5754
rect 9926 5726 11550 5754
rect 11578 5726 11583 5754
rect 11657 5726 11662 5754
rect 11690 5726 13482 5754
rect 2417 5670 2422 5698
rect 2450 5670 2870 5698
rect 2898 5670 2903 5698
rect 4153 5670 4158 5698
rect 4186 5670 6286 5698
rect 6314 5670 6319 5698
rect 10425 5670 10430 5698
rect 10458 5670 11494 5698
rect 11522 5670 11527 5698
rect 11606 5670 13846 5698
rect 13874 5670 13879 5698
rect 0 5642 56 5656
rect 11606 5642 11634 5670
rect 15792 5642 15848 5656
rect 0 5614 686 5642
rect 714 5614 719 5642
rect 1801 5614 1806 5642
rect 1834 5614 2702 5642
rect 2730 5614 2735 5642
rect 3873 5614 3878 5642
rect 3906 5614 4438 5642
rect 4466 5614 4471 5642
rect 5665 5614 5670 5642
rect 5698 5614 7294 5642
rect 7322 5614 7327 5642
rect 7905 5614 7910 5642
rect 7938 5614 9030 5642
rect 9058 5614 9063 5642
rect 10467 5614 10486 5642
rect 10514 5614 10519 5642
rect 10649 5614 10654 5642
rect 10682 5614 11634 5642
rect 11769 5614 11774 5642
rect 11802 5614 12558 5642
rect 12586 5614 12591 5642
rect 13617 5614 13622 5642
rect 13650 5614 15848 5642
rect 0 5600 56 5614
rect 15792 5600 15848 5614
rect 5217 5558 5222 5586
rect 5250 5558 9310 5586
rect 9338 5558 9343 5586
rect 10089 5558 10094 5586
rect 10122 5558 10430 5586
rect 10458 5558 10463 5586
rect 11825 5558 11830 5586
rect 11858 5558 12614 5586
rect 12642 5558 12647 5586
rect 3089 5502 3094 5530
rect 3122 5502 3486 5530
rect 3514 5502 3519 5530
rect 4186 5502 8302 5530
rect 8330 5502 8335 5530
rect 9361 5502 9366 5530
rect 9394 5502 11662 5530
rect 11690 5502 11695 5530
rect 1897 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2039 5502
rect 4153 5446 4158 5474
rect 4186 5446 4214 5502
rect 11897 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12039 5502
rect 7121 5446 7126 5474
rect 7154 5446 7462 5474
rect 7490 5446 7630 5474
rect 7658 5446 7663 5474
rect 12105 5446 12110 5474
rect 12138 5446 12558 5474
rect 12586 5446 12591 5474
rect 0 5418 56 5432
rect 15792 5418 15848 5432
rect 0 5390 2114 5418
rect 3481 5390 3486 5418
rect 3514 5390 4046 5418
rect 4074 5390 4079 5418
rect 7401 5390 7406 5418
rect 7434 5390 7686 5418
rect 7714 5390 7966 5418
rect 7994 5390 7999 5418
rect 9977 5390 9982 5418
rect 10010 5390 10150 5418
rect 10178 5390 10183 5418
rect 11433 5390 11438 5418
rect 11466 5390 11830 5418
rect 11858 5390 11863 5418
rect 14401 5390 14406 5418
rect 14434 5390 15848 5418
rect 0 5376 56 5390
rect 2086 5306 2114 5390
rect 15792 5376 15848 5390
rect 2585 5334 2590 5362
rect 2618 5334 2758 5362
rect 2786 5334 5222 5362
rect 5250 5334 5255 5362
rect 5329 5334 5334 5362
rect 5362 5334 11326 5362
rect 11354 5334 11359 5362
rect 11433 5334 11438 5362
rect 11466 5334 14686 5362
rect 14714 5334 14719 5362
rect 2086 5278 4214 5306
rect 4242 5278 4247 5306
rect 4825 5278 4830 5306
rect 4858 5278 5222 5306
rect 5250 5278 5255 5306
rect 6449 5278 6454 5306
rect 6482 5278 6734 5306
rect 6762 5278 6767 5306
rect 10369 5278 10374 5306
rect 10402 5278 10654 5306
rect 10682 5278 10687 5306
rect 10985 5278 10990 5306
rect 11018 5278 11158 5306
rect 11186 5278 11191 5306
rect 11769 5278 11774 5306
rect 11802 5278 12278 5306
rect 12306 5278 12311 5306
rect 13841 5278 13846 5306
rect 13874 5278 14238 5306
rect 14266 5278 14271 5306
rect 6113 5222 6118 5250
rect 6146 5222 9254 5250
rect 9282 5222 9287 5250
rect 11097 5222 11102 5250
rect 11130 5222 12334 5250
rect 12362 5222 12367 5250
rect 0 5194 56 5208
rect 15792 5194 15848 5208
rect 0 5166 406 5194
rect 434 5166 439 5194
rect 1353 5166 1358 5194
rect 1386 5166 7182 5194
rect 7210 5166 7215 5194
rect 11153 5166 11158 5194
rect 11186 5166 13902 5194
rect 13930 5166 13935 5194
rect 14289 5166 14294 5194
rect 14322 5166 15848 5194
rect 0 5152 56 5166
rect 15792 5152 15848 5166
rect 6169 5110 6174 5138
rect 6202 5110 7518 5138
rect 7546 5110 7551 5138
rect 8409 5110 8414 5138
rect 8442 5110 11438 5138
rect 11466 5110 11471 5138
rect 2227 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2369 5110
rect 12227 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12369 5110
rect 9921 5054 9926 5082
rect 9954 5054 11774 5082
rect 11802 5054 11807 5082
rect 2137 4998 2142 5026
rect 2170 4998 4438 5026
rect 4466 4998 4471 5026
rect 10817 4998 10822 5026
rect 10850 4998 11718 5026
rect 11746 4998 11751 5026
rect 12609 4998 12614 5026
rect 12642 4998 13062 5026
rect 13090 4998 13095 5026
rect 0 4970 56 4984
rect 15792 4970 15848 4984
rect 0 4942 5054 4970
rect 5082 4942 5087 4970
rect 7961 4942 7966 4970
rect 7994 4942 14686 4970
rect 14714 4942 14719 4970
rect 15185 4942 15190 4970
rect 15218 4942 15848 4970
rect 0 4928 56 4942
rect 15792 4928 15848 4942
rect 401 4886 406 4914
rect 434 4886 2646 4914
rect 2674 4886 2679 4914
rect 3313 4886 3318 4914
rect 3346 4886 5950 4914
rect 5978 4886 5983 4914
rect 6113 4886 6118 4914
rect 6146 4886 10878 4914
rect 10906 4886 10911 4914
rect 11601 4886 11606 4914
rect 11634 4886 12278 4914
rect 12306 4886 12311 4914
rect 2529 4830 2534 4858
rect 2562 4830 6902 4858
rect 6930 4830 6935 4858
rect 7457 4830 7462 4858
rect 7490 4830 7686 4858
rect 7714 4830 7719 4858
rect 7961 4830 7966 4858
rect 7994 4830 8134 4858
rect 8162 4830 8167 4858
rect 11377 4830 11382 4858
rect 11410 4830 11662 4858
rect 11690 4830 11942 4858
rect 11970 4830 11975 4858
rect 12105 4830 12110 4858
rect 12138 4830 14518 4858
rect 14546 4830 14551 4858
rect 3593 4774 3598 4802
rect 3626 4774 3878 4802
rect 3906 4774 3911 4802
rect 8297 4774 8302 4802
rect 8330 4774 13902 4802
rect 13930 4774 13935 4802
rect 0 4746 56 4760
rect 15792 4746 15848 4760
rect 0 4718 910 4746
rect 938 4718 943 4746
rect 4097 4718 4102 4746
rect 4130 4718 5726 4746
rect 5754 4718 5759 4746
rect 15073 4718 15078 4746
rect 15106 4718 15848 4746
rect 0 4704 56 4718
rect 1897 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2039 4718
rect 11897 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12039 4718
rect 15792 4704 15848 4718
rect 6673 4662 6678 4690
rect 6706 4662 6902 4690
rect 6930 4662 6935 4690
rect 4769 4606 4774 4634
rect 4802 4606 7854 4634
rect 7882 4606 7887 4634
rect 10033 4606 10038 4634
rect 10066 4606 12446 4634
rect 12474 4606 12479 4634
rect 5329 4550 5334 4578
rect 5362 4550 12110 4578
rect 12138 4550 12143 4578
rect 0 4522 56 4536
rect 15792 4522 15848 4536
rect 0 4494 7462 4522
rect 7490 4494 7495 4522
rect 14009 4494 14014 4522
rect 14042 4494 14294 4522
rect 14322 4494 14327 4522
rect 15185 4494 15190 4522
rect 15218 4494 15848 4522
rect 0 4480 56 4494
rect 15792 4480 15848 4494
rect 1857 4438 1862 4466
rect 1890 4438 2590 4466
rect 2618 4438 2623 4466
rect 4153 4438 4158 4466
rect 4186 4438 5726 4466
rect 5754 4438 5759 4466
rect 8353 4438 8358 4466
rect 8386 4438 14686 4466
rect 14714 4438 14719 4466
rect 905 4382 910 4410
rect 938 4382 7406 4410
rect 7434 4382 7574 4410
rect 7602 4382 7607 4410
rect 10649 4382 10654 4410
rect 10682 4382 11326 4410
rect 11354 4382 11359 4410
rect 11545 4382 11550 4410
rect 11578 4382 12614 4410
rect 12642 4382 12647 4410
rect 5273 4326 5278 4354
rect 5306 4326 5614 4354
rect 5642 4326 6790 4354
rect 6818 4326 6823 4354
rect 7294 4326 11830 4354
rect 11858 4326 11863 4354
rect 0 4298 56 4312
rect 2227 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2369 4326
rect 7294 4298 7322 4326
rect 12227 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12369 4326
rect 15792 4298 15848 4312
rect 0 4270 2114 4298
rect 3257 4270 3262 4298
rect 3290 4270 5502 4298
rect 5530 4270 5535 4298
rect 5833 4270 5838 4298
rect 5866 4270 7322 4298
rect 7546 4270 7966 4298
rect 7994 4270 7999 4298
rect 9585 4270 9590 4298
rect 9618 4270 10934 4298
rect 10962 4270 10967 4298
rect 15073 4270 15078 4298
rect 15106 4270 15848 4298
rect 0 4256 56 4270
rect 2086 4242 2114 4270
rect 7546 4242 7574 4270
rect 15792 4256 15848 4270
rect 2086 4214 7574 4242
rect 7849 4214 7854 4242
rect 7882 4214 14742 4242
rect 14770 4214 14775 4242
rect 6225 4158 6230 4186
rect 6258 4158 6398 4186
rect 6426 4158 7630 4186
rect 7658 4158 7663 4186
rect 1577 4102 1582 4130
rect 1610 4102 3486 4130
rect 3514 4102 3519 4130
rect 5777 4102 5782 4130
rect 5810 4102 7070 4130
rect 7098 4102 7103 4130
rect 8465 4102 8470 4130
rect 8498 4102 14686 4130
rect 14714 4102 14719 4130
rect 0 4074 56 4088
rect 5950 4074 5978 4102
rect 15792 4074 15848 4088
rect 0 4046 2534 4074
rect 2562 4046 2567 4074
rect 3985 4046 3990 4074
rect 4018 4046 5054 4074
rect 5082 4046 5087 4074
rect 5945 4046 5950 4074
rect 5978 4046 5983 4074
rect 8073 4046 8078 4074
rect 8106 4046 14630 4074
rect 14658 4046 14663 4074
rect 15129 4046 15134 4074
rect 15162 4046 15848 4074
rect 0 4032 56 4046
rect 15792 4032 15848 4046
rect 5553 3990 5558 4018
rect 5586 3990 10766 4018
rect 10794 3990 10799 4018
rect 2585 3934 2590 3962
rect 2618 3934 2758 3962
rect 2786 3934 6846 3962
rect 6874 3934 6879 3962
rect 7546 3934 9926 3962
rect 9954 3934 9959 3962
rect 1897 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2039 3934
rect 7546 3906 7574 3934
rect 11897 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12039 3934
rect 2473 3878 2478 3906
rect 2506 3878 5166 3906
rect 5194 3878 5199 3906
rect 6897 3878 6902 3906
rect 6930 3878 7574 3906
rect 9025 3878 9030 3906
rect 9058 3878 11186 3906
rect 0 3850 56 3864
rect 11158 3850 11186 3878
rect 15792 3850 15848 3864
rect 0 3822 2534 3850
rect 2562 3822 2567 3850
rect 7966 3822 9310 3850
rect 9338 3822 9343 3850
rect 10033 3822 10038 3850
rect 10066 3822 11046 3850
rect 11074 3822 11079 3850
rect 11158 3822 14686 3850
rect 14714 3822 14719 3850
rect 15185 3822 15190 3850
rect 15218 3822 15848 3850
rect 0 3808 56 3822
rect 5049 3766 5054 3794
rect 5082 3766 7686 3794
rect 7714 3766 7798 3794
rect 7826 3766 7831 3794
rect 7966 3738 7994 3822
rect 15792 3808 15848 3822
rect 8073 3766 8078 3794
rect 8106 3766 8414 3794
rect 8442 3766 8447 3794
rect 12105 3766 12110 3794
rect 12138 3766 13174 3794
rect 13202 3766 13207 3794
rect 3817 3710 3822 3738
rect 3850 3710 6958 3738
rect 6986 3710 6991 3738
rect 7546 3710 7994 3738
rect 8241 3710 8246 3738
rect 8274 3710 12894 3738
rect 12922 3710 12927 3738
rect 7546 3682 7574 3710
rect 4321 3654 4326 3682
rect 4354 3654 4438 3682
rect 4466 3654 7574 3682
rect 8913 3654 8918 3682
rect 8946 3654 13342 3682
rect 13370 3654 13375 3682
rect 0 3626 56 3640
rect 15792 3626 15848 3640
rect 0 3598 2450 3626
rect 7625 3598 7630 3626
rect 7658 3598 14742 3626
rect 14770 3598 14775 3626
rect 15185 3598 15190 3626
rect 15218 3598 15848 3626
rect 0 3584 56 3598
rect 2227 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2369 3542
rect 2422 3514 2450 3598
rect 15792 3584 15848 3598
rect 2529 3542 2534 3570
rect 2562 3542 7126 3570
rect 7154 3542 7159 3570
rect 12227 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12369 3542
rect 2422 3486 7574 3514
rect 7602 3486 7607 3514
rect 12945 3486 12950 3514
rect 12978 3486 14350 3514
rect 14378 3486 14383 3514
rect 681 3430 686 3458
rect 714 3430 3374 3458
rect 3402 3430 3407 3458
rect 3873 3430 3878 3458
rect 3906 3430 4942 3458
rect 4970 3430 4975 3458
rect 9193 3430 9198 3458
rect 9226 3430 11102 3458
rect 11130 3430 11135 3458
rect 0 3402 56 3416
rect 15792 3402 15848 3416
rect 0 3374 7238 3402
rect 7266 3374 7271 3402
rect 10481 3374 10486 3402
rect 10514 3374 13118 3402
rect 13146 3374 13151 3402
rect 15129 3374 15134 3402
rect 15162 3374 15848 3402
rect 0 3360 56 3374
rect 15792 3360 15848 3374
rect 4433 3318 4438 3346
rect 4466 3318 7966 3346
rect 7994 3318 7999 3346
rect 8073 3318 8078 3346
rect 8106 3318 8358 3346
rect 8386 3318 8391 3346
rect 1806 3262 7014 3290
rect 7042 3262 7182 3290
rect 7210 3262 7215 3290
rect 7457 3262 7462 3290
rect 7490 3262 13902 3290
rect 13930 3262 13935 3290
rect 0 3178 56 3192
rect 1806 3178 1834 3262
rect 4153 3206 4158 3234
rect 4186 3206 4438 3234
rect 4466 3206 4471 3234
rect 15792 3178 15848 3192
rect 0 3150 1834 3178
rect 14401 3150 14406 3178
rect 14434 3150 15848 3178
rect 0 3136 56 3150
rect 1897 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2039 3150
rect 11897 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12039 3150
rect 15792 3136 15848 3150
rect 121 3038 126 3066
rect 154 3038 13846 3066
rect 13874 3038 13879 3066
rect 7513 2982 7518 3010
rect 7546 2982 8302 3010
rect 8330 2982 8335 3010
rect 0 2954 56 2968
rect 15792 2954 15848 2968
rect 0 2926 7182 2954
rect 7210 2926 7215 2954
rect 7457 2926 7462 2954
rect 7490 2926 7574 2954
rect 8129 2926 8134 2954
rect 8162 2926 13230 2954
rect 13258 2926 13263 2954
rect 15073 2926 15078 2954
rect 15106 2926 15848 2954
rect 0 2912 56 2926
rect 7546 2898 7574 2926
rect 15792 2912 15848 2926
rect 7546 2870 13006 2898
rect 13034 2870 13039 2898
rect 2641 2814 2646 2842
rect 2674 2814 7070 2842
rect 7098 2814 7238 2842
rect 7266 2814 7271 2842
rect 9137 2814 9142 2842
rect 9170 2814 14014 2842
rect 14042 2814 14047 2842
rect 0 2730 56 2744
rect 2227 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2369 2758
rect 12227 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12369 2758
rect 15792 2730 15848 2744
rect 0 2702 2114 2730
rect 4209 2702 4214 2730
rect 4242 2702 8750 2730
rect 8778 2702 8862 2730
rect 8890 2702 8895 2730
rect 15129 2702 15134 2730
rect 15162 2702 15848 2730
rect 0 2688 56 2702
rect 2086 2674 2114 2702
rect 15792 2688 15848 2702
rect 2086 2646 8022 2674
rect 8050 2646 8055 2674
rect 8689 2646 8694 2674
rect 8722 2646 13902 2674
rect 13930 2646 13935 2674
rect 8073 2590 8078 2618
rect 8106 2590 14742 2618
rect 14770 2590 14775 2618
rect 7513 2534 7518 2562
rect 7546 2534 14686 2562
rect 14714 2534 14719 2562
rect 0 2506 56 2520
rect 15792 2506 15848 2520
rect 0 2478 1414 2506
rect 1442 2478 1447 2506
rect 2529 2478 2534 2506
rect 2562 2478 8190 2506
rect 8218 2478 8223 2506
rect 14401 2478 14406 2506
rect 14434 2478 15848 2506
rect 0 2464 56 2478
rect 15792 2464 15848 2478
rect 121 2422 126 2450
rect 154 2422 10654 2450
rect 10682 2422 10687 2450
rect 1897 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2039 2366
rect 11897 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12039 2366
rect 0 2282 56 2296
rect 15792 2282 15848 2296
rect 0 2254 7630 2282
rect 7658 2254 7663 2282
rect 15185 2254 15190 2282
rect 15218 2254 15848 2282
rect 0 2240 56 2254
rect 15792 2240 15848 2254
rect 7065 2198 7070 2226
rect 7098 2198 14014 2226
rect 14042 2198 14047 2226
rect 1409 2142 1414 2170
rect 1442 2142 8302 2170
rect 8330 2142 8335 2170
rect 8633 2142 8638 2170
rect 8666 2142 14686 2170
rect 14714 2142 14719 2170
rect 7513 2086 7518 2114
rect 7546 2086 13902 2114
rect 13930 2086 13935 2114
rect 0 2058 56 2072
rect 15792 2058 15848 2072
rect 0 2030 6622 2058
rect 6650 2030 6655 2058
rect 7009 2030 7014 2058
rect 7042 2030 7294 2058
rect 7322 2030 7327 2058
rect 15129 2030 15134 2058
rect 15162 2030 15848 2058
rect 0 2016 56 2030
rect 15792 2016 15848 2030
rect 3369 1974 3374 2002
rect 3402 1974 7686 2002
rect 7714 1974 7719 2002
rect 2227 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2369 1974
rect 12227 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12369 1974
rect 1241 1862 1246 1890
rect 1274 1862 9478 1890
rect 9506 1862 9511 1890
rect 0 1834 56 1848
rect 15792 1834 15848 1848
rect 0 1806 7014 1834
rect 7042 1806 7047 1834
rect 10873 1806 10878 1834
rect 10906 1806 14182 1834
rect 14210 1806 14215 1834
rect 14289 1806 14294 1834
rect 14322 1806 15848 1834
rect 0 1792 56 1806
rect 15792 1792 15848 1806
rect 13281 1750 13286 1778
rect 13314 1750 13678 1778
rect 13706 1750 13711 1778
rect 7233 1694 7238 1722
rect 7266 1694 13846 1722
rect 13874 1694 13879 1722
rect 13953 1694 13958 1722
rect 13986 1694 14294 1722
rect 14322 1694 14327 1722
rect 1806 1638 6846 1666
rect 6874 1638 6879 1666
rect 7289 1638 7294 1666
rect 7322 1638 14742 1666
rect 14770 1638 14775 1666
rect 0 1610 56 1624
rect 1806 1610 1834 1638
rect 15792 1610 15848 1624
rect 0 1582 1834 1610
rect 15073 1582 15078 1610
rect 15106 1582 15848 1610
rect 0 1568 56 1582
rect 1897 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2039 1582
rect 11897 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12039 1582
rect 15792 1568 15848 1582
rect 1073 1470 1078 1498
rect 1106 1470 8638 1498
rect 8666 1470 8671 1498
rect 8073 1414 8078 1442
rect 8106 1414 13118 1442
rect 13146 1414 13151 1442
rect 0 1386 56 1400
rect 15792 1386 15848 1400
rect 0 1358 7518 1386
rect 7546 1358 7686 1386
rect 7714 1358 7719 1386
rect 8353 1358 8358 1386
rect 8386 1358 13902 1386
rect 13930 1358 13935 1386
rect 14009 1358 14014 1386
rect 14042 1358 14686 1386
rect 14714 1358 14719 1386
rect 15185 1358 15190 1386
rect 15218 1358 15848 1386
rect 0 1344 56 1358
rect 15792 1344 15848 1358
rect 2086 1246 8022 1274
rect 8050 1246 8134 1274
rect 8162 1246 8167 1274
rect 10705 1246 10710 1274
rect 10738 1246 10822 1274
rect 10850 1246 10855 1274
rect 0 1162 56 1176
rect 2086 1162 2114 1246
rect 2227 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2369 1190
rect 12227 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12369 1190
rect 15792 1162 15848 1176
rect 0 1134 2114 1162
rect 10593 1134 10598 1162
rect 10626 1134 11662 1162
rect 11690 1134 11695 1162
rect 14401 1134 14406 1162
rect 14434 1134 15848 1162
rect 0 1120 56 1134
rect 15792 1120 15848 1134
rect 7961 1078 7966 1106
rect 7994 1078 14686 1106
rect 14714 1078 14719 1106
rect 2086 1022 6790 1050
rect 6818 1022 6823 1050
rect 7401 1022 7406 1050
rect 7434 1022 13342 1050
rect 13370 1022 13375 1050
rect 0 938 56 952
rect 2086 938 2114 1022
rect 3145 966 3150 994
rect 3178 966 10206 994
rect 10234 966 10374 994
rect 10402 966 10407 994
rect 12553 966 12558 994
rect 12586 966 12591 994
rect 12558 938 12586 966
rect 15792 938 15848 952
rect 0 910 2114 938
rect 2142 910 9142 938
rect 9170 910 9310 938
rect 9338 910 9343 938
rect 11209 910 11214 938
rect 11242 910 12390 938
rect 12418 910 12586 938
rect 14345 910 14350 938
rect 14378 910 15848 938
rect 0 896 56 910
rect 2142 882 2170 910
rect 15792 896 15848 910
rect 1801 854 1806 882
rect 1834 854 2170 882
rect 3817 854 3822 882
rect 3850 854 10822 882
rect 10850 854 10855 882
rect 3481 798 3486 826
rect 3514 798 5166 826
rect 5194 798 5199 826
rect 6953 798 6958 826
rect 6986 798 7126 826
rect 7154 798 7159 826
rect 1897 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2039 798
rect 11897 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12039 798
rect 6337 742 6342 770
rect 6370 742 8246 770
rect 8274 742 8279 770
rect 0 714 56 728
rect 15792 714 15848 728
rect 0 686 7630 714
rect 7658 686 7663 714
rect 13617 686 13622 714
rect 13650 686 15848 714
rect 0 672 56 686
rect 15792 672 15848 686
rect 5553 630 5558 658
rect 5586 630 7462 658
rect 7490 630 7495 658
rect 8129 630 8134 658
rect 8162 630 8526 658
rect 8554 630 8559 658
rect 7849 574 7854 602
rect 7882 574 12166 602
rect 12194 574 12199 602
rect 4186 518 8134 546
rect 8162 518 8167 546
rect 8353 518 8358 546
rect 8386 518 12950 546
rect 12978 518 12983 546
rect 0 490 56 504
rect 4186 490 4214 518
rect 15792 490 15848 504
rect 0 462 4214 490
rect 7849 462 7854 490
rect 7882 462 8806 490
rect 8834 462 8918 490
rect 8946 462 8951 490
rect 11097 462 11102 490
rect 11130 462 11382 490
rect 11410 462 11415 490
rect 13337 462 13342 490
rect 13370 462 15848 490
rect 0 448 56 462
rect 15792 448 15848 462
rect 3593 406 3598 434
rect 3626 406 12110 434
rect 12138 406 12143 434
rect 2227 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2369 406
rect 12227 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12369 406
rect 8521 350 8526 378
rect 8554 350 11158 378
rect 11186 350 11326 378
rect 11354 350 11359 378
rect 4489 294 4494 322
rect 4522 294 9366 322
rect 9394 294 9399 322
rect 9865 294 9870 322
rect 9898 294 10430 322
rect 10458 294 10463 322
rect 0 266 56 280
rect 15792 266 15848 280
rect 0 238 7462 266
rect 7490 238 7495 266
rect 9193 238 9198 266
rect 9226 238 11102 266
rect 11130 238 11135 266
rect 12441 238 12446 266
rect 12474 238 15848 266
rect 0 224 56 238
rect 15792 224 15848 238
rect 1022 126 6958 154
rect 6986 126 6991 154
rect 0 42 56 56
rect 1022 42 1050 126
rect 1129 70 1134 98
rect 1162 70 1167 98
rect 2473 70 2478 98
rect 2506 70 9646 98
rect 9674 70 9679 98
rect 13729 70 13734 98
rect 13762 70 13767 98
rect 13897 70 13902 98
rect 13930 70 14070 98
rect 14098 70 14103 98
rect 0 14 1050 42
rect 1134 42 1162 70
rect 13734 42 13762 70
rect 15792 42 15848 56
rect 1134 14 9758 42
rect 9786 14 9791 42
rect 13734 14 15848 42
rect 0 0 56 14
rect 15792 0 15848 14
<< via3 >>
rect 2232 6650 2260 6678
rect 2284 6650 2312 6678
rect 2336 6650 2364 6678
rect 12232 6650 12260 6678
rect 12284 6650 12312 6678
rect 12336 6650 12364 6678
rect 5782 6510 5810 6538
rect 8862 6510 8890 6538
rect 9758 6454 9786 6482
rect 1902 6258 1930 6286
rect 1954 6258 1982 6286
rect 2006 6258 2034 6286
rect 11902 6258 11930 6286
rect 11954 6258 11982 6286
rect 12006 6258 12034 6286
rect 8862 6062 8890 6090
rect 5782 5950 5810 5978
rect 9758 5894 9786 5922
rect 2232 5866 2260 5894
rect 2284 5866 2312 5894
rect 2336 5866 2364 5894
rect 12232 5866 12260 5894
rect 12284 5866 12312 5894
rect 12336 5866 12364 5894
rect 11662 5726 11690 5754
rect 10486 5614 10514 5642
rect 5222 5558 5250 5586
rect 11662 5502 11690 5530
rect 1902 5474 1930 5502
rect 1954 5474 1982 5502
rect 2006 5474 2034 5502
rect 11902 5474 11930 5502
rect 11954 5474 11982 5502
rect 12006 5474 12034 5502
rect 5222 5334 5250 5362
rect 11438 5334 11466 5362
rect 4214 5278 4242 5306
rect 11438 5110 11466 5138
rect 2232 5082 2260 5110
rect 2284 5082 2312 5110
rect 2336 5082 2364 5110
rect 12232 5082 12260 5110
rect 12284 5082 12312 5110
rect 12336 5082 12364 5110
rect 5054 4942 5082 4970
rect 12110 4830 12138 4858
rect 1902 4690 1930 4718
rect 1954 4690 1982 4718
rect 2006 4690 2034 4718
rect 11902 4690 11930 4718
rect 11954 4690 11982 4718
rect 12006 4690 12034 4718
rect 12110 4550 12138 4578
rect 2232 4298 2260 4326
rect 2284 4298 2312 4326
rect 2336 4298 2364 4326
rect 12232 4298 12260 4326
rect 12284 4298 12312 4326
rect 12336 4298 12364 4326
rect 2534 4046 2562 4074
rect 1902 3906 1930 3934
rect 1954 3906 1982 3934
rect 2006 3906 2034 3934
rect 11902 3906 11930 3934
rect 11954 3906 11982 3934
rect 12006 3906 12034 3934
rect 5054 3766 5082 3794
rect 2232 3514 2260 3542
rect 2284 3514 2312 3542
rect 2336 3514 2364 3542
rect 2534 3542 2562 3570
rect 12232 3514 12260 3542
rect 12284 3514 12312 3542
rect 12336 3514 12364 3542
rect 10486 3374 10514 3402
rect 1902 3122 1930 3150
rect 1954 3122 1982 3150
rect 2006 3122 2034 3150
rect 11902 3122 11930 3150
rect 11954 3122 11982 3150
rect 12006 3122 12034 3150
rect 2232 2730 2260 2758
rect 2284 2730 2312 2758
rect 2336 2730 2364 2758
rect 12232 2730 12260 2758
rect 12284 2730 12312 2758
rect 12336 2730 12364 2758
rect 4214 2702 4242 2730
rect 1902 2338 1930 2366
rect 1954 2338 1982 2366
rect 2006 2338 2034 2366
rect 11902 2338 11930 2366
rect 11954 2338 11982 2366
rect 12006 2338 12034 2366
rect 2232 1946 2260 1974
rect 2284 1946 2312 1974
rect 2336 1946 2364 1974
rect 12232 1946 12260 1974
rect 12284 1946 12312 1974
rect 12336 1946 12364 1974
rect 1902 1554 1930 1582
rect 1954 1554 1982 1582
rect 2006 1554 2034 1582
rect 11902 1554 11930 1582
rect 11954 1554 11982 1582
rect 12006 1554 12034 1582
rect 2232 1162 2260 1190
rect 2284 1162 2312 1190
rect 2336 1162 2364 1190
rect 12232 1162 12260 1190
rect 12284 1162 12312 1190
rect 12336 1162 12364 1190
rect 1902 770 1930 798
rect 1954 770 1982 798
rect 2006 770 2034 798
rect 11902 770 11930 798
rect 11954 770 11982 798
rect 12006 770 12034 798
rect 2232 378 2260 406
rect 2284 378 2312 406
rect 2336 378 2364 406
rect 12232 378 12260 406
rect 12284 378 12312 406
rect 12336 378 12364 406
<< metal4 >>
rect 1888 6286 2048 7112
rect 1888 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2048 6286
rect 1888 5502 2048 6258
rect 1888 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2048 5502
rect 1888 4718 2048 5474
rect 1888 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2048 4718
rect 1888 3934 2048 4690
rect 1888 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2048 3934
rect 1888 3150 2048 3906
rect 1888 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2048 3150
rect 1888 2366 2048 3122
rect 1888 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2048 2366
rect 1888 1582 2048 2338
rect 1888 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2048 1582
rect 1888 798 2048 1554
rect 1888 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2048 798
rect 1888 0 2048 770
rect 2218 6678 2378 7112
rect 2218 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2378 6678
rect 2218 5894 2378 6650
rect 5782 6538 5810 6543
rect 5782 5978 5810 6510
rect 8862 6538 8890 6543
rect 8862 6090 8890 6510
rect 8862 6057 8890 6062
rect 9758 6482 9786 6487
rect 5782 5945 5810 5950
rect 2218 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2378 5894
rect 9758 5922 9786 6454
rect 9758 5889 9786 5894
rect 11888 6286 12048 7112
rect 11888 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12048 6286
rect 2218 5110 2378 5866
rect 11662 5754 11690 5759
rect 10486 5642 10514 5647
rect 5222 5586 5250 5591
rect 5222 5362 5250 5558
rect 5222 5329 5250 5334
rect 2218 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2378 5110
rect 2218 4326 2378 5082
rect 2218 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2378 4326
rect 2218 3542 2378 4298
rect 4214 5306 4242 5311
rect 2218 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2378 3542
rect 2534 4074 2562 4079
rect 2534 3570 2562 4046
rect 2534 3537 2562 3542
rect 2218 2758 2378 3514
rect 2218 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2378 2758
rect 2218 1974 2378 2730
rect 4214 2730 4242 5278
rect 5054 4970 5082 4975
rect 5054 3794 5082 4942
rect 5054 3761 5082 3766
rect 10486 3402 10514 5614
rect 11662 5530 11690 5726
rect 11662 5497 11690 5502
rect 11888 5502 12048 6258
rect 11888 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12048 5502
rect 11438 5362 11466 5367
rect 11438 5138 11466 5334
rect 11438 5105 11466 5110
rect 10486 3369 10514 3374
rect 11888 4718 12048 5474
rect 12218 6678 12378 7112
rect 12218 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12378 6678
rect 12218 5894 12378 6650
rect 12218 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12378 5894
rect 12218 5110 12378 5866
rect 12218 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12378 5110
rect 11888 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12048 4718
rect 11888 3934 12048 4690
rect 12110 4858 12138 4863
rect 12110 4578 12138 4830
rect 12110 4545 12138 4550
rect 11888 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12048 3934
rect 4214 2697 4242 2702
rect 11888 3150 12048 3906
rect 11888 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12048 3150
rect 2218 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2378 1974
rect 2218 1190 2378 1946
rect 2218 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2378 1190
rect 2218 406 2378 1162
rect 2218 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2378 406
rect 2218 0 2378 378
rect 11888 2366 12048 3122
rect 11888 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12048 2366
rect 11888 1582 12048 2338
rect 11888 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12048 1582
rect 11888 798 12048 1554
rect 11888 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12048 798
rect 11888 0 12048 770
rect 12218 4326 12378 5082
rect 12218 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12378 4326
rect 12218 3542 12378 4298
rect 12218 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12378 3542
rect 12218 2758 12378 3514
rect 12218 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12378 2758
rect 12218 1974 12378 2730
rect 12218 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12378 1974
rect 12218 1190 12378 1946
rect 12218 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12378 1190
rect 12218 406 12378 1162
rect 12218 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12378 406
rect 12218 0 12378 378
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _00_
timestamp 1486834041
transform 1 0 7056 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _01_
timestamp 1486834041
transform 1 0 7504 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _02_
timestamp 1486834041
transform 1 0 8064 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _03_
timestamp 1486834041
transform 1 0 7728 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _04_
timestamp 1486834041
transform 1 0 6888 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _05_
timestamp 1486834041
transform 1 0 8064 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _06_
timestamp 1486834041
transform 1 0 7616 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _07_
timestamp 1486834041
transform 1 0 6944 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _08_
timestamp 1486834041
transform 1 0 7224 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _09_
timestamp 1486834041
transform 1 0 6720 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _10_
timestamp 1486834041
transform 1 0 7728 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _11_
timestamp 1486834041
transform 1 0 8344 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _12_
timestamp 1486834041
transform 1 0 8288 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _13_
timestamp 1486834041
transform 1 0 7168 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _14_
timestamp 1486834041
transform 1 0 7112 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _15_
timestamp 1486834041
transform 1 0 7280 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _16_
timestamp 1486834041
transform 1 0 7728 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _17_
timestamp 1486834041
transform 1 0 8120 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _18_
timestamp 1486834041
transform 1 0 7560 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _19_
timestamp 1486834041
transform 1 0 8064 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _20_
timestamp 1486834041
transform 1 0 7616 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _21_
timestamp 1486834041
transform 1 0 7504 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _22_
timestamp 1486834041
transform 1 0 7728 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _23_
timestamp 1486834041
transform 1 0 7168 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _24_
timestamp 1486834041
transform 1 0 8792 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _25_
timestamp 1486834041
transform 1 0 7784 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _26_
timestamp 1486834041
transform 1 0 8568 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _27_
timestamp 1486834041
transform 1 0 11424 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _28_
timestamp 1486834041
transform 1 0 9688 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _29_
timestamp 1486834041
transform 1 0 10136 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _30_
timestamp 1486834041
transform 1 0 10640 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _31_
timestamp 1486834041
transform 1 0 14952 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _32_
timestamp 1486834041
transform 1 0 9240 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _33_
timestamp 1486834041
transform 1 0 9744 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _34_
timestamp 1486834041
transform 1 0 10304 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _35_
timestamp 1486834041
transform 1 0 10752 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _36_
timestamp 1486834041
transform 1 0 13384 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _37_
timestamp 1486834041
transform 1 0 1456 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _38_
timestamp 1486834041
transform -1 0 5880 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _39_
timestamp 1486834041
transform -1 0 6664 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _40_
timestamp 1486834041
transform -1 0 7056 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _41_
timestamp 1486834041
transform 1 0 8848 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _42_
timestamp 1486834041
transform 1 0 11256 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _43_
timestamp 1486834041
transform 1 0 11312 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _44_
timestamp 1486834041
transform 1 0 10472 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _45_
timestamp 1486834041
transform 1 0 11704 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _46_
timestamp 1486834041
transform 1 0 12488 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _47_
timestamp 1486834041
transform -1 0 11480 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _48_
timestamp 1486834041
transform 1 0 12656 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _49_
timestamp 1486834041
transform 1 0 13216 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _50_
timestamp 1486834041
transform 1 0 14168 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _51_
timestamp 1486834041
transform -1 0 14616 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _52_
timestamp 1486834041
transform -1 0 4816 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _53_
timestamp 1486834041
transform -1 0 3808 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _54_
timestamp 1486834041
transform -1 0 2688 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _55_
timestamp 1486834041
transform -1 0 2240 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _56_
timestamp 1486834041
transform -1 0 7560 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _57_
timestamp 1486834041
transform -1 0 7280 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _58_
timestamp 1486834041
transform -1 0 4872 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _59_
timestamp 1486834041
transform -1 0 6328 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _60_
timestamp 1486834041
transform -1 0 6104 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _61_
timestamp 1486834041
transform -1 0 5376 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _62_
timestamp 1486834041
transform -1 0 5544 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _63_
timestamp 1486834041
transform -1 0 5880 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _64_
timestamp 1486834041
transform -1 0 9128 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _65_
timestamp 1486834041
transform -1 0 8680 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _66_
timestamp 1486834041
transform -1 0 8232 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _67_
timestamp 1486834041
transform -1 0 7952 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _68_
timestamp 1486834041
transform -1 0 6664 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _69_
timestamp 1486834041
transform -1 0 7784 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _70_
timestamp 1486834041
transform 1 0 2632 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _71_
timestamp 1486834041
transform -1 0 4256 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _72_
timestamp 1486834041
transform 1 0 14168 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _73_
timestamp 1486834041
transform 1 0 11872 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _74_
timestamp 1486834041
transform 1 0 11480 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _75_
timestamp 1486834041
transform 1 0 11032 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _76_
timestamp 1486834041
transform 1 0 10584 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _77_
timestamp 1486834041
transform 1 0 10472 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _78_
timestamp 1486834041
transform -1 0 10136 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _79_
timestamp 1486834041
transform -1 0 9632 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _80_
timestamp 1486834041
transform -1 0 9184 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _81_
timestamp 1486834041
transform -1 0 9576 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _82_
timestamp 1486834041
transform -1 0 4424 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _83_
timestamp 1486834041
transform 1 0 2632 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _84_
timestamp 1486834041
transform 1 0 9688 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _85_
timestamp 1486834041
transform 1 0 9408 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _86_
timestamp 1486834041
transform -1 0 9240 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _87_
timestamp 1486834041
transform -1 0 6832 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _88_
timestamp 1486834041
transform 1 0 9968 0 1 392
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__00__I
timestamp 1486834041
transform 1 0 6944 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__01__I
timestamp 1486834041
transform -1 0 7504 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__02__I
timestamp 1486834041
transform 1 0 8512 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__03__I
timestamp 1486834041
transform 1 0 7616 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__04__I
timestamp 1486834041
transform 1 0 6776 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__05__I
timestamp 1486834041
transform -1 0 8064 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__06__I
timestamp 1486834041
transform 1 0 7504 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__07__I
timestamp 1486834041
transform 1 0 6832 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__08__I
timestamp 1486834041
transform -1 0 7056 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__09__I
timestamp 1486834041
transform 1 0 6608 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__10__I
timestamp 1486834041
transform 1 0 7616 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__11__I
timestamp 1486834041
transform -1 0 8344 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__12__I
timestamp 1486834041
transform 1 0 8064 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__13__I
timestamp 1486834041
transform -1 0 7168 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__14__I
timestamp 1486834041
transform 1 0 7000 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__15__I
timestamp 1486834041
transform -1 0 7280 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__16__I
timestamp 1486834041
transform 1 0 7616 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__17__I
timestamp 1486834041
transform -1 0 8120 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__18__I
timestamp 1486834041
transform 1 0 7448 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__19__I
timestamp 1486834041
transform 1 0 7952 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__20__I
timestamp 1486834041
transform 1 0 7448 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__21__I
timestamp 1486834041
transform 1 0 7392 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__22__I
timestamp 1486834041
transform -1 0 7728 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__23__I
timestamp 1486834041
transform 1 0 7056 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__24__I
timestamp 1486834041
transform -1 0 8792 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__25__I
timestamp 1486834041
transform 1 0 7672 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__26__I
timestamp 1486834041
transform -1 0 8568 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__27__I
timestamp 1486834041
transform 1 0 11312 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__28__I
timestamp 1486834041
transform -1 0 9688 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__29__I
timestamp 1486834041
transform -1 0 9464 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__30__I
timestamp 1486834041
transform 1 0 11088 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__31__I
timestamp 1486834041
transform 1 0 13944 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__32__I
timestamp 1486834041
transform 1 0 9128 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__33__I
timestamp 1486834041
transform 1 0 9632 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__34__I
timestamp 1486834041
transform 1 0 10192 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__35__I
timestamp 1486834041
transform -1 0 10752 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__36__I
timestamp 1486834041
transform 1 0 13440 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__37__I
timestamp 1486834041
transform -1 0 1456 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__38__I
timestamp 1486834041
transform 1 0 5880 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__39__I
timestamp 1486834041
transform 1 0 6664 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__40__I
timestamp 1486834041
transform 1 0 7056 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__41__I
timestamp 1486834041
transform -1 0 8848 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__42__I
timestamp 1486834041
transform 1 0 11144 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__43__I
timestamp 1486834041
transform -1 0 11144 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__44__I
timestamp 1486834041
transform -1 0 10472 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__45__I
timestamp 1486834041
transform -1 0 11704 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__46__I
timestamp 1486834041
transform 1 0 12376 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__47__I
timestamp 1486834041
transform 1 0 11928 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__48__I
timestamp 1486834041
transform -1 0 12656 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__49__I
timestamp 1486834041
transform 1 0 13664 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__50__I
timestamp 1486834041
transform -1 0 14056 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__51__I
timestamp 1486834041
transform -1 0 14616 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__52__I
timestamp 1486834041
transform -1 0 4928 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__53__I
timestamp 1486834041
transform 1 0 3808 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__54__I
timestamp 1486834041
transform -1 0 2800 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__55__I
timestamp 1486834041
transform 1 0 2408 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__56__I
timestamp 1486834041
transform -1 0 7672 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__57__I
timestamp 1486834041
transform -1 0 7392 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__58__I
timestamp 1486834041
transform -1 0 4648 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__59__I
timestamp 1486834041
transform -1 0 6440 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__60__I
timestamp 1486834041
transform 1 0 6104 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__61__I
timestamp 1486834041
transform -1 0 5656 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__62__I
timestamp 1486834041
transform 1 0 5656 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__63__I
timestamp 1486834041
transform -1 0 5992 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__64__I
timestamp 1486834041
transform 1 0 9128 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__65__I
timestamp 1486834041
transform -1 0 8792 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__66__I
timestamp 1486834041
transform 1 0 8232 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__67__I
timestamp 1486834041
transform -1 0 8176 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__68__I
timestamp 1486834041
transform -1 0 6552 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__69__I
timestamp 1486834041
transform -1 0 8120 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__70__I
timestamp 1486834041
transform -1 0 2632 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__71__I
timestamp 1486834041
transform -1 0 4480 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__72__I
timestamp 1486834041
transform 1 0 13832 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__73__I
timestamp 1486834041
transform -1 0 11872 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__74__I
timestamp 1486834041
transform -1 0 11312 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__75__I
timestamp 1486834041
transform -1 0 11032 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__76__I
timestamp 1486834041
transform -1 0 10360 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__77__I
timestamp 1486834041
transform -1 0 10472 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__78__I
timestamp 1486834041
transform 1 0 10136 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__79__I
timestamp 1486834041
transform -1 0 9744 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__80__I
timestamp 1486834041
transform -1 0 9296 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__81__I
timestamp 1486834041
transform 1 0 9576 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__82__I
timestamp 1486834041
transform 1 0 4424 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__83__I
timestamp 1486834041
transform -1 0 2632 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__84__I
timestamp 1486834041
transform -1 0 9576 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__85__I
timestamp 1486834041
transform -1 0 8792 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__86__I
timestamp 1486834041
transform 1 0 9240 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__87__I
timestamp 1486834041
transform -1 0 6944 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__88__I
timestamp 1486834041
transform -1 0 9856 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2
timestamp 1486834041
transform 1 0 448 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36
timestamp 1486834041
transform 1 0 2352 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70
timestamp 1486834041
transform 1 0 4256 0 1 392
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86
timestamp 1486834041
transform 1 0 5152 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90
timestamp 1486834041
transform 1 0 5376 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101
timestamp 1486834041
transform 1 0 5992 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1486834041
transform 1 0 6160 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115
timestamp 1486834041
transform 1 0 6776 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_117
timestamp 1486834041
transform 1 0 6888 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_122
timestamp 1486834041
transform 1 0 7168 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_148
timestamp 1486834041
transform 1 0 8624 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_160
timestamp 1486834041
transform 1 0 9296 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_164
timestamp 1486834041
transform 1 0 9520 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_178
timestamp 1486834041
transform 1 0 10304 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_189
timestamp 1486834041
transform 1 0 10920 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195
timestamp 1486834041
transform 1 0 11256 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_206
timestamp 1486834041
transform 1 0 11872 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_240
timestamp 1486834041
transform 1 0 13776 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2
timestamp 1486834041
transform 1 0 448 0 -1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1486834041
transform 1 0 4032 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_72
timestamp 1486834041
transform 1 0 4368 0 -1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_104
timestamp 1486834041
transform 1 0 6160 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_128
timestamp 1486834041
transform 1 0 7504 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_142
timestamp 1486834041
transform 1 0 8288 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_144
timestamp 1486834041
transform 1 0 8400 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_147
timestamp 1486834041
transform 1 0 8568 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_155
timestamp 1486834041
transform 1 0 9016 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_167
timestamp 1486834041
transform 1 0 9688 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_194
timestamp 1486834041
transform 1 0 11200 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_203
timestamp 1486834041
transform 1 0 11704 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_207
timestamp 1486834041
transform 1 0 11928 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_209
timestamp 1486834041
transform 1 0 12040 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_212
timestamp 1486834041
transform 1 0 12208 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_214
timestamp 1486834041
transform 1 0 12320 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_225
timestamp 1486834041
transform 1 0 12936 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1486834041
transform 1 0 448 0 1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1486834041
transform 1 0 2240 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1486834041
transform 1 0 2408 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1486834041
transform 1 0 5992 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_107
timestamp 1486834041
transform 1 0 6328 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_115
timestamp 1486834041
transform 1 0 6776 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_126
timestamp 1486834041
transform 1 0 7392 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_146
timestamp 1486834041
transform 1 0 8512 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_155
timestamp 1486834041
transform 1 0 9016 0 1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 9912 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_177
timestamp 1486834041
transform 1 0 10248 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_181
timestamp 1486834041
transform 1 0 10472 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_183
timestamp 1486834041
transform 1 0 10584 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_186
timestamp 1486834041
transform 1 0 10752 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_194
timestamp 1486834041
transform 1 0 11200 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_198
timestamp 1486834041
transform 1 0 11424 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_200
timestamp 1486834041
transform 1 0 11536 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_211
timestamp 1486834041
transform 1 0 12152 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_215
timestamp 1486834041
transform 1 0 12376 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_217
timestamp 1486834041
transform 1 0 12488 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_228
timestamp 1486834041
transform 1 0 13104 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_230
timestamp 1486834041
transform 1 0 13216 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1486834041
transform 1 0 448 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1486834041
transform 1 0 4032 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_72
timestamp 1486834041
transform 1 0 4368 0 -1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_104
timestamp 1486834041
transform 1 0 6160 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_112
timestamp 1486834041
transform 1 0 6608 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_114
timestamp 1486834041
transform 1 0 6720 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_125
timestamp 1486834041
transform 1 0 7336 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_133
timestamp 1486834041
transform 1 0 7784 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_135
timestamp 1486834041
transform 1 0 7896 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_138
timestamp 1486834041
transform 1 0 8064 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_142
timestamp 1486834041
transform 1 0 8288 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_206
timestamp 1486834041
transform 1 0 11872 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_212
timestamp 1486834041
transform 1 0 12208 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_228
timestamp 1486834041
transform 1 0 13104 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_240
timestamp 1486834041
transform 1 0 13776 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1486834041
transform 1 0 448 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 2240 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1486834041
transform 1 0 2408 0 1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1486834041
transform 1 0 5992 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_107
timestamp 1486834041
transform 1 0 6328 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_115
timestamp 1486834041
transform 1 0 6776 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_117
timestamp 1486834041
transform 1 0 6888 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_122
timestamp 1486834041
transform 1 0 7168 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_143
timestamp 1486834041
transform 1 0 8344 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_147
timestamp 1486834041
transform 1 0 8568 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_151
timestamp 1486834041
transform 1 0 8792 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_167
timestamp 1486834041
transform 1 0 9688 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_177
timestamp 1486834041
transform 1 0 10248 0 1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_241
timestamp 1486834041
transform 1 0 13832 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_247
timestamp 1486834041
transform 1 0 14168 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_251
timestamp 1486834041
transform 1 0 14392 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1486834041
transform 1 0 448 0 -1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1486834041
transform 1 0 4032 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_72
timestamp 1486834041
transform 1 0 4368 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_104
timestamp 1486834041
transform 1 0 6160 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_142
timestamp 1486834041
transform 1 0 8288 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_159
timestamp 1486834041
transform 1 0 9240 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_191
timestamp 1486834041
transform 1 0 11032 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_207
timestamp 1486834041
transform 1 0 11928 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_209
timestamp 1486834041
transform 1 0 12040 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_212
timestamp 1486834041
transform 1 0 12208 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_228
timestamp 1486834041
transform 1 0 13104 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_236
timestamp 1486834041
transform 1 0 13552 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_240
timestamp 1486834041
transform 1 0 13776 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1486834041
transform 1 0 448 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 2240 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1486834041
transform 1 0 2408 0 1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1486834041
transform 1 0 5992 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_107
timestamp 1486834041
transform 1 0 6328 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_115
timestamp 1486834041
transform 1 0 6776 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_119
timestamp 1486834041
transform 1 0 7000 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_130
timestamp 1486834041
transform 1 0 7616 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_162
timestamp 1486834041
transform 1 0 9408 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_170
timestamp 1486834041
transform 1 0 9856 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_174
timestamp 1486834041
transform 1 0 10080 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_177
timestamp 1486834041
transform 1 0 10248 0 1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_241
timestamp 1486834041
transform 1 0 13832 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_247
timestamp 1486834041
transform 1 0 14168 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_2
timestamp 1486834041
transform 1 0 448 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_34
timestamp 1486834041
transform 1 0 2240 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_50
timestamp 1486834041
transform 1 0 3136 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_58
timestamp 1486834041
transform 1 0 3584 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_74
timestamp 1486834041
transform 1 0 4480 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_106
timestamp 1486834041
transform 1 0 6272 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_114
timestamp 1486834041
transform 1 0 6720 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_118
timestamp 1486834041
transform 1 0 6944 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_129
timestamp 1486834041
transform 1 0 7560 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_132
timestamp 1486834041
transform 1 0 7728 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_136
timestamp 1486834041
transform 1 0 7952 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_150
timestamp 1486834041
transform 1 0 8736 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_182
timestamp 1486834041
transform 1 0 10528 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_198
timestamp 1486834041
transform 1 0 11424 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_206
timestamp 1486834041
transform 1 0 11872 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_212
timestamp 1486834041
transform 1 0 12208 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_220
timestamp 1486834041
transform 1 0 12656 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_224
timestamp 1486834041
transform 1 0 12880 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_226
timestamp 1486834041
transform 1 0 12992 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1486834041
transform 1 0 448 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 2240 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_37
timestamp 1486834041
transform 1 0 2408 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_41
timestamp 1486834041
transform 1 0 2632 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_44
timestamp 1486834041
transform 1 0 2800 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_52
timestamp 1486834041
transform 1 0 3248 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_64
timestamp 1486834041
transform 1 0 3920 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_75
timestamp 1486834041
transform 1 0 4536 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_83
timestamp 1486834041
transform 1 0 4984 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_97
timestamp 1486834041
transform 1 0 5768 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1486834041
transform 1 0 5992 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_107
timestamp 1486834041
transform 1 0 6328 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_115
timestamp 1486834041
transform 1 0 6776 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_119
timestamp 1486834041
transform 1 0 7000 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_121
timestamp 1486834041
transform 1 0 7112 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_140
timestamp 1486834041
transform 1 0 8176 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_172
timestamp 1486834041
transform 1 0 9968 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_174
timestamp 1486834041
transform 1 0 10080 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_177
timestamp 1486834041
transform 1 0 10248 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_209
timestamp 1486834041
transform 1 0 12040 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_247
timestamp 1486834041
transform 1 0 14168 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_2
timestamp 1486834041
transform 1 0 448 0 -1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_90
timestamp 1486834041
transform 1 0 5376 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_109
timestamp 1486834041
transform 1 0 6440 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_125
timestamp 1486834041
transform 1 0 7336 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_129
timestamp 1486834041
transform 1 0 7560 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_142
timestamp 1486834041
transform 1 0 8288 0 -1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_174
timestamp 1486834041
transform 1 0 10080 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_190
timestamp 1486834041
transform 1 0 10976 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_198
timestamp 1486834041
transform 1 0 11424 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_202
timestamp 1486834041
transform 1 0 11648 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_206
timestamp 1486834041
transform 1 0 11872 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1486834041
transform 1 0 12208 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_2
timestamp 1486834041
transform 1 0 448 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_18
timestamp 1486834041
transform 1 0 1344 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1486834041
transform 1 0 2240 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_107
timestamp 1486834041
transform 1 0 6328 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_115
timestamp 1486834041
transform 1 0 6776 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_118
timestamp 1486834041
transform 1 0 6944 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_136
timestamp 1486834041
transform 1 0 7952 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_147
timestamp 1486834041
transform 1 0 8568 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_163
timestamp 1486834041
transform 1 0 9464 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_171
timestamp 1486834041
transform 1 0 9912 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_177
timestamp 1486834041
transform 1 0 10248 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_193
timestamp 1486834041
transform 1 0 11144 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_214
timestamp 1486834041
transform 1 0 12320 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_216
timestamp 1486834041
transform 1 0 12432 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_2
timestamp 1486834041
transform 1 0 448 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_18
timestamp 1486834041
transform 1 0 1344 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_26
timestamp 1486834041
transform 1 0 1792 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_72
timestamp 1486834041
transform 1 0 4368 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_74
timestamp 1486834041
transform 1 0 4480 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_105
timestamp 1486834041
transform 1 0 6216 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_107
timestamp 1486834041
transform 1 0 6328 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_126
timestamp 1486834041
transform 1 0 7392 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_131
timestamp 1486834041
transform 1 0 7672 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_135
timestamp 1486834041
transform 1 0 7896 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_138
timestamp 1486834041
transform 1 0 8064 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_142
timestamp 1486834041
transform 1 0 8288 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_160
timestamp 1486834041
transform 1 0 9296 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_164
timestamp 1486834041
transform 1 0 9520 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_168
timestamp 1486834041
transform 1 0 9744 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_172
timestamp 1486834041
transform 1 0 9968 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_174
timestamp 1486834041
transform 1 0 10080 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_209
timestamp 1486834041
transform 1 0 12040 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_240
timestamp 1486834041
transform 1 0 13776 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_2
timestamp 1486834041
transform 1 0 448 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_18
timestamp 1486834041
transform 1 0 1344 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_20
timestamp 1486834041
transform 1 0 1456 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_37
timestamp 1486834041
transform 1 0 2408 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_129
timestamp 1486834041
transform 1 0 7560 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_146
timestamp 1486834041
transform 1 0 8512 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_166
timestamp 1486834041
transform 1 0 9632 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_2
timestamp 1486834041
transform 1 0 448 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_72
timestamp 1486834041
transform 1 0 4368 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_123
timestamp 1486834041
transform 1 0 7224 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_139
timestamp 1486834041
transform 1 0 8120 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_142
timestamp 1486834041
transform 1 0 8288 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_146
timestamp 1486834041
transform 1 0 8512 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_148
timestamp 1486834041
transform 1 0 8624 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_151
timestamp 1486834041
transform 1 0 8792 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_155
timestamp 1486834041
transform 1 0 9016 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_159
timestamp 1486834041
transform 1 0 9240 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_183
timestamp 1486834041
transform 1 0 10584 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_194
timestamp 1486834041
transform 1 0 11200 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_209
timestamp 1486834041
transform 1 0 12040 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_254
timestamp 1486834041
transform 1 0 14560 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_2
timestamp 1486834041
transform 1 0 448 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_18
timestamp 1486834041
transform 1 0 1344 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_20
timestamp 1486834041
transform 1 0 1456 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_37
timestamp 1486834041
transform 1 0 2408 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_107
timestamp 1486834041
transform 1 0 6328 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_241
timestamp 1486834041
transform 1 0 13832 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_2
timestamp 1486834041
transform 1 0 448 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_36
timestamp 1486834041
transform 1 0 2352 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_70
timestamp 1486834041
transform 1 0 4256 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_104
timestamp 1486834041
transform 1 0 6160 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_127
timestamp 1486834041
transform 1 0 7448 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_140
timestamp 1486834041
transform 1 0 8176 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_143
timestamp 1486834041
transform 1 0 8344 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_147
timestamp 1486834041
transform 1 0 8568 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_161
timestamp 1486834041
transform 1 0 9352 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_172
timestamp 1486834041
transform 1 0 9968 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_174
timestamp 1486834041
transform 1 0 10080 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_203
timestamp 1486834041
transform 1 0 11704 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_236
timestamp 1486834041
transform 1 0 13552 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_268
timestamp 1486834041
transform 1 0 15344 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform 1 0 13272 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform 1 0 14616 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform 1 0 13832 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform 1 0 14616 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform 1 0 14616 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform 1 0 13832 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform 1 0 14616 0 1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform 1 0 14616 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform 1 0 14616 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform 1 0 14616 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform 1 0 14616 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform 1 0 12096 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform 1 0 14616 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform 1 0 14616 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 14616 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 13832 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform 1 0 13832 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 13048 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform 1 0 13272 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform -1 0 10920 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform 1 0 12264 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform 1 0 13048 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 12880 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform -1 0 11032 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform -1 0 13272 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 13048 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 13832 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 13832 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 14616 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 14616 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform 1 0 13832 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 14616 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform 1 0 10920 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform 1 0 12992 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform 1 0 12208 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform 1 0 13776 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform 1 0 13048 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform -1 0 13272 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform 1 0 13776 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform 1 0 14168 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform -1 0 13776 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform 1 0 14560 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform -1 0 14056 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform 1 0 11032 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform 1 0 11872 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform 1 0 11256 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform -1 0 12600 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform 1 0 11480 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform 1 0 12656 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform 1 0 12600 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform 1 0 12208 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform 1 0 12264 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform -1 0 2296 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform -1 0 3472 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform 1 0 1904 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform 1 0 2520 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform -1 0 1456 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform -1 0 2688 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform -1 0 2296 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform -1 0 3472 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform -1 0 4256 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform -1 0 4088 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform -1 0 2240 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform -1 0 3472 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform -1 0 3864 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform -1 0 4256 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform -1 0 4872 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform -1 0 3360 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform -1 0 4256 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform -1 0 4648 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform 1 0 3080 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform 1 0 4872 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform -1 0 5432 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform 1 0 5656 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform 1 0 5432 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform -1 0 6048 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform -1 0 7224 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform -1 0 7336 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform 1 0 6664 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform -1 0 4144 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform -1 0 4648 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform -1 0 5432 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform -1 0 6216 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform -1 0 5656 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform -1 0 5432 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform -1 0 6216 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform -1 0 5264 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform -1 0 7112 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output89
timestamp 1486834041
transform 1 0 10248 0 1 5096
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_16
timestamp 1486834041
transform 1 0 336 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 15512 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_17
timestamp 1486834041
transform 1 0 336 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 15512 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_18
timestamp 1486834041
transform 1 0 336 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 15512 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_19
timestamp 1486834041
transform 1 0 336 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 15512 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_20
timestamp 1486834041
transform 1 0 336 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 15512 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_21
timestamp 1486834041
transform 1 0 336 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 15512 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_22
timestamp 1486834041
transform 1 0 336 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 15512 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_23
timestamp 1486834041
transform 1 0 336 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 15512 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_24
timestamp 1486834041
transform 1 0 336 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 15512 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_25
timestamp 1486834041
transform 1 0 336 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 15512 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_26
timestamp 1486834041
transform 1 0 336 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 15512 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_27
timestamp 1486834041
transform 1 0 336 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 15512 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_28
timestamp 1486834041
transform 1 0 336 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 15512 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_29
timestamp 1486834041
transform 1 0 336 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 15512 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_30
timestamp 1486834041
transform 1 0 336 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 15512 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_31
timestamp 1486834041
transform 1 0 336 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 15512 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_32
timestamp 1486834041
transform 1 0 2240 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_33
timestamp 1486834041
transform 1 0 4144 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34
timestamp 1486834041
transform 1 0 6048 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1486834041
transform 1 0 7952 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1486834041
transform 1 0 9856 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1486834041
transform 1 0 11760 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1486834041
transform 1 0 13664 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_39
timestamp 1486834041
transform 1 0 4256 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_40
timestamp 1486834041
transform 1 0 8176 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_41
timestamp 1486834041
transform 1 0 12096 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_42
timestamp 1486834041
transform 1 0 2296 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_43
timestamp 1486834041
transform 1 0 6216 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_44
timestamp 1486834041
transform 1 0 10136 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_45
timestamp 1486834041
transform 1 0 14056 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_46
timestamp 1486834041
transform 1 0 4256 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_47
timestamp 1486834041
transform 1 0 8176 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_48
timestamp 1486834041
transform 1 0 12096 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_49
timestamp 1486834041
transform 1 0 2296 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_50
timestamp 1486834041
transform 1 0 6216 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_51
timestamp 1486834041
transform 1 0 10136 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_52
timestamp 1486834041
transform 1 0 14056 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_53
timestamp 1486834041
transform 1 0 4256 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_54
timestamp 1486834041
transform 1 0 8176 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_55
timestamp 1486834041
transform 1 0 12096 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_56
timestamp 1486834041
transform 1 0 2296 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_57
timestamp 1486834041
transform 1 0 6216 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_58
timestamp 1486834041
transform 1 0 10136 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_59
timestamp 1486834041
transform 1 0 14056 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_60
timestamp 1486834041
transform 1 0 4256 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_61
timestamp 1486834041
transform 1 0 8176 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_62
timestamp 1486834041
transform 1 0 12096 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_63
timestamp 1486834041
transform 1 0 2296 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_64
timestamp 1486834041
transform 1 0 6216 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_65
timestamp 1486834041
transform 1 0 10136 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_66
timestamp 1486834041
transform 1 0 14056 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_67
timestamp 1486834041
transform 1 0 4256 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_68
timestamp 1486834041
transform 1 0 8176 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_69
timestamp 1486834041
transform 1 0 12096 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_70
timestamp 1486834041
transform 1 0 2296 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_71
timestamp 1486834041
transform 1 0 6216 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_72
timestamp 1486834041
transform 1 0 10136 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_73
timestamp 1486834041
transform 1 0 14056 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_74
timestamp 1486834041
transform 1 0 4256 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_75
timestamp 1486834041
transform 1 0 8176 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_76
timestamp 1486834041
transform 1 0 12096 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_77
timestamp 1486834041
transform 1 0 2296 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_78
timestamp 1486834041
transform 1 0 6216 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_79
timestamp 1486834041
transform 1 0 10136 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_80
timestamp 1486834041
transform 1 0 14056 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_81
timestamp 1486834041
transform 1 0 4256 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_82
timestamp 1486834041
transform 1 0 8176 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_83
timestamp 1486834041
transform 1 0 12096 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_84
timestamp 1486834041
transform 1 0 2296 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_85
timestamp 1486834041
transform 1 0 6216 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_86
timestamp 1486834041
transform 1 0 10136 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_87
timestamp 1486834041
transform 1 0 14056 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_88
timestamp 1486834041
transform 1 0 2240 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_89
timestamp 1486834041
transform 1 0 4144 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_90
timestamp 1486834041
transform 1 0 6048 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_91
timestamp 1486834041
transform 1 0 7952 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_92
timestamp 1486834041
transform 1 0 9856 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_93
timestamp 1486834041
transform 1 0 11760 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_94
timestamp 1486834041
transform 1 0 13664 0 -1 6664
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 0 56 56 0 FreeSans 224 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 2240 56 2296 0 FreeSans 224 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 2464 56 2520 0 FreeSans 224 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 2688 56 2744 0 FreeSans 224 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 2912 56 2968 0 FreeSans 224 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 3136 56 3192 0 FreeSans 224 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 3360 56 3416 0 FreeSans 224 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 3584 56 3640 0 FreeSans 224 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 3808 56 3864 0 FreeSans 224 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 4032 56 4088 0 FreeSans 224 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 4256 56 4312 0 FreeSans 224 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 224 56 280 0 FreeSans 224 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 4480 56 4536 0 FreeSans 224 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 4704 56 4760 0 FreeSans 224 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 4928 56 4984 0 FreeSans 224 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 5152 56 5208 0 FreeSans 224 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 5376 56 5432 0 FreeSans 224 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 5600 56 5656 0 FreeSans 224 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 5824 56 5880 0 FreeSans 224 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 6048 56 6104 0 FreeSans 224 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 6272 56 6328 0 FreeSans 224 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 6496 56 6552 0 FreeSans 224 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 448 56 504 0 FreeSans 224 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 6720 56 6776 0 FreeSans 224 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 6944 56 7000 0 FreeSans 224 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 672 56 728 0 FreeSans 224 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 896 56 952 0 FreeSans 224 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 1120 56 1176 0 FreeSans 224 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 1344 56 1400 0 FreeSans 224 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 1568 56 1624 0 FreeSans 224 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 1792 56 1848 0 FreeSans 224 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 2016 56 2072 0 FreeSans 224 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 15792 0 15848 56 0 FreeSans 224 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 15792 2240 15848 2296 0 FreeSans 224 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 15792 2464 15848 2520 0 FreeSans 224 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 15792 2688 15848 2744 0 FreeSans 224 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 15792 2912 15848 2968 0 FreeSans 224 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 15792 3136 15848 3192 0 FreeSans 224 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 15792 3360 15848 3416 0 FreeSans 224 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 15792 3584 15848 3640 0 FreeSans 224 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 15792 3808 15848 3864 0 FreeSans 224 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 15792 4032 15848 4088 0 FreeSans 224 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 15792 4256 15848 4312 0 FreeSans 224 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 15792 224 15848 280 0 FreeSans 224 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 15792 4480 15848 4536 0 FreeSans 224 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 15792 4704 15848 4760 0 FreeSans 224 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 15792 4928 15848 4984 0 FreeSans 224 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 15792 5152 15848 5208 0 FreeSans 224 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 15792 5376 15848 5432 0 FreeSans 224 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 15792 5600 15848 5656 0 FreeSans 224 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 15792 5824 15848 5880 0 FreeSans 224 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 15792 6048 15848 6104 0 FreeSans 224 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 15792 6272 15848 6328 0 FreeSans 224 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 15792 6496 15848 6552 0 FreeSans 224 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 15792 448 15848 504 0 FreeSans 224 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 15792 6720 15848 6776 0 FreeSans 224 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 15792 6944 15848 7000 0 FreeSans 224 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 15792 672 15848 728 0 FreeSans 224 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 15792 896 15848 952 0 FreeSans 224 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 15792 1120 15848 1176 0 FreeSans 224 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 15792 1344 15848 1400 0 FreeSans 224 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 15792 1568 15848 1624 0 FreeSans 224 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 15792 1792 15848 1848 0 FreeSans 224 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 15792 2016 15848 2072 0 FreeSans 224 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 1792 0 1848 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 8512 0 8568 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 9184 0 9240 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 9856 0 9912 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 10528 0 10584 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 11200 0 11256 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 11872 0 11928 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 12544 0 12600 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 13216 0 13272 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 13888 0 13944 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 14560 0 14616 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 2464 0 2520 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 3136 0 3192 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 3808 0 3864 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 4480 0 4536 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 5152 0 5208 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 5824 0 5880 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 6496 0 6552 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 7168 0 7224 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 7840 0 7896 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 10864 7056 10920 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 11984 7056 12040 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 12096 7056 12152 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 12208 7056 12264 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 12320 7056 12376 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 12432 7056 12488 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 12544 7056 12600 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 12656 7056 12712 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 12768 7056 12824 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 12880 7056 12936 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 12992 7056 13048 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 10976 7056 11032 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 11088 7056 11144 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 11200 7056 11256 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 11312 7056 11368 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 11424 7056 11480 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 11536 7056 11592 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 11648 7056 11704 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 11760 7056 11816 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 11872 7056 11928 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 2688 7056 2744 7112 0 FreeSans 224 0 0 0 N1BEG[0]
port 104 nsew signal output
flabel metal2 s 2800 7056 2856 7112 0 FreeSans 224 0 0 0 N1BEG[1]
port 105 nsew signal output
flabel metal2 s 2912 7056 2968 7112 0 FreeSans 224 0 0 0 N1BEG[2]
port 106 nsew signal output
flabel metal2 s 3024 7056 3080 7112 0 FreeSans 224 0 0 0 N1BEG[3]
port 107 nsew signal output
flabel metal2 s 3136 7056 3192 7112 0 FreeSans 224 0 0 0 N2BEG[0]
port 108 nsew signal output
flabel metal2 s 3248 7056 3304 7112 0 FreeSans 224 0 0 0 N2BEG[1]
port 109 nsew signal output
flabel metal2 s 3360 7056 3416 7112 0 FreeSans 224 0 0 0 N2BEG[2]
port 110 nsew signal output
flabel metal2 s 3472 7056 3528 7112 0 FreeSans 224 0 0 0 N2BEG[3]
port 111 nsew signal output
flabel metal2 s 3584 7056 3640 7112 0 FreeSans 224 0 0 0 N2BEG[4]
port 112 nsew signal output
flabel metal2 s 3696 7056 3752 7112 0 FreeSans 224 0 0 0 N2BEG[5]
port 113 nsew signal output
flabel metal2 s 3808 7056 3864 7112 0 FreeSans 224 0 0 0 N2BEG[6]
port 114 nsew signal output
flabel metal2 s 3920 7056 3976 7112 0 FreeSans 224 0 0 0 N2BEG[7]
port 115 nsew signal output
flabel metal2 s 4032 7056 4088 7112 0 FreeSans 224 0 0 0 N2BEGb[0]
port 116 nsew signal output
flabel metal2 s 4144 7056 4200 7112 0 FreeSans 224 0 0 0 N2BEGb[1]
port 117 nsew signal output
flabel metal2 s 4256 7056 4312 7112 0 FreeSans 224 0 0 0 N2BEGb[2]
port 118 nsew signal output
flabel metal2 s 4368 7056 4424 7112 0 FreeSans 224 0 0 0 N2BEGb[3]
port 119 nsew signal output
flabel metal2 s 4480 7056 4536 7112 0 FreeSans 224 0 0 0 N2BEGb[4]
port 120 nsew signal output
flabel metal2 s 4592 7056 4648 7112 0 FreeSans 224 0 0 0 N2BEGb[5]
port 121 nsew signal output
flabel metal2 s 4704 7056 4760 7112 0 FreeSans 224 0 0 0 N2BEGb[6]
port 122 nsew signal output
flabel metal2 s 4816 7056 4872 7112 0 FreeSans 224 0 0 0 N2BEGb[7]
port 123 nsew signal output
flabel metal2 s 4928 7056 4984 7112 0 FreeSans 224 0 0 0 N4BEG[0]
port 124 nsew signal output
flabel metal2 s 6048 7056 6104 7112 0 FreeSans 224 0 0 0 N4BEG[10]
port 125 nsew signal output
flabel metal2 s 6160 7056 6216 7112 0 FreeSans 224 0 0 0 N4BEG[11]
port 126 nsew signal output
flabel metal2 s 6272 7056 6328 7112 0 FreeSans 224 0 0 0 N4BEG[12]
port 127 nsew signal output
flabel metal2 s 6384 7056 6440 7112 0 FreeSans 224 0 0 0 N4BEG[13]
port 128 nsew signal output
flabel metal2 s 6496 7056 6552 7112 0 FreeSans 224 0 0 0 N4BEG[14]
port 129 nsew signal output
flabel metal2 s 6608 7056 6664 7112 0 FreeSans 224 0 0 0 N4BEG[15]
port 130 nsew signal output
flabel metal2 s 5040 7056 5096 7112 0 FreeSans 224 0 0 0 N4BEG[1]
port 131 nsew signal output
flabel metal2 s 5152 7056 5208 7112 0 FreeSans 224 0 0 0 N4BEG[2]
port 132 nsew signal output
flabel metal2 s 5264 7056 5320 7112 0 FreeSans 224 0 0 0 N4BEG[3]
port 133 nsew signal output
flabel metal2 s 5376 7056 5432 7112 0 FreeSans 224 0 0 0 N4BEG[4]
port 134 nsew signal output
flabel metal2 s 5488 7056 5544 7112 0 FreeSans 224 0 0 0 N4BEG[5]
port 135 nsew signal output
flabel metal2 s 5600 7056 5656 7112 0 FreeSans 224 0 0 0 N4BEG[6]
port 136 nsew signal output
flabel metal2 s 5712 7056 5768 7112 0 FreeSans 224 0 0 0 N4BEG[7]
port 137 nsew signal output
flabel metal2 s 5824 7056 5880 7112 0 FreeSans 224 0 0 0 N4BEG[8]
port 138 nsew signal output
flabel metal2 s 5936 7056 5992 7112 0 FreeSans 224 0 0 0 N4BEG[9]
port 139 nsew signal output
flabel metal2 s 6720 7056 6776 7112 0 FreeSans 224 0 0 0 S1END[0]
port 140 nsew signal input
flabel metal2 s 6832 7056 6888 7112 0 FreeSans 224 0 0 0 S1END[1]
port 141 nsew signal input
flabel metal2 s 6944 7056 7000 7112 0 FreeSans 224 0 0 0 S1END[2]
port 142 nsew signal input
flabel metal2 s 7056 7056 7112 7112 0 FreeSans 224 0 0 0 S1END[3]
port 143 nsew signal input
flabel metal2 s 8064 7056 8120 7112 0 FreeSans 224 0 0 0 S2END[0]
port 144 nsew signal input
flabel metal2 s 8176 7056 8232 7112 0 FreeSans 224 0 0 0 S2END[1]
port 145 nsew signal input
flabel metal2 s 8288 7056 8344 7112 0 FreeSans 224 0 0 0 S2END[2]
port 146 nsew signal input
flabel metal2 s 8400 7056 8456 7112 0 FreeSans 224 0 0 0 S2END[3]
port 147 nsew signal input
flabel metal2 s 8512 7056 8568 7112 0 FreeSans 224 0 0 0 S2END[4]
port 148 nsew signal input
flabel metal2 s 8624 7056 8680 7112 0 FreeSans 224 0 0 0 S2END[5]
port 149 nsew signal input
flabel metal2 s 8736 7056 8792 7112 0 FreeSans 224 0 0 0 S2END[6]
port 150 nsew signal input
flabel metal2 s 8848 7056 8904 7112 0 FreeSans 224 0 0 0 S2END[7]
port 151 nsew signal input
flabel metal2 s 7168 7056 7224 7112 0 FreeSans 224 0 0 0 S2MID[0]
port 152 nsew signal input
flabel metal2 s 7280 7056 7336 7112 0 FreeSans 224 0 0 0 S2MID[1]
port 153 nsew signal input
flabel metal2 s 7392 7056 7448 7112 0 FreeSans 224 0 0 0 S2MID[2]
port 154 nsew signal input
flabel metal2 s 7504 7056 7560 7112 0 FreeSans 224 0 0 0 S2MID[3]
port 155 nsew signal input
flabel metal2 s 7616 7056 7672 7112 0 FreeSans 224 0 0 0 S2MID[4]
port 156 nsew signal input
flabel metal2 s 7728 7056 7784 7112 0 FreeSans 224 0 0 0 S2MID[5]
port 157 nsew signal input
flabel metal2 s 7840 7056 7896 7112 0 FreeSans 224 0 0 0 S2MID[6]
port 158 nsew signal input
flabel metal2 s 7952 7056 8008 7112 0 FreeSans 224 0 0 0 S2MID[7]
port 159 nsew signal input
flabel metal2 s 8960 7056 9016 7112 0 FreeSans 224 0 0 0 S4END[0]
port 160 nsew signal input
flabel metal2 s 10080 7056 10136 7112 0 FreeSans 224 0 0 0 S4END[10]
port 161 nsew signal input
flabel metal2 s 10192 7056 10248 7112 0 FreeSans 224 0 0 0 S4END[11]
port 162 nsew signal input
flabel metal2 s 10304 7056 10360 7112 0 FreeSans 224 0 0 0 S4END[12]
port 163 nsew signal input
flabel metal2 s 10416 7056 10472 7112 0 FreeSans 224 0 0 0 S4END[13]
port 164 nsew signal input
flabel metal2 s 10528 7056 10584 7112 0 FreeSans 224 0 0 0 S4END[14]
port 165 nsew signal input
flabel metal2 s 10640 7056 10696 7112 0 FreeSans 224 0 0 0 S4END[15]
port 166 nsew signal input
flabel metal2 s 9072 7056 9128 7112 0 FreeSans 224 0 0 0 S4END[1]
port 167 nsew signal input
flabel metal2 s 9184 7056 9240 7112 0 FreeSans 224 0 0 0 S4END[2]
port 168 nsew signal input
flabel metal2 s 9296 7056 9352 7112 0 FreeSans 224 0 0 0 S4END[3]
port 169 nsew signal input
flabel metal2 s 9408 7056 9464 7112 0 FreeSans 224 0 0 0 S4END[4]
port 170 nsew signal input
flabel metal2 s 9520 7056 9576 7112 0 FreeSans 224 0 0 0 S4END[5]
port 171 nsew signal input
flabel metal2 s 9632 7056 9688 7112 0 FreeSans 224 0 0 0 S4END[6]
port 172 nsew signal input
flabel metal2 s 9744 7056 9800 7112 0 FreeSans 224 0 0 0 S4END[7]
port 173 nsew signal input
flabel metal2 s 9856 7056 9912 7112 0 FreeSans 224 0 0 0 S4END[8]
port 174 nsew signal input
flabel metal2 s 9968 7056 10024 7112 0 FreeSans 224 0 0 0 S4END[9]
port 175 nsew signal input
flabel metal2 s 1120 0 1176 56 0 FreeSans 224 0 0 0 UserCLK
port 176 nsew signal input
flabel metal2 s 10752 7056 10808 7112 0 FreeSans 224 0 0 0 UserCLKo
port 177 nsew signal output
flabel metal4 s 1888 0 2048 7112 0 FreeSans 736 90 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 1888 0 2048 28 0 FreeSans 184 0 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 1888 7084 2048 7112 0 FreeSans 184 0 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 11888 0 12048 7112 0 FreeSans 736 90 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 11888 0 12048 28 0 FreeSans 184 0 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 11888 7084 12048 7112 0 FreeSans 184 0 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 2218 0 2378 7112 0 FreeSans 736 90 0 0 VSS
port 179 nsew ground bidirectional
flabel metal4 s 2218 0 2378 28 0 FreeSans 184 0 0 0 VSS
port 179 nsew ground bidirectional
flabel metal4 s 2218 7084 2378 7112 0 FreeSans 184 0 0 0 VSS
port 179 nsew ground bidirectional
flabel metal4 s 12218 0 12378 7112 0 FreeSans 736 90 0 0 VSS
port 179 nsew ground bidirectional
flabel metal4 s 12218 0 12378 28 0 FreeSans 184 0 0 0 VSS
port 179 nsew ground bidirectional
flabel metal4 s 12218 7084 12378 7112 0 FreeSans 184 0 0 0 VSS
port 179 nsew ground bidirectional
rlabel metal1 7924 6272 7924 6272 0 VDD
rlabel metal1 7924 6664 7924 6664 0 VSS
rlabel metal3 539 28 539 28 0 FrameData[0]
rlabel metal2 7644 2408 7644 2408 0 FrameData[10]
rlabel metal3 735 2492 735 2492 0 FrameData[11]
rlabel metal3 1071 2716 1071 2716 0 FrameData[12]
rlabel metal2 7224 2660 7224 2660 0 FrameData[13]
rlabel metal3 931 3164 931 3164 0 FrameData[14]
rlabel metal2 7252 3500 7252 3500 0 FrameData[15]
rlabel metal3 1239 3612 1239 3612 0 FrameData[16]
rlabel metal3 1295 3836 1295 3836 0 FrameData[17]
rlabel metal3 1295 4060 1295 4060 0 FrameData[18]
rlabel metal3 1071 4284 1071 4284 0 FrameData[19]
rlabel metal2 7476 364 7476 364 0 FrameData[1]
rlabel metal2 7476 4676 7476 4676 0 FrameData[20]
rlabel metal3 483 4732 483 4732 0 FrameData[21]
rlabel metal3 2555 4956 2555 4956 0 FrameData[22]
rlabel metal3 231 5180 231 5180 0 FrameData[23]
rlabel metal3 1071 5404 1071 5404 0 FrameData[24]
rlabel metal3 2044 3444 2044 3444 0 FrameData[25]
rlabel metal3 567 5852 567 5852 0 FrameData[26]
rlabel metal2 112 2436 112 2436 0 FrameData[27]
rlabel metal3 651 6300 651 6300 0 FrameData[28]
rlabel metal4 5796 6244 5796 6244 0 FrameData[29]
rlabel metal3 2121 476 2121 476 0 FrameData[2]
rlabel metal2 10724 5880 10724 5880 0 FrameData[30]
rlabel metal3 91 6972 91 6972 0 FrameData[31]
rlabel metal2 7644 812 7644 812 0 FrameData[3]
rlabel metal3 1071 924 1071 924 0 FrameData[4]
rlabel metal3 1071 1148 1071 1148 0 FrameData[5]
rlabel metal3 7616 1372 7616 1372 0 FrameData[6]
rlabel metal3 931 1596 931 1596 0 FrameData[7]
rlabel metal2 7028 1932 7028 1932 0 FrameData[8]
rlabel metal2 6636 2296 6636 2296 0 FrameData[9]
rlabel metal3 14777 28 14777 28 0 FrameData_O[0]
rlabel metal2 15204 1988 15204 1988 0 FrameData_O[10]
rlabel metal3 15113 2492 15113 2492 0 FrameData_O[11]
rlabel metal2 15148 2464 15148 2464 0 FrameData_O[12]
rlabel metal2 15092 2772 15092 2772 0 FrameData_O[13]
rlabel metal3 15113 3164 15113 3164 0 FrameData_O[14]
rlabel metal2 15148 3192 15148 3192 0 FrameData_O[15]
rlabel metal2 15204 3444 15204 3444 0 FrameData_O[16]
rlabel metal3 15505 3836 15505 3836 0 FrameData_O[17]
rlabel metal2 15148 3920 15148 3920 0 FrameData_O[18]
rlabel metal3 15449 4284 15449 4284 0 FrameData_O[19]
rlabel metal3 14133 252 14133 252 0 FrameData_O[1]
rlabel metal3 15505 4508 15505 4508 0 FrameData_O[20]
rlabel metal3 15449 4732 15449 4732 0 FrameData_O[21]
rlabel metal3 15505 4956 15505 4956 0 FrameData_O[22]
rlabel metal2 14308 5068 14308 5068 0 FrameData_O[23]
rlabel metal3 15113 5404 15113 5404 0 FrameData_O[24]
rlabel metal3 14721 5628 14721 5628 0 FrameData_O[25]
rlabel metal3 14749 5852 14749 5852 0 FrameData_O[26]
rlabel metal2 10500 6244 10500 6244 0 FrameData_O[27]
rlabel metal2 12740 5236 12740 5236 0 FrameData_O[28]
rlabel metal2 13636 3472 13636 3472 0 FrameData_O[29]
rlabel metal3 14581 476 14581 476 0 FrameData_O[2]
rlabel metal3 15421 6748 15421 6748 0 FrameData_O[30]
rlabel metal2 12852 5376 12852 5376 0 FrameData_O[31]
rlabel metal3 14721 700 14721 700 0 FrameData_O[3]
rlabel metal2 14364 784 14364 784 0 FrameData_O[4]
rlabel metal2 14420 1036 14420 1036 0 FrameData_O[5]
rlabel metal2 15204 1036 15204 1036 0 FrameData_O[6]
rlabel metal2 15092 1316 15092 1316 0 FrameData_O[7]
rlabel metal3 15057 1820 15057 1820 0 FrameData_O[8]
rlabel metal2 15148 1736 15148 1736 0 FrameData_O[9]
rlabel metal2 1820 455 1820 455 0 FrameStrobe[0]
rlabel metal2 11172 420 11172 420 0 FrameStrobe[10]
rlabel metal2 11116 364 11116 364 0 FrameStrobe[11]
rlabel metal2 10444 392 10444 392 0 FrameStrobe[12]
rlabel metal2 11676 1204 11676 1204 0 FrameStrobe[13]
rlabel metal3 11816 924 11816 924 0 FrameStrobe[14]
rlabel metal2 11900 371 11900 371 0 FrameStrobe[15]
rlabel metal2 12628 1064 12628 1064 0 FrameStrobe[16]
rlabel metal2 13244 861 13244 861 0 FrameStrobe[17]
rlabel metal2 13916 63 13916 63 0 FrameStrobe[18]
rlabel metal2 14560 1260 14560 1260 0 FrameStrobe[19]
rlabel metal2 2492 63 2492 63 0 FrameStrobe[1]
rlabel metal2 3164 511 3164 511 0 FrameStrobe[2]
rlabel metal2 3836 455 3836 455 0 FrameStrobe[3]
rlabel metal2 13468 5908 13468 5908 0 FrameStrobe[4]
rlabel metal3 2548 4116 2548 4116 0 FrameStrobe[5]
rlabel metal2 5824 476 5824 476 0 FrameStrobe[6]
rlabel metal2 6524 315 6524 315 0 FrameStrobe[7]
rlabel metal2 7084 812 7084 812 0 FrameStrobe[8]
rlabel metal3 8344 476 8344 476 0 FrameStrobe[9]
rlabel metal2 10892 6825 10892 6825 0 FrameStrobe_O[0]
rlabel metal2 13580 6104 13580 6104 0 FrameStrobe_O[10]
rlabel metal2 12124 6265 12124 6265 0 FrameStrobe_O[11]
rlabel metal2 14140 6692 14140 6692 0 FrameStrobe_O[12]
rlabel metal2 13524 6104 13524 6104 0 FrameStrobe_O[13]
rlabel metal2 12684 5180 12684 5180 0 FrameStrobe_O[14]
rlabel metal2 14140 6076 14140 6076 0 FrameStrobe_O[15]
rlabel metal2 12684 6629 12684 6629 0 FrameStrobe_O[16]
rlabel metal2 12796 6517 12796 6517 0 FrameStrobe_O[17]
rlabel metal2 14924 6664 14924 6664 0 FrameStrobe_O[18]
rlabel metal2 13468 5180 13468 5180 0 FrameStrobe_O[19]
rlabel metal2 11004 6853 11004 6853 0 FrameStrobe_O[1]
rlabel metal2 11116 6797 11116 6797 0 FrameStrobe_O[2]
rlabel metal2 11228 6433 11228 6433 0 FrameStrobe_O[3]
rlabel metal3 11676 6188 11676 6188 0 FrameStrobe_O[4]
rlabel metal2 11452 6237 11452 6237 0 FrameStrobe_O[5]
rlabel metal2 11564 6993 11564 6993 0 FrameStrobe_O[6]
rlabel metal2 11676 6769 11676 6769 0 FrameStrobe_O[7]
rlabel metal2 11788 6349 11788 6349 0 FrameStrobe_O[8]
rlabel metal2 11900 6713 11900 6713 0 FrameStrobe_O[9]
rlabel metal2 2716 6349 2716 6349 0 N1BEG[0]
rlabel metal2 2940 4130 2940 4130 0 N1BEG[1]
rlabel metal2 2436 5264 2436 5264 0 N1BEG[2]
rlabel metal2 2940 5348 2940 5348 0 N1BEG[3]
rlabel metal3 2128 6580 2128 6580 0 N2BEG[0]
rlabel metal2 2324 5768 2324 5768 0 N2BEG[1]
rlabel metal2 3388 6629 3388 6629 0 N2BEG[2]
rlabel metal2 3108 5264 3108 5264 0 N2BEG[3]
rlabel metal2 3836 4130 3836 4130 0 N2BEG[4]
rlabel metal2 3724 5845 3724 5845 0 N2BEG[5]
rlabel metal2 1876 6720 1876 6720 0 N2BEG[6]
rlabel metal2 3108 5824 3108 5824 0 N2BEG[7]
rlabel metal2 4060 6237 4060 6237 0 N2BEGb[0]
rlabel metal2 3892 5152 3892 5152 0 N2BEGb[1]
rlabel metal2 4340 5152 4340 5152 0 N2BEGb[2]
rlabel metal2 2996 6608 2996 6608 0 N2BEGb[3]
rlabel metal2 4508 6713 4508 6713 0 N2BEGb[4]
rlabel metal2 4228 5768 4228 5768 0 N2BEGb[5]
rlabel metal2 3668 6216 3668 6216 0 N2BEGb[6]
rlabel metal2 4844 6181 4844 6181 0 N2BEGb[7]
rlabel metal2 4956 6013 4956 6013 0 N4BEG[0]
rlabel metal2 6076 6349 6076 6349 0 N4BEG[10]
rlabel metal3 6104 6188 6104 6188 0 N4BEG[11]
rlabel metal2 5684 6608 5684 6608 0 N4BEG[12]
rlabel metal2 6412 6349 6412 6349 0 N4BEG[13]
rlabel metal3 6664 6132 6664 6132 0 N4BEG[14]
rlabel metal2 6636 6825 6636 6825 0 N4BEG[15]
rlabel metal2 3780 6692 3780 6692 0 N4BEG[1]
rlabel metal2 4172 6412 4172 6412 0 N4BEG[2]
rlabel metal2 5292 6237 5292 6237 0 N4BEG[3]
rlabel metal2 5404 6461 5404 6461 0 N4BEG[4]
rlabel metal2 5180 5936 5180 5936 0 N4BEG[5]
rlabel metal2 5628 6629 5628 6629 0 N4BEG[6]
rlabel metal2 5796 5600 5796 5600 0 N4BEG[7]
rlabel metal2 4900 6720 4900 6720 0 N4BEG[8]
rlabel metal2 6524 5488 6524 5488 0 N4BEG[9]
rlabel metal2 2156 4704 2156 4704 0 S1END[0]
rlabel metal2 2772 3864 2772 3864 0 S1END[1]
rlabel metal2 3780 3724 3780 3724 0 S1END[2]
rlabel metal2 4816 4172 4816 4172 0 S1END[3]
rlabel metal2 4172 3276 4172 3276 0 S2END[0]
rlabel metal2 2772 6104 2772 6104 0 S2END[1]
rlabel metal2 8092 5880 8092 5880 0 S2END[2]
rlabel metal2 6580 6692 6580 6692 0 S2END[3]
rlabel metal3 8344 6580 8344 6580 0 S2END[4]
rlabel metal2 8260 6748 8260 6748 0 S2END[5]
rlabel metal2 8596 6440 8596 6440 0 S2END[6]
rlabel metal3 8932 6076 8932 6076 0 S2END[7]
rlabel metal3 6440 4116 6440 4116 0 S2MID[0]
rlabel metal2 5572 3668 5572 3668 0 S2MID[1]
rlabel metal3 6216 4340 6216 4340 0 S2MID[2]
rlabel metal2 6160 4564 6160 4564 0 S2MID[3]
rlabel metal3 6328 4172 6328 4172 0 S2MID[4]
rlabel metal2 4788 6384 4788 6384 0 S2MID[5]
rlabel metal2 7364 5852 7364 5852 0 S2MID[6]
rlabel metal2 7420 5348 7420 5348 0 S2MID[7]
rlabel metal2 6692 5656 6692 5656 0 S4END[0]
rlabel metal2 10444 5292 10444 5292 0 S4END[10]
rlabel metal2 10360 5012 10360 5012 0 S4END[11]
rlabel metal2 11172 5572 11172 5572 0 S4END[12]
rlabel metal2 11536 5012 11536 5012 0 S4END[13]
rlabel metal2 12012 4564 12012 4564 0 S4END[14]
rlabel metal2 13860 5516 13860 5516 0 S4END[15]
rlabel metal2 9100 6769 9100 6769 0 S4END[1]
rlabel metal2 9492 6608 9492 6608 0 S4END[2]
rlabel metal2 9772 5936 9772 5936 0 S4END[3]
rlabel metal2 2772 5320 2772 5320 0 S4END[4]
rlabel metal3 4396 3668 4396 3668 0 S4END[5]
rlabel metal2 9604 6244 9604 6244 0 S4END[6]
rlabel metal2 9100 5516 9100 5516 0 S4END[7]
rlabel metal2 9548 5404 9548 5404 0 S4END[8]
rlabel metal2 10164 5208 10164 5208 0 S4END[9]
rlabel metal2 1148 63 1148 63 0 UserCLK
rlabel metal2 10528 5236 10528 5236 0 UserCLKo
rlabel metal2 13356 1176 13356 1176 0 net1
rlabel metal2 14700 3780 14700 3780 0 net10
rlabel metal2 8372 4900 8372 4900 0 net11
rlabel metal3 10024 588 10024 588 0 net12
rlabel metal2 7980 5096 7980 5096 0 net13
rlabel metal2 14756 4760 14756 4760 0 net14
rlabel metal2 14700 5516 14700 5516 0 net15
rlabel metal2 13916 4844 13916 4844 0 net16
rlabel metal2 14028 3472 14028 3472 0 net17
rlabel metal2 8148 2576 8148 2576 0 net18
rlabel metal3 11144 3668 11144 3668 0 net19
rlabel metal2 14756 2184 14756 2184 0 net2
rlabel metal2 11788 4732 11788 4732 0 net20
rlabel metal2 10052 5124 10052 5124 0 net21
rlabel metal4 10500 4508 10500 4508 0 net22
rlabel metal2 8372 588 8372 588 0 net23
rlabel metal2 10948 5824 10948 5824 0 net24
rlabel metal2 15316 5964 15316 5964 0 net25
rlabel metal2 13132 1232 13132 1232 0 net26
rlabel metal2 13860 1148 13860 1148 0 net27
rlabel metal2 13916 1204 13916 1204 0 net28
rlabel metal2 14700 840 14700 840 0 net29
rlabel metal2 13916 2632 13916 2632 0 net3
rlabel metal2 14756 1316 14756 1316 0 net30
rlabel metal2 13916 1960 13916 1960 0 net31
rlabel metal2 14028 1792 14028 1792 0 net32
rlabel metal3 10276 4284 10276 4284 0 net33
rlabel metal3 12096 4396 12096 4396 0 net34
rlabel metal3 11956 4900 11956 4900 0 net35
rlabel metal2 10864 644 10864 644 0 net36
rlabel metal2 12096 1428 12096 1428 0 net37
rlabel metal2 12964 1036 12964 1036 0 net38
rlabel metal2 13916 5432 13916 5432 0 net39
rlabel metal2 8652 2716 8652 2716 0 net4
rlabel metal2 14364 4788 14364 4788 0 net40
rlabel metal2 13580 3360 13580 3360 0 net41
rlabel metal2 14560 4564 14560 4564 0 net42
rlabel metal2 14308 1568 14308 1568 0 net43
rlabel metal3 10556 3836 10556 3836 0 net44
rlabel metal2 10724 1036 10724 1036 0 net45
rlabel metal2 11116 1358 11116 1358 0 net46
rlabel metal3 13132 6020 13132 6020 0 net47
rlabel metal2 1820 5768 1820 5768 0 net48
rlabel metal3 6524 644 6524 644 0 net49
rlabel metal3 11116 2548 11116 2548 0 net5
rlabel metal2 6356 700 6356 700 0 net50
rlabel metal2 6748 1372 6748 1372 0 net51
rlabel metal3 10164 3444 10164 3444 0 net52
rlabel metal2 2156 5152 2156 5152 0 net53
rlabel metal2 3416 3780 3416 3780 0 net54
rlabel metal2 2324 4186 2324 4186 0 net55
rlabel metal3 2240 4452 2240 4452 0 net56
rlabel metal2 1372 5824 1372 5824 0 net57
rlabel metal2 2548 5264 2548 5264 0 net58
rlabel metal2 4508 5880 4508 5880 0 net59
rlabel metal2 13916 3304 13916 3304 0 net6
rlabel metal3 4648 4900 4648 4900 0 net60
rlabel metal2 4172 4312 4172 4312 0 net61
rlabel metal2 4004 4256 4004 4256 0 net62
rlabel metal2 2324 6468 2324 6468 0 net63
rlabel metal2 3276 4984 3276 4984 0 net64
rlabel metal2 3780 5684 3780 5684 0 net65
rlabel metal2 4172 5208 4172 5208 0 net66
rlabel metal2 4788 4564 4788 4564 0 net67
rlabel metal2 3276 6552 3276 6552 0 net68
rlabel metal2 6300 6048 6300 6048 0 net69
rlabel metal2 14756 3276 14756 3276 0 net7
rlabel metal2 4564 5600 4564 5600 0 net70
rlabel metal2 3080 6020 3080 6020 0 net71
rlabel metal2 3892 3388 3892 3388 0 net72
rlabel metal2 14532 5040 14532 5040 0 net73
rlabel metal2 4116 4256 4116 4256 0 net74
rlabel metal2 2996 5628 2996 5628 0 net75
rlabel metal2 5964 6356 5964 6356 0 net76
rlabel metal2 7140 6048 7140 6048 0 net77
rlabel metal2 7252 6132 7252 6132 0 net78
rlabel metal2 6468 5124 6468 5124 0 net79
rlabel metal2 14644 3724 14644 3724 0 net8
rlabel metal2 12124 560 12124 560 0 net80
rlabel metal3 7308 4312 7308 4312 0 net81
rlabel metal2 5348 5320 5348 5320 0 net82
rlabel metal2 10892 5124 10892 5124 0 net83
rlabel metal2 5572 4844 5572 4844 0 net84
rlabel metal2 9828 5404 9828 5404 0 net85
rlabel metal3 7700 5236 7700 5236 0 net86
rlabel metal2 5180 6384 5180 6384 0 net87
rlabel metal2 7028 5712 7028 5712 0 net88
rlabel metal2 10248 532 10248 532 0 net89
rlabel metal2 8484 4284 8484 4284 0 net9
<< properties >>
string FIXED_BBOX 0 0 15848 7112
<< end >>
