module DSP (Tile_X0Y0_UserCLKo,
    Tile_X0Y1_UserCLK,
    Tile_X0Y0_E1BEG,
    Tile_X0Y0_E1END,
    Tile_X0Y0_E2BEG,
    Tile_X0Y0_E2BEGb,
    Tile_X0Y0_E2END,
    Tile_X0Y0_E2MID,
    Tile_X0Y0_E6BEG,
    Tile_X0Y0_E6END,
    Tile_X0Y0_EE4BEG,
    Tile_X0Y0_EE4END,
    Tile_X0Y0_FrameData,
    Tile_X0Y0_FrameData_O,
    Tile_X0Y0_FrameStrobe_O,
    Tile_X0Y0_N1BEG,
    Tile_X0Y0_N2BEG,
    Tile_X0Y0_N2BEGb,
    Tile_X0Y0_N4BEG,
    Tile_X0Y0_NN4BEG,
    Tile_X0Y0_S1END,
    Tile_X0Y0_S2END,
    Tile_X0Y0_S2MID,
    Tile_X0Y0_S4END,
    Tile_X0Y0_SS4END,
    Tile_X0Y0_W1BEG,
    Tile_X0Y0_W1END,
    Tile_X0Y0_W2BEG,
    Tile_X0Y0_W2BEGb,
    Tile_X0Y0_W2END,
    Tile_X0Y0_W2MID,
    Tile_X0Y0_W6BEG,
    Tile_X0Y0_W6END,
    Tile_X0Y0_WW4BEG,
    Tile_X0Y0_WW4END,
    Tile_X0Y1_E1BEG,
    Tile_X0Y1_E1END,
    Tile_X0Y1_E2BEG,
    Tile_X0Y1_E2BEGb,
    Tile_X0Y1_E2END,
    Tile_X0Y1_E2MID,
    Tile_X0Y1_E6BEG,
    Tile_X0Y1_E6END,
    Tile_X0Y1_EE4BEG,
    Tile_X0Y1_EE4END,
    Tile_X0Y1_FrameData,
    Tile_X0Y1_FrameData_O,
    Tile_X0Y1_FrameStrobe,
    Tile_X0Y1_N1END,
    Tile_X0Y1_N2END,
    Tile_X0Y1_N2MID,
    Tile_X0Y1_N4END,
    Tile_X0Y1_NN4END,
    Tile_X0Y1_S1BEG,
    Tile_X0Y1_S2BEG,
    Tile_X0Y1_S2BEGb,
    Tile_X0Y1_S4BEG,
    Tile_X0Y1_SS4BEG,
    Tile_X0Y1_W1BEG,
    Tile_X0Y1_W1END,
    Tile_X0Y1_W2BEG,
    Tile_X0Y1_W2BEGb,
    Tile_X0Y1_W2END,
    Tile_X0Y1_W2MID,
    Tile_X0Y1_W6BEG,
    Tile_X0Y1_W6END,
    Tile_X0Y1_WW4BEG,
    Tile_X0Y1_WW4END);
 output Tile_X0Y0_UserCLKo;
 input Tile_X0Y1_UserCLK;
 output [3:0] Tile_X0Y0_E1BEG;
 input [3:0] Tile_X0Y0_E1END;
 output [7:0] Tile_X0Y0_E2BEG;
 output [7:0] Tile_X0Y0_E2BEGb;
 input [7:0] Tile_X0Y0_E2END;
 input [7:0] Tile_X0Y0_E2MID;
 output [11:0] Tile_X0Y0_E6BEG;
 input [11:0] Tile_X0Y0_E6END;
 output [15:0] Tile_X0Y0_EE4BEG;
 input [15:0] Tile_X0Y0_EE4END;
 input [31:0] Tile_X0Y0_FrameData;
 output [31:0] Tile_X0Y0_FrameData_O;
 output [19:0] Tile_X0Y0_FrameStrobe_O;
 output [3:0] Tile_X0Y0_N1BEG;
 output [7:0] Tile_X0Y0_N2BEG;
 output [7:0] Tile_X0Y0_N2BEGb;
 output [15:0] Tile_X0Y0_N4BEG;
 output [15:0] Tile_X0Y0_NN4BEG;
 input [3:0] Tile_X0Y0_S1END;
 input [7:0] Tile_X0Y0_S2END;
 input [7:0] Tile_X0Y0_S2MID;
 input [15:0] Tile_X0Y0_S4END;
 input [15:0] Tile_X0Y0_SS4END;
 output [3:0] Tile_X0Y0_W1BEG;
 input [3:0] Tile_X0Y0_W1END;
 output [7:0] Tile_X0Y0_W2BEG;
 output [7:0] Tile_X0Y0_W2BEGb;
 input [7:0] Tile_X0Y0_W2END;
 input [7:0] Tile_X0Y0_W2MID;
 output [11:0] Tile_X0Y0_W6BEG;
 input [11:0] Tile_X0Y0_W6END;
 output [15:0] Tile_X0Y0_WW4BEG;
 input [15:0] Tile_X0Y0_WW4END;
 output [3:0] Tile_X0Y1_E1BEG;
 input [3:0] Tile_X0Y1_E1END;
 output [7:0] Tile_X0Y1_E2BEG;
 output [7:0] Tile_X0Y1_E2BEGb;
 input [7:0] Tile_X0Y1_E2END;
 input [7:0] Tile_X0Y1_E2MID;
 output [11:0] Tile_X0Y1_E6BEG;
 input [11:0] Tile_X0Y1_E6END;
 output [15:0] Tile_X0Y1_EE4BEG;
 input [15:0] Tile_X0Y1_EE4END;
 input [31:0] Tile_X0Y1_FrameData;
 output [31:0] Tile_X0Y1_FrameData_O;
 input [19:0] Tile_X0Y1_FrameStrobe;
 input [3:0] Tile_X0Y1_N1END;
 input [7:0] Tile_X0Y1_N2END;
 input [7:0] Tile_X0Y1_N2MID;
 input [15:0] Tile_X0Y1_N4END;
 input [15:0] Tile_X0Y1_NN4END;
 output [3:0] Tile_X0Y1_S1BEG;
 output [7:0] Tile_X0Y1_S2BEG;
 output [7:0] Tile_X0Y1_S2BEGb;
 output [15:0] Tile_X0Y1_S4BEG;
 output [15:0] Tile_X0Y1_SS4BEG;
 output [3:0] Tile_X0Y1_W1BEG;
 input [3:0] Tile_X0Y1_W1END;
 output [7:0] Tile_X0Y1_W2BEG;
 output [7:0] Tile_X0Y1_W2BEGb;
 input [7:0] Tile_X0Y1_W2END;
 input [7:0] Tile_X0Y1_W2MID;
 output [11:0] Tile_X0Y1_W6BEG;
 input [11:0] Tile_X0Y1_W6END;
 output [15:0] Tile_X0Y1_WW4BEG;
 input [15:0] Tile_X0Y1_WW4END;

 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire \Tile_X0Y1_DSP_bot.A0 ;
 wire \Tile_X0Y1_DSP_bot.A1 ;
 wire \Tile_X0Y1_DSP_bot.A2 ;
 wire \Tile_X0Y1_DSP_bot.A3 ;
 wire \Tile_X0Y1_DSP_bot.B0 ;
 wire \Tile_X0Y1_DSP_bot.B1 ;
 wire \Tile_X0Y1_DSP_bot.B2 ;
 wire \Tile_X0Y1_DSP_bot.B3 ;
 wire \Tile_X0Y1_DSP_bot.C0 ;
 wire \Tile_X0Y1_DSP_bot.C1 ;
 wire \Tile_X0Y1_DSP_bot.C2 ;
 wire \Tile_X0Y1_DSP_bot.C3 ;
 wire \Tile_X0Y1_DSP_bot.C4 ;
 wire \Tile_X0Y1_DSP_bot.C5 ;
 wire \Tile_X0Y1_DSP_bot.C6 ;
 wire \Tile_X0Y1_DSP_bot.C7 ;
 wire \Tile_X0Y1_DSP_bot.C8 ;
 wire \Tile_X0Y1_DSP_bot.C9 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[10] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[11] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[12] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[13] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[14] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[15] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[16] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[17] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[18] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[8] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[9] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[10] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[11] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[12] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[13] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[14] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[15] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[16] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[17] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[18] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[19] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[8] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[9] ;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire Tile_X0Y1_UserCLK_regs;
 wire clknet_0_Tile_X0Y1_UserCLK;
 wire clknet_1_0__leaf_Tile_X0Y1_UserCLK;
 wire clknet_0_Tile_X0Y1_UserCLK_regs;
 wire clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs;
 wire clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs;
 wire clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs;
 wire clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs;

 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2267_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2268_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2269_ (.A1(_0069_),
    .A2(_0610_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2270_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ),
    .A2(_0609_),
    .B(_0070_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2271_ (.I0(Tile_X0Y1_N2MID[4]),
    .I1(Tile_X0Y0_E2END[4]),
    .I2(Tile_X0Y0_E1END[2]),
    .I3(Tile_X0Y0_E6END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2272_ (.A1(_0069_),
    .A2(_0613_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2273_ (.I0(Tile_X0Y0_S2END[4]),
    .I1(Tile_X0Y0_W2END[4]),
    .I2(Tile_X0Y0_S4END[0]),
    .I3(Tile_X0Y0_WW4END[2]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2274_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ),
    .A2(_0615_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2275_ (.A1(_0611_),
    .A2(_0612_),
    .B1(_0614_),
    .B2(_0616_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2276_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2277_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2278_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2279_ (.I0(_0618_),
    .I1(_0619_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2280_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0620_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2281_ (.I(_0621_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2282_ (.A1(_0499_),
    .A2(_0502_),
    .B(_0509_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2283_ (.A1(_0498_),
    .A2(_0503_),
    .B(_0508_),
    .C(_0062_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2284_ (.A1(_0061_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2285_ (.A1(Tile_X0Y0_E2MID[7]),
    .A2(_0062_),
    .B(_0065_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2286_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ),
    .A2(_0064_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2287_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ),
    .A2(Tile_X0Y0_S2MID[7]),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ),
    .C(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2288_ (.I(_0628_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2289_ (.A1(_0623_),
    .A2(_0626_),
    .B(_0628_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2290_ (.A1(_0624_),
    .A2(_0625_),
    .B(_0629_),
    .C(_0099_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2291_ (.A1(_0623_),
    .A2(_0626_),
    .B(_0628_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2292_ (.A1(_0099_),
    .A2(_0208_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q ),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2293_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .B(_0102_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2294_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2295_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .A2(_0208_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2296_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .B(_0636_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2297_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2298_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .A2(_0211_),
    .B(_0638_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2299_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ),
    .A2(_0639_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2300_ (.A1(_0637_),
    .A2(_0640_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2301_ (.A1(_0101_),
    .A2(_0635_),
    .B(_0641_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2302_ (.I0(_0456_),
    .I1(Tile_X0Y1_N4END[5]),
    .I2(Tile_X0Y1_N2MID[1]),
    .I3(Tile_X0Y0_EE4END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2303_ (.A1(_0101_),
    .A2(_0643_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2304_ (.I0(Tile_X0Y0_E6END[1]),
    .I1(Tile_X0Y0_S2END[1]),
    .I2(Tile_X0Y0_W2END[1]),
    .I3(Tile_X0Y0_W6END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2305_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ),
    .A2(_0645_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2306_ (.A1(_0644_),
    .A2(_0646_),
    .B(_0642_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2307_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2308_ (.A1(Tile_X0Y0_W2END[4]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q ),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2309_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q ),
    .A2(_0617_),
    .B(_0648_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2310_ (.A1(Tile_X0Y1_N4END[5]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q ),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2311_ (.A1(_0068_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q ),
    .C(_0650_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2312_ (.A1(_0649_),
    .A2(_0651_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2313_ (.I(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2314_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ),
    .A2(_0652_),
    .B(_0647_),
    .C(_0102_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2315_ (.I(_0654_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2316_ (.A1(_0632_),
    .A2(_0633_),
    .B(_0654_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2317_ (.I(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2318_ (.A1(_0632_),
    .A2(_0633_),
    .B(_0654_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2319_ (.A1(_0631_),
    .A2(_0634_),
    .B(_0655_),
    .C(_0098_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2320_ (.A1(Tile_X0Y0_S2MID[5]),
    .A2(_0098_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2321_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .A2(_0660_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2322_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .A2(_0660_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2323_ (.A1(Tile_X0Y1_W1END[3]),
    .A2(_0098_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2324_ (.A1(Tile_X0Y1_W1END[1]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2325_ (.A1(_0663_),
    .A2(_0664_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2326_ (.A1(_0659_),
    .A2(_0661_),
    .B(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2327_ (.A1(_0658_),
    .A2(_0662_),
    .B1(_0663_),
    .B2(_0664_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2328_ (.I0(Tile_X0Y1_N1END[1]),
    .I1(Tile_X0Y1_N2END[5]),
    .I2(Tile_X0Y1_E1END[1]),
    .I3(Tile_X0Y1_E2END[5]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2329_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(_0668_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2330_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0669_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2331_ (.I(_0670_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2332_ (.A1(_0667_),
    .A2(_0670_),
    .B(_0621_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2333_ (.I(_0672_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2334_ (.I0(_0672_),
    .I1(_0104_),
    .I2(_0103_),
    .I3(_0617_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2335_ (.I(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2336_ (.A1(_0105_),
    .A2(_0374_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2337_ (.A1(_0105_),
    .A2(_0673_),
    .B(_0675_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q ),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2338_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q ),
    .A2(_0608_),
    .B(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2339_ (.I(_0677_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2340_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[6] ),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2341_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(_0677_),
    .B(_0678_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2342_ (.I(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2343_ (.A1(_0375_),
    .A2(_0377_),
    .B(_0410_),
    .C(_0138_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2344_ (.A1(_0632_),
    .A2(_0633_),
    .B(_0654_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2345_ (.A1(_0096_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2346_ (.A1(Tile_X0Y0_S2MID[5]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .C(_0683_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2347_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .A2(_0684_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2348_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .A2(_0681_),
    .A3(_0682_),
    .B(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2349_ (.I0(Tile_X0Y1_N1END[1]),
    .I1(Tile_X0Y1_N2END[5]),
    .I2(Tile_X0Y1_E1END[1]),
    .I3(Tile_X0Y1_E2END[5]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2350_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .A2(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2351_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2352_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2353_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2354_ (.I0(_0691_),
    .I1(_0690_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2355_ (.A1(_0686_),
    .A2(_0689_),
    .B1(_0692_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2356_ (.A1(_0686_),
    .A2(_0689_),
    .B1(_0692_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .C(_0137_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2357_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .A2(Tile_X0Y1_W2MID[0]),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2358_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2359_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2360_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2361_ (.A1(_0092_),
    .A2(_0698_),
    .B(_0093_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2362_ (.I0(Tile_X0Y1_NN4END[5]),
    .I1(Tile_X0Y0_E1END[3]),
    .I2(Tile_X0Y0_E2END[1]),
    .I3(Tile_X0Y0_E6END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2363_ (.A1(_0092_),
    .A2(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2364_ (.I0(Tile_X0Y0_S2END[1]),
    .I1(Tile_X0Y0_S4END[1]),
    .I2(Tile_X0Y0_W2END[1]),
    .I3(Tile_X0Y0_W6END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2365_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(_0702_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2366_ (.A1(_0697_),
    .A2(_0699_),
    .B1(_0701_),
    .B2(_0703_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2367_ (.A1(_0046_),
    .A2(_0137_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2368_ (.A1(_0137_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .B(_0704_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2369_ (.A1(_0694_),
    .A2(_0695_),
    .B1(_0705_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .C(_0139_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2370_ (.A1(_0139_),
    .A2(_0254_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2371_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ),
    .A2(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2372_ (.A1(_0706_),
    .A2(_0708_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2373_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .A2(_0445_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2374_ (.A1(Tile_X0Y1_W6END[0]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q ),
    .C(_0710_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2375_ (.A1(_0140_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q ),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2376_ (.A1(Tile_X0Y1_N4END[0]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .B(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2377_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ),
    .A2(_0711_),
    .A3(_0713_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2378_ (.I0(Tile_X0Y1_N2END[0]),
    .I1(Tile_X0Y0_S2MID[0]),
    .I2(Tile_X0Y1_EE4END[1]),
    .I3(Tile_X0Y1_W2END[0]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q ),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2379_ (.I(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2380_ (.A1(_0139_),
    .A2(_0716_),
    .B(_0141_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2381_ (.A1(_0714_),
    .A2(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2382_ (.A1(_0709_),
    .A2(_0718_),
    .ZN(\Tile_X0Y1_DSP_bot.B3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2383_ (.A1(_0706_),
    .A2(_0708_),
    .B1(_0714_),
    .B2(_0717_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2384_ (.A1(_0131_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[3] ),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2385_ (.A1(_0719_),
    .A2(_0720_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2386_ (.A1(_0679_),
    .A2(_0721_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2387_ (.A1(_0551_),
    .A2(_0679_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2388_ (.A1(_0598_),
    .A2(_0721_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2389_ (.A1(_0723_),
    .A2(_0724_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2390_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .A2(_0241_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2391_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .B(_0726_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2392_ (.A1(Tile_X0Y1_N2MID[0]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2393_ (.A1(_0133_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .C(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2394_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .A2(_0729_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2395_ (.I0(_0033_),
    .I1(_0034_),
    .I2(_0253_),
    .I3(_0038_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q ),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2396_ (.A1(_0727_),
    .A2(_0730_),
    .B1(_0731_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q ),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2397_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2398_ (.A1(_0135_),
    .A2(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2399_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2400_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .A2(_0735_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2401_ (.I0(Tile_X0Y1_N1END[0]),
    .I1(Tile_X0Y1_N2END[2]),
    .I2(Tile_X0Y1_E2END[2]),
    .I3(Tile_X0Y1_E6END[0]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2402_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .A2(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2403_ (.I0(Tile_X0Y0_S2MID[2]),
    .I1(Tile_X0Y1_W2END[2]),
    .I2(Tile_X0Y0_S4END[6]),
    .I3(Tile_X0Y1_W6END[0]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2404_ (.A1(_0135_),
    .A2(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2405_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .A2(_0738_),
    .A3(_0740_),
    .B1(_0734_),
    .B2(_0736_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2406_ (.I0(Tile_X0Y1_N4END[0]),
    .I1(Tile_X0Y0_S4END[4]),
    .I2(Tile_X0Y1_E6END[0]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2407_ (.I0(Tile_X0Y1_N2END[0]),
    .I1(Tile_X0Y0_S2MID[0]),
    .I2(Tile_X0Y1_E2END[0]),
    .I3(Tile_X0Y1_WW4END[3]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q ),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2408_ (.I(_0742_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2409_ (.I0(_0742_),
    .I1(_0741_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2410_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q ),
    .A2(_0744_),
    .B(_0732_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2411_ (.I(_0745_),
    .ZN(\Tile_X0Y1_DSP_bot.A3 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2412_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[3] ),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2413_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(_0745_),
    .B(_0746_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2414_ (.I(_0747_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2415_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .I1(Tile_X0Y0_W2MID[0]),
    .I2(Tile_X0Y0_S2MID[0]),
    .I3(_0316_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2416_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0483_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q ),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2417_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0749_),
    .B(_0750_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2418_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2419_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .A2(_0210_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2420_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .B(_0753_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2421_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .A2(_0213_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2422_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .B(_0755_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2423_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .A2(_0754_),
    .B(_0756_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2424_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ),
    .A2(_0752_),
    .B(_0757_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2425_ (.I0(_0306_),
    .I1(Tile_X0Y0_E2END[3]),
    .I2(Tile_X0Y1_N2MID[3]),
    .I3(Tile_X0Y0_E6END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2426_ (.I0(Tile_X0Y0_S2END[3]),
    .I1(Tile_X0Y0_W2END[3]),
    .I2(Tile_X0Y0_S4END[3]),
    .I3(Tile_X0Y0_W6END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2427_ (.I(_0760_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2428_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ),
    .A2(_0761_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2429_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ),
    .A2(_0759_),
    .B(_0762_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2430_ (.A1(_0758_),
    .A2(_0763_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2431_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2432_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ),
    .A2(_0764_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2433_ (.A1(Tile_X0Y0_W6END[0]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q ),
    .C(_0765_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2434_ (.A1(_0118_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q ),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2435_ (.A1(Tile_X0Y1_N4END[4]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ),
    .B(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2436_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0766_),
    .A3(_0768_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2437_ (.I0(Tile_X0Y1_N2MID[0]),
    .I1(Tile_X0Y0_S2END[0]),
    .I2(Tile_X0Y0_EE4END[1]),
    .I3(Tile_X0Y0_W2END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q ),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2438_ (.I(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2439_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0770_),
    .B(_0769_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q ),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2440_ (.A1(_0751_),
    .A2(_0772_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2441_ (.I(_0773_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2442_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[7] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2443_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .A2(_0773_),
    .B(_0774_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2444_ (.I(_0775_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2445_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2446_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .A2(_0209_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2447_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .B(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2448_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .A2(_0215_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2449_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .B(_0780_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2450_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ),
    .A2(_0779_),
    .A3(_0781_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2451_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ),
    .A2(_0777_),
    .B(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2452_ (.I0(Tile_X0Y1_NN4END[7]),
    .I1(Tile_X0Y0_E1END[1]),
    .I2(Tile_X0Y0_E2END[3]),
    .I3(Tile_X0Y0_E6END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2453_ (.I0(Tile_X0Y0_S2END[3]),
    .I1(Tile_X0Y0_W2END[3]),
    .I2(Tile_X0Y0_S4END[3]),
    .I3(Tile_X0Y0_W6END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2454_ (.I0(_0784_),
    .I1(_0785_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2455_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ),
    .A2(_0786_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2456_ (.A1(_0783_),
    .A2(_0787_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2457_ (.I(_0788_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2458_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ),
    .A2(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2459_ (.A1(Tile_X0Y0_S4END[1]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q ),
    .C(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2460_ (.A1(Tile_X0Y1_NN4END[5]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2461_ (.A1(_0100_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q ),
    .C(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2462_ (.A1(_0116_),
    .A2(_0792_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2463_ (.I0(Tile_X0Y1_N2MID[4]),
    .I1(Tile_X0Y0_E2END[4]),
    .I2(Tile_X0Y0_SS4END[2]),
    .I3(Tile_X0Y0_W2END[4]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q ),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2464_ (.I(_0794_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2465_ (.A1(_0790_),
    .A2(_0793_),
    .B1(_0795_),
    .B2(_0116_),
    .C(_0117_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2466_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2467_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .A2(_0208_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2468_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .B(_0798_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2469_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2470_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .A2(_0211_),
    .B(_0800_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2471_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2472_ (.A1(_0799_),
    .A2(_0802_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2473_ (.A1(_0115_),
    .A2(_0797_),
    .B(_0803_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2474_ (.I0(_0306_),
    .I1(Tile_X0Y0_E1END[1]),
    .I2(Tile_X0Y1_N2MID[5]),
    .I3(Tile_X0Y0_E2END[5]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2475_ (.A1(_0115_),
    .A2(_0805_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2476_ (.I0(Tile_X0Y0_S1END[1]),
    .I1(Tile_X0Y0_W1END[1]),
    .I2(Tile_X0Y0_S2END[5]),
    .I3(Tile_X0Y0_W1END[3]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2477_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(_0807_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2478_ (.A1(_0806_),
    .A2(_0808_),
    .B(_0804_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2479_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2480_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ),
    .A2(_0809_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2481_ (.A1(Tile_X0Y0_S2MID[4]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ),
    .C(_0810_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2482_ (.A1(_0667_),
    .A2(_0670_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ),
    .C(_0621_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2483_ (.A1(_0103_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2484_ (.I(_0813_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2485_ (.A1(_0812_),
    .A2(_0814_),
    .B(_0811_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2486_ (.I(_0815_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2487_ (.A1(_0812_),
    .A2(_0814_),
    .B(_0116_),
    .C(_0811_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2488_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .I1(Tile_X0Y0_S2MID[5]),
    .I2(Tile_X0Y0_E2MID[5]),
    .I3(Tile_X0Y0_W2MID[5]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2489_ (.A1(_0116_),
    .A2(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2490_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q ),
    .A2(_0819_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2491_ (.A1(_0817_),
    .A2(_0820_),
    .B(_0796_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2492_ (.I(_0821_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X ));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2493_ (.A1(_0817_),
    .A2(_0820_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .C(_0796_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2494_ (.A1(_0131_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[6] ),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2495_ (.A1(_0822_),
    .A2(_0823_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2496_ (.I(_0824_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2497_ (.I0(Tile_X0Y1_N2MID[4]),
    .I1(Tile_X0Y1_E2MID[4]),
    .I2(Tile_X0Y1_W2MID[4]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q ),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2498_ (.I(_0826_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2499_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2500_ (.A1(_0136_),
    .A2(_0828_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2501_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2502_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .A2(_0830_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2503_ (.I0(Tile_X0Y1_NN4END[2]),
    .I1(Tile_X0Y1_EE4END[2]),
    .I2(Tile_X0Y1_E1END[0]),
    .I3(Tile_X0Y1_E6END[0]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2504_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .A2(_0832_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2505_ (.I0(Tile_X0Y0_S4END[6]),
    .I1(Tile_X0Y0_SS4END[6]),
    .I2(Tile_X0Y1_W2END[2]),
    .I3(Tile_X0Y1_W6END[0]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2506_ (.A1(_0136_),
    .A2(_0834_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2507_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .A2(_0833_),
    .A3(_0835_),
    .B1(_0829_),
    .B2(_0831_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2508_ (.I0(Tile_X0Y1_N4END[1]),
    .I1(Tile_X0Y1_W6END[1]),
    .I2(Tile_X0Y1_E6END[1]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q ),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2509_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0836_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2510_ (.I0(Tile_X0Y1_N2END[4]),
    .I1(Tile_X0Y0_S2MID[4]),
    .I2(Tile_X0Y1_EE4END[0]),
    .I3(Tile_X0Y1_W2END[4]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q ),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2511_ (.I(_0838_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2512_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0455_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q ),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2513_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0827_),
    .B(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2514_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0839_),
    .B(_0837_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q ),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2515_ (.A1(_0841_),
    .A2(_0842_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2516_ (.I(_0843_),
    .ZN(\Tile_X0Y1_DSP_bot.A2 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2517_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(_0843_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2518_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[2] ),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2519_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(_0843_),
    .B(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2520_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[2] ),
    .B(_0844_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2521_ (.A1(_0822_),
    .A2(_0823_),
    .A3(_0847_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2522_ (.A1(_0748_),
    .A2(_0822_),
    .A3(_0823_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2523_ (.A1(_0776_),
    .A2(_0847_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2524_ (.I(_0850_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2525_ (.A1(_0849_),
    .A2(_0850_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2526_ (.A1(_0849_),
    .A2(_0850_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2527_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2528_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .A2(_0208_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2529_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .B(_0855_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2530_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2531_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .A2(_0211_),
    .B(_0857_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2532_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_0858_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2533_ (.A1(_0856_),
    .A2(_0859_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2534_ (.A1(_0113_),
    .A2(_0854_),
    .B(_0860_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2535_ (.I0(_0306_),
    .I1(Tile_X0Y0_E1END[1]),
    .I2(Tile_X0Y1_N2MID[5]),
    .I3(Tile_X0Y0_E2END[5]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2536_ (.A1(_0113_),
    .A2(_0862_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2537_ (.I0(Tile_X0Y0_S1END[1]),
    .I1(Tile_X0Y0_S2END[5]),
    .I2(Tile_X0Y0_S1END[3]),
    .I3(Tile_X0Y0_W1END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2538_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_0864_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2539_ (.A1(_0863_),
    .A2(_0865_),
    .B(_0861_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2540_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2541_ (.A1(_0111_),
    .A2(_0866_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2542_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2543_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .A2(_0868_),
    .B(_0112_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2544_ (.I0(Tile_X0Y1_N2END[3]),
    .I1(Tile_X0Y1_N4END[3]),
    .I2(Tile_X0Y1_E1END[1]),
    .I3(Tile_X0Y1_E2END[3]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2545_ (.A1(_0111_),
    .A2(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2546_ (.I0(Tile_X0Y1_E6END[1]),
    .I1(Tile_X0Y0_S2MID[3]),
    .I2(Tile_X0Y1_W2END[3]),
    .I3(Tile_X0Y1_WW4END[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2547_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .A2(_0872_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q ),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2548_ (.A1(_0867_),
    .A2(_0869_),
    .B1(_0871_),
    .B2(_0873_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2549_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .I1(Tile_X0Y0_W2MID[2]),
    .I2(Tile_X0Y0_E2MID[2]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q ),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2550_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .I1(Tile_X0Y0_E2MID[3]),
    .I2(Tile_X0Y0_S2MID[3]),
    .I3(Tile_X0Y0_W2MID[3]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q ),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2551_ (.A1(_0114_),
    .A2(_0875_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2552_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ),
    .A2(_0874_),
    .B(_0876_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2553_ (.A1(_0114_),
    .A2(_0468_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2554_ (.I0(Tile_X0Y1_N2MID[2]),
    .I1(Tile_X0Y0_S2END[2]),
    .I2(Tile_X0Y0_E2END[2]),
    .I3(Tile_X0Y0_WW4END[2]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q ),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2555_ (.I(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2556_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ),
    .A2(_0879_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q ),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2557_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q ),
    .A2(_0877_),
    .B1(_0878_),
    .B2(_0881_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2558_ (.I0(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[5] ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ),
    .S(_0131_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2559_ (.I(_0882_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2560_ (.I0(Tile_X0Y1_N2MID[6]),
    .I1(Tile_X0Y0_E2END[6]),
    .I2(Tile_X0Y0_SS4END[3]),
    .I3(Tile_X0Y0_W2END[6]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q ),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2561_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0884_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q ),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2562_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0408_),
    .B(_0885_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2563_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0218_),
    .B1(_0417_),
    .B2(_0420_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2564_ (.A1(_0083_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2565_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .Z(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2566_ (.A1(_0089_),
    .A2(_0889_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2567_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2568_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ),
    .A2(_0891_),
    .B(_0090_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2569_ (.I0(Tile_X0Y1_N2MID[4]),
    .I1(Tile_X0Y1_N4END[4]),
    .I2(Tile_X0Y0_E1END[2]),
    .I3(Tile_X0Y0_E2END[4]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2570_ (.A1(_0089_),
    .A2(_0893_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2571_ (.I0(Tile_X0Y0_E6END[0]),
    .I1(Tile_X0Y0_S2END[4]),
    .I2(Tile_X0Y0_W2END[4]),
    .I3(Tile_X0Y0_W6END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2572_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ),
    .A2(_0895_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2573_ (.A1(_0890_),
    .A2(_0892_),
    .B1(_0894_),
    .B2(_0896_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2574_ (.I0(Tile_X0Y0_W2MID[6]),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2575_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q ),
    .A2(_0897_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2576_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q ),
    .A2(_0887_),
    .A3(_0888_),
    .B(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2577_ (.A1(_0061_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q ),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2578_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ),
    .B(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2579_ (.A1(_0064_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2580_ (.A1(Tile_X0Y0_S2MID[7]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q ),
    .C(_0902_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2581_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0903_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2582_ (.A1(_0901_),
    .A2(_0904_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q ),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2583_ (.A1(_0899_),
    .A2(_0905_),
    .B(_0886_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2584_ (.I(_0906_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2585_ (.I0(_0906_),
    .I1(_0132_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2586_ (.A1(_0883_),
    .A2(_0907_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2587_ (.A1(_0853_),
    .A2(_0908_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2588_ (.A1(_0852_),
    .A2(_0909_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2589_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2590_ (.A1(_0071_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q ),
    .C(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2591_ (.A1(Tile_X0Y0_S2MID[3]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q ),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2592_ (.A1(_0074_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q ),
    .B(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2593_ (.A1(_0912_),
    .A2(_0914_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2594_ (.A1(_0912_),
    .A2(_0914_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2595_ (.I0(Tile_X0Y0_E2MID[2]),
    .I1(Tile_X0Y0_W2MID[2]),
    .I2(Tile_X0Y0_S2MID[2]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q ),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2596_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ),
    .A2(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2597_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ),
    .A2(_0916_),
    .B(_0918_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q ),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2598_ (.I0(Tile_X0Y0_EE4END[2]),
    .I1(Tile_X0Y0_S4END[2]),
    .I2(Tile_X0Y0_W2END[7]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q ),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2599_ (.I0(Tile_X0Y1_NN4END[4]),
    .I1(Tile_X0Y0_S2END[2]),
    .I2(Tile_X0Y0_E2END[2]),
    .I3(Tile_X0Y0_W2END[2]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q ),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2600_ (.I(_0921_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2601_ (.I0(_0921_),
    .I1(_0920_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2602_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q ),
    .A2(_0923_),
    .B(_0919_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2603_ (.I(_0924_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2604_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2605_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[5] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .B(_0925_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2606_ (.I(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2607_ (.A1(_0882_),
    .A2(_0927_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2608_ (.A1(_0776_),
    .A2(_0907_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2609_ (.A1(_0849_),
    .A2(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2610_ (.A1(_0748_),
    .A2(_0776_),
    .B1(_0825_),
    .B2(_0907_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2611_ (.A1(_0930_),
    .A2(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2612_ (.A1(_0928_),
    .A2(_0932_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2613_ (.A1(_0910_),
    .A2(_0933_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2614_ (.A1(_0723_),
    .A2(_0724_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2615_ (.A1(_0910_),
    .A2(_0933_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2616_ (.A1(_0935_),
    .A2(_0936_),
    .B(_0934_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2617_ (.A1(_0928_),
    .A2(_0932_),
    .B(_0930_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2618_ (.A1(_0680_),
    .A2(_0883_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2619_ (.A1(_0775_),
    .A2(_0927_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2620_ (.A1(_0825_),
    .A2(_0926_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2621_ (.A1(_0929_),
    .A2(_0941_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2622_ (.A1(_0929_),
    .A2(_0941_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2623_ (.A1(_0939_),
    .A2(_0943_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2624_ (.A1(_0939_),
    .A2(_0943_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2625_ (.A1(_0938_),
    .A2(_0945_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2626_ (.A1(_0938_),
    .A2(_0945_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2627_ (.I(_0947_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2628_ (.A1(_0600_),
    .A2(_0947_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2629_ (.A1(_0937_),
    .A2(_0949_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2630_ (.A1(_0725_),
    .A2(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2631_ (.I0(Tile_X0Y1_N2MID[3]),
    .I1(Tile_X0Y1_E2MID[3]),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2632_ (.A1(_0144_),
    .A2(_0952_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2633_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .I1(Tile_X0Y1_W2MID[3]),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2634_ (.I0(_0952_),
    .I1(_0954_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q ),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2635_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q ),
    .A2(_0954_),
    .B(_0953_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2636_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2637_ (.A1(_0145_),
    .A2(_0957_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2638_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2639_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .A2(_0959_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2640_ (.I0(Tile_X0Y1_N1END[0]),
    .I1(Tile_X0Y1_N2END[2]),
    .I2(Tile_X0Y1_N4END[2]),
    .I3(Tile_X0Y1_E2END[2]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2641_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .A2(_0961_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2642_ (.I0(Tile_X0Y1_E6END[0]),
    .I1(Tile_X0Y1_W2END[2]),
    .I2(Tile_X0Y0_S2MID[2]),
    .I3(Tile_X0Y1_WW4END[3]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2643_ (.A1(_0145_),
    .A2(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2644_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ),
    .A2(_0962_),
    .A3(_0964_),
    .B1(_0958_),
    .B2(_0960_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2645_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2646_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .A2(_0965_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2647_ (.A1(Tile_X0Y1_W2END[7]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q ),
    .C(_0966_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2648_ (.A1(_0134_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q ),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2649_ (.A1(Tile_X0Y1_EE4END[2]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .B(_0968_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2650_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2651_ (.A1(_0142_),
    .A2(_0970_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2652_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2653_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .A2(_0972_),
    .B(_0143_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2654_ (.I0(Tile_X0Y1_N1END[2]),
    .I1(Tile_X0Y1_N2END[4]),
    .I2(Tile_X0Y1_N4END[0]),
    .I3(Tile_X0Y1_E2END[4]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2655_ (.A1(_0142_),
    .A2(_0974_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2656_ (.I0(Tile_X0Y1_E6END[0]),
    .I1(Tile_X0Y0_S2MID[4]),
    .I2(Tile_X0Y1_W2END[4]),
    .I3(Tile_X0Y1_W6END[0]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2657_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .A2(_0976_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q ),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2658_ (.A1(_0971_),
    .A2(_0973_),
    .B1(_0975_),
    .B2(_0977_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2659_ (.I0(Tile_X0Y1_NN4END[0]),
    .I1(Tile_X0Y0_S2MID[2]),
    .I2(Tile_X0Y1_E2END[2]),
    .I3(Tile_X0Y1_W2END[2]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q ),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2660_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_0956_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2661_ (.I0(Tile_X0Y1_W2MID[2]),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2662_ (.A1(Tile_X0Y1_E2MID[2]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2663_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ),
    .A2(_0788_),
    .B(_0981_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q ),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2664_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q ),
    .A2(_0980_),
    .B(_0982_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2665_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_0967_),
    .A3(_0969_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2666_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_0978_),
    .B(_0984_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2667_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ),
    .A2(_0979_),
    .A3(_0983_),
    .B(_0985_),
    .ZN(\Tile_X0Y1_DSP_bot.A1 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2668_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(\Tile_X0Y1_DSP_bot.A1 ),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2669_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(_0146_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2670_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(_0146_),
    .B(_0986_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2671_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(\Tile_X0Y1_DSP_bot.A1 ),
    .B(_0987_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2672_ (.A1(_0822_),
    .A2(_0823_),
    .A3(_0989_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2673_ (.A1(_0775_),
    .A2(_0988_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2674_ (.A1(_0848_),
    .A2(_0991_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2675_ (.A1(_0747_),
    .A2(_0882_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2676_ (.A1(_0882_),
    .A2(_0992_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2677_ (.A1(_0851_),
    .A2(_0990_),
    .B1(_0994_),
    .B2(_0748_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2678_ (.A1(_0853_),
    .A2(_0908_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2679_ (.A1(_0995_),
    .A2(_0996_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2680_ (.A1(_0995_),
    .A2(_0996_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2681_ (.A1(_0632_),
    .A2(_0633_),
    .B(_0654_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2682_ (.A1(_0631_),
    .A2(_0634_),
    .B(_0655_),
    .C(_0148_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2683_ (.A1(Tile_X0Y0_S2MID[5]),
    .A2(_0148_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2684_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .A2(_1001_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2685_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .A2(_1001_),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2686_ (.A1(Tile_X0Y1_W1END[3]),
    .A2(_0148_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2687_ (.A1(Tile_X0Y1_W1END[1]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2688_ (.A1(_1004_),
    .A2(_1005_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2689_ (.A1(_1000_),
    .A2(_1002_),
    .B(_1006_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2690_ (.A1(_0999_),
    .A2(_1003_),
    .B1(_1004_),
    .B2(_1005_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2691_ (.I0(Tile_X0Y1_N1END[1]),
    .I1(Tile_X0Y1_N2END[5]),
    .I2(Tile_X0Y1_E1END[1]),
    .I3(Tile_X0Y1_E2END[5]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2692_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2693_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q ),
    .A2(_1010_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2694_ (.I(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2695_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2696_ (.I(_1013_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2697_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(_1014_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2698_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2699_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(_1016_),
    .B(_1015_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q ),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2700_ (.I(_1017_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2701_ (.A1(_1007_),
    .A2(_1012_),
    .B(_1017_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2702_ (.A1(_1008_),
    .A2(_1011_),
    .B(_1018_),
    .C(_0147_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2703_ (.A1(_1007_),
    .A2(_1012_),
    .B(_1017_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2704_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2705_ (.I(_1021_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2706_ (.A1(_0027_),
    .A2(_0147_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2707_ (.A1(Tile_X0Y1_E2MID[4]),
    .A2(_0147_),
    .B(_1023_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2708_ (.I(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2709_ (.A1(_1019_),
    .A2(_1021_),
    .B(_1024_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2710_ (.A1(_1020_),
    .A2(_1022_),
    .B(_1025_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2711_ (.A1(_1019_),
    .A2(_1021_),
    .B(_1024_),
    .C(_0150_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2712_ (.A1(_0149_),
    .A2(_0454_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2713_ (.A1(Tile_X0Y1_W2MID[5]),
    .A2(_0149_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q ),
    .C(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2714_ (.A1(Tile_X0Y1_N2MID[5]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q ),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2715_ (.A1(Tile_X0Y1_E2MID[5]),
    .A2(_0149_),
    .B(_1031_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2716_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q ),
    .A2(_1032_),
    .B(_1030_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2717_ (.A1(_0152_),
    .A2(_1033_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2718_ (.A1(_0152_),
    .A2(_1033_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2719_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2720_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .A2(_1036_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2721_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2722_ (.A1(_0151_),
    .A2(_1038_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2723_ (.I0(Tile_X0Y1_NN4END[3]),
    .I1(Tile_X0Y1_E1END[1]),
    .I2(Tile_X0Y1_E2END[3]),
    .I3(Tile_X0Y1_E6END[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2724_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .A2(_1040_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2725_ (.I0(Tile_X0Y0_S2MID[3]),
    .I1(Tile_X0Y1_W2END[3]),
    .I2(Tile_X0Y0_S4END[7]),
    .I3(Tile_X0Y1_W6END[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2726_ (.A1(_0151_),
    .A2(_1042_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2727_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .A2(_1041_),
    .A3(_1043_),
    .B1(_1037_),
    .B2(_1039_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2728_ (.I0(Tile_X0Y1_NN4END[1]),
    .I1(Tile_X0Y1_EE4END[1]),
    .I2(Tile_X0Y0_S4END[5]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q ),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2729_ (.I0(Tile_X0Y1_N2END[4]),
    .I1(Tile_X0Y1_E2END[4]),
    .I2(Tile_X0Y0_SS4END[6]),
    .I3(Tile_X0Y1_W2END[4]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q ),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2730_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .A2(_1045_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2731_ (.A1(_0150_),
    .A2(_1044_),
    .B(_1046_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q ),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2732_ (.I(_1047_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2733_ (.A1(_1027_),
    .A2(_1035_),
    .B(_1047_),
    .ZN(\Tile_X0Y1_DSP_bot.B2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2734_ (.A1(_1028_),
    .A2(_1034_),
    .B(_1048_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2735_ (.A1(_1027_),
    .A2(_1035_),
    .B(_1047_),
    .C(_0131_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2736_ (.A1(_0131_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[2] ),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2737_ (.I(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2738_ (.A1(_1049_),
    .A2(_1052_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2739_ (.A1(_1050_),
    .A2(_1051_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2740_ (.A1(_0598_),
    .A2(_1053_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2741_ (.I(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2742_ (.A1(_0552_),
    .A2(_0926_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2743_ (.A1(_0552_),
    .A2(_0926_),
    .B(_0722_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2744_ (.A1(_0721_),
    .A2(_0927_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2745_ (.A1(_0723_),
    .A2(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2746_ (.A1(_0722_),
    .A2(_1055_),
    .A3(_1057_),
    .Z(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2747_ (.A1(_0998_),
    .A2(_1061_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2748_ (.A1(_0997_),
    .A2(_1062_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2749_ (.A1(_0935_),
    .A2(_0936_),
    .Z(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2750_ (.A1(_0997_),
    .A2(_1062_),
    .B(_1064_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2751_ (.A1(_1056_),
    .A2(_1058_),
    .B(_1060_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2752_ (.A1(_1063_),
    .A2(_1064_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2753_ (.A1(_1066_),
    .A2(_1067_),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2754_ (.A1(_1065_),
    .A2(_1068_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2755_ (.A1(_1065_),
    .A2(_1068_),
    .B(_0951_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2756_ (.A1(_0942_),
    .A2(_0944_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2757_ (.A1(_0679_),
    .A2(_0824_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2758_ (.A1(_0679_),
    .A2(_0775_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2759_ (.A1(_0940_),
    .A2(_1072_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2760_ (.A1(_0598_),
    .A2(_0882_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2761_ (.A1(_0598_),
    .A2(_0882_),
    .A3(_1074_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2762_ (.A1(_1074_),
    .A2(_1075_),
    .Z(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2763_ (.I(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2764_ (.A1(_1071_),
    .A2(_1078_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2765_ (.A1(_0942_),
    .A2(_0944_),
    .A3(_1077_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2766_ (.A1(_1079_),
    .A2(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2767_ (.A1(_0600_),
    .A2(_0948_),
    .B(_0946_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2768_ (.A1(_1079_),
    .A2(_1080_),
    .A3(_1082_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2769_ (.A1(_1081_),
    .A2(_1082_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2770_ (.A1(_0937_),
    .A2(_0949_),
    .B1(_0950_),
    .B2(_0725_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2771_ (.A1(_1084_),
    .A2(_1085_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2772_ (.A1(_1084_),
    .A2(_1085_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2773_ (.A1(_1070_),
    .A2(_1087_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2774_ (.A1(_1070_),
    .A2(_1087_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2775_ (.A1(_0951_),
    .A2(_1069_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2776_ (.I0(Tile_X0Y1_N2END[6]),
    .I1(Tile_X0Y1_E2END[6]),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q ),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2777_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q ),
    .A2(Tile_X0Y1_W2END[6]),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2778_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q ),
    .A2(_0153_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q ),
    .C(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2779_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q ),
    .A2(_1091_),
    .B(_1093_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2780_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .A2(_0436_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2781_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .A2(_1094_),
    .B(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2782_ (.A1(_0048_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2783_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .B(_1097_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2784_ (.A1(_0032_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2785_ (.A1(Tile_X0Y1_N2MID[7]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .B(_1099_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2786_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .A2(_1100_),
    .B(_1098_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2787_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2788_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2789_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2790_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .A2(_0211_),
    .B(_1104_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2791_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .A2(_1103_),
    .B(_1105_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2792_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ),
    .A2(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2793_ (.A1(_0127_),
    .A2(_1102_),
    .B(_1107_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2794_ (.I0(_0456_),
    .I1(Tile_X0Y0_E1END[3]),
    .I2(Tile_X0Y1_N2MID[7]),
    .I3(Tile_X0Y0_E2END[7]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2795_ (.A1(_0127_),
    .A2(_1109_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2796_ (.I0(Tile_X0Y0_S1END[3]),
    .I1(Tile_X0Y0_W1END[1]),
    .I2(Tile_X0Y0_S2END[7]),
    .I3(Tile_X0Y0_W1END[3]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2797_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(_1111_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2798_ (.A1(_1110_),
    .A2(_1112_),
    .B(_1108_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2799_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2800_ (.A1(Tile_X0Y1_N2MID[6]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2801_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .A2(_1113_),
    .B(_1114_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q ),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2802_ (.I0(Tile_X0Y1_W2MID[6]),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2803_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q ),
    .A2(_1116_),
    .B(_1115_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2804_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q ),
    .A2(_1117_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2805_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q ),
    .A2(_1096_),
    .B1(_1101_),
    .B2(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2806_ (.I(_1119_),
    .ZN(\Tile_X0Y1_DSP_bot.A0 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2807_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[0] ),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2808_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(_1119_),
    .B(_1120_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2809_ (.I(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2810_ (.A1(_0775_),
    .A2(_1121_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2811_ (.A1(_0990_),
    .A2(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2812_ (.A1(_0846_),
    .A2(_0882_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2813_ (.A1(_0990_),
    .A2(_1123_),
    .B1(_1124_),
    .B2(_1125_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2814_ (.A1(_0992_),
    .A2(_0993_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2815_ (.A1(_1126_),
    .A2(_1127_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2816_ (.A1(_1126_),
    .A2(_1127_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2817_ (.A1(_0679_),
    .A2(_1053_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2818_ (.A1(_0552_),
    .A2(_0907_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2819_ (.A1(_0719_),
    .A2(_0720_),
    .A3(_0907_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2820_ (.A1(_1059_),
    .A2(_1131_),
    .Z(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2821_ (.A1(_1130_),
    .A2(_1133_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2822_ (.A1(_1130_),
    .A2(_1133_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2823_ (.A1(_1129_),
    .A2(_1135_),
    .B(_1128_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2824_ (.A1(_0998_),
    .A2(_1061_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2825_ (.A1(_1062_),
    .A2(_1136_),
    .A3(_1137_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2826_ (.A1(_1057_),
    .A2(_1132_),
    .B(_1134_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2827_ (.A1(_0998_),
    .A2(_1061_),
    .A3(_1136_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2828_ (.A1(_1139_),
    .A2(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2829_ (.A1(_1138_),
    .A2(_1141_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2830_ (.I(_1142_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2831_ (.A1(_1066_),
    .A2(_1067_),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2832_ (.A1(_1143_),
    .A2(_1144_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2833_ (.A1(_1090_),
    .A2(_1145_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2834_ (.A1(_1090_),
    .A2(_1145_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2835_ (.A1(_0882_),
    .A2(_1121_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2836_ (.A1(_0990_),
    .A2(_1148_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2837_ (.A1(_1124_),
    .A2(_1125_),
    .Z(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2838_ (.A1(_1149_),
    .A2(_1150_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2839_ (.A1(_0927_),
    .A2(_1053_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2840_ (.A1(_0721_),
    .A2(_0747_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2841_ (.A1(_0551_),
    .A2(_0747_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2842_ (.A1(_0551_),
    .A2(_0747_),
    .A3(_1132_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2843_ (.A1(_0551_),
    .A2(_0747_),
    .B(_1132_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2844_ (.A1(_1132_),
    .A2(_1152_),
    .A3(_1154_),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2845_ (.A1(_1149_),
    .A2(_1150_),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2846_ (.A1(_1151_),
    .A2(_1157_),
    .A3(_1158_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2847_ (.A1(_1151_),
    .A2(_1159_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2848_ (.A1(_1129_),
    .A2(_1135_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2849_ (.A1(_1151_),
    .A2(_1159_),
    .B(_1161_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2850_ (.A1(_0926_),
    .A2(_1054_),
    .A3(_1156_),
    .B(_1155_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2851_ (.I0(Tile_X0Y1_N2END[2]),
    .I1(Tile_X0Y1_E2END[2]),
    .I2(Tile_X0Y0_S2MID[2]),
    .I3(Tile_X0Y1_WW4END[2]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q ),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2852_ (.I0(_0231_),
    .I1(_1164_),
    .S(_0157_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2853_ (.A1(_0375_),
    .A2(_0377_),
    .B(_0410_),
    .C(_0155_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2854_ (.A1(_0632_),
    .A2(_0633_),
    .B(_0654_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2855_ (.A1(_0096_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2856_ (.A1(Tile_X0Y0_S2MID[5]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .C(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2857_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_1169_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2858_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .A2(_1166_),
    .A3(_1167_),
    .B(_1170_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2859_ (.I0(Tile_X0Y1_N1END[1]),
    .I1(Tile_X0Y1_N2END[5]),
    .I2(Tile_X0Y1_E1END[1]),
    .I3(Tile_X0Y1_E2END[5]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2860_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2861_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ),
    .A2(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2862_ (.A1(_1171_),
    .A2(_1174_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2863_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2864_ (.I(_1176_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2865_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_1177_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2866_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2867_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_1179_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2868_ (.A1(_0156_),
    .A2(_1180_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2869_ (.A1(_1178_),
    .A2(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2870_ (.A1(_1175_),
    .A2(_1182_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2871_ (.A1(_1171_),
    .A2(_1174_),
    .B1(_1178_),
    .B2(_1181_),
    .C(_0154_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2872_ (.A1(Tile_X0Y1_W2MID[2]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2873_ (.A1(Tile_X0Y1_N2MID[2]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2874_ (.A1(Tile_X0Y1_E2MID[2]),
    .A2(_0154_),
    .B(_1185_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2875_ (.A1(_1183_),
    .A2(_1184_),
    .B1(_1186_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ),
    .C(_0157_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2876_ (.I0(Tile_X0Y1_N2MID[3]),
    .I1(Tile_X0Y1_E2MID[3]),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .I3(Tile_X0Y1_W2MID[3]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q ),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2877_ (.A1(_0157_),
    .A2(_1188_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2878_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ),
    .A2(_1189_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2879_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ),
    .A2(_1165_),
    .B1(_1187_),
    .B2(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2880_ (.I(_1191_),
    .ZN(\Tile_X0Y1_DSP_bot.B1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2881_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ),
    .A2(_1165_),
    .B1(_1187_),
    .B2(_1190_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2882_ (.A1(_0131_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[1] ),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2883_ (.A1(_1192_),
    .A2(_1193_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2884_ (.A1(_0599_),
    .A2(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2885_ (.A1(_1163_),
    .A2(_1195_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2886_ (.A1(_1163_),
    .A2(_1195_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2887_ (.A1(_1151_),
    .A2(_1159_),
    .A3(_1161_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2888_ (.A1(_1197_),
    .A2(_1198_),
    .B(_1162_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2889_ (.I(_1199_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2890_ (.A1(_1139_),
    .A2(_1140_),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2891_ (.A1(_1200_),
    .A2(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2892_ (.A1(_1199_),
    .A2(_1201_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2893_ (.A1(_1196_),
    .A2(_1203_),
    .B(_1202_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2894_ (.A1(_1143_),
    .A2(_1144_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2895_ (.A1(_1204_),
    .A2(_1205_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2896_ (.A1(_1204_),
    .A2(_1205_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2897_ (.A1(_0882_),
    .A2(_0988_),
    .B1(_1121_),
    .B2(_0824_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2898_ (.A1(_1149_),
    .A2(_1208_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2899_ (.A1(_0907_),
    .A2(_1054_),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2900_ (.A1(_0552_),
    .A2(_0847_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2901_ (.A1(_0721_),
    .A2(_0747_),
    .B(_1211_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2902_ (.A1(_0719_),
    .A2(_0720_),
    .A3(_0847_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2903_ (.A1(_0551_),
    .A2(_0747_),
    .A3(_1213_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2904_ (.A1(_1153_),
    .A2(_1210_),
    .A3(_1211_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2905_ (.A1(_1209_),
    .A2(_1215_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2906_ (.A1(_1149_),
    .A2(_1150_),
    .A3(_1157_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2907_ (.A1(_1216_),
    .A2(_1217_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2908_ (.A1(_1216_),
    .A2(_1217_),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2909_ (.A1(_0680_),
    .A2(_1194_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2910_ (.A1(_1210_),
    .A2(_1212_),
    .B(_1214_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2911_ (.I0(Tile_X0Y1_NN4END[3]),
    .I1(Tile_X0Y1_E2END[6]),
    .I2(Tile_X0Y0_S2MID[6]),
    .I3(Tile_X0Y1_W2END[6]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q ),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2912_ (.I0(Tile_X0Y1_E2END[3]),
    .I1(Tile_X0Y1_WW4END[2]),
    .I2(Tile_X0Y0_SS4END[7]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2913_ (.I0(_1222_),
    .I1(_1223_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2914_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ),
    .A2(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2915_ (.A1(_0667_),
    .A2(_0670_),
    .B(_0158_),
    .C(_0621_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2916_ (.A1(_0666_),
    .A2(_0671_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .C(_0622_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2917_ (.A1(Tile_X0Y1_W2MID[6]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2918_ (.I(_1228_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2919_ (.A1(Tile_X0Y1_E2MID[6]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2920_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .A2(_1113_),
    .B(_1230_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2921_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2922_ (.A1(_1227_),
    .A2(_1229_),
    .B(_1231_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2923_ (.A1(_1226_),
    .A2(_1228_),
    .B(_1232_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2924_ (.I0(Tile_X0Y1_N2MID[7]),
    .I1(Tile_X0Y1_E2MID[7]),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .I3(Tile_X0Y1_W2MID[7]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q ),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2925_ (.A1(_0159_),
    .A2(_1235_),
    .B(_0160_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2926_ (.I(_1236_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2927_ (.A1(_1233_),
    .A2(_1236_),
    .B(_1225_),
    .ZN(\Tile_X0Y1_DSP_bot.B0 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2928_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ),
    .A2(_1224_),
    .B1(_1234_),
    .B2(_1237_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2929_ (.A1(_1233_),
    .A2(_1236_),
    .B(_0131_),
    .C(_1225_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2930_ (.A1(_0131_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[0] ),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2931_ (.I(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2932_ (.A1(_1238_),
    .A2(_1241_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2933_ (.A1(_0598_),
    .A2(_1242_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2934_ (.A1(_0598_),
    .A2(_1221_),
    .A3(_1242_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2935_ (.I(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2936_ (.A1(_1221_),
    .A2(_1243_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2937_ (.A1(_1220_),
    .A2(_1246_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2938_ (.A1(_1219_),
    .A2(_1247_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2939_ (.A1(_1218_),
    .A2(_1248_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2940_ (.A1(_1160_),
    .A2(_1161_),
    .A3(_1197_),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2941_ (.I(_1250_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2942_ (.A1(_1249_),
    .A2(_1251_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2943_ (.A1(_1220_),
    .A2(_1246_),
    .B(_1245_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2944_ (.A1(_1249_),
    .A2(_1250_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2945_ (.A1(_1253_),
    .A2(_1254_),
    .B(_1252_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2946_ (.A1(_1196_),
    .A2(_1203_),
    .Z(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2947_ (.A1(_1255_),
    .A2(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2948_ (.A1(_0747_),
    .A2(_1050_),
    .A3(_1051_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2949_ (.A1(_0552_),
    .A2(_0989_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2950_ (.A1(_1213_),
    .A2(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2951_ (.A1(_1213_),
    .A2(_1259_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2952_ (.A1(_1213_),
    .A2(_1258_),
    .A3(_1259_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2953_ (.A1(_0882_),
    .A2(_1121_),
    .A3(_1262_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2954_ (.A1(_1209_),
    .A2(_1215_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2955_ (.A1(_1263_),
    .A2(_1264_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2956_ (.A1(_1209_),
    .A2(_1215_),
    .A3(_1263_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2957_ (.A1(_0926_),
    .A2(_1194_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2958_ (.A1(_1258_),
    .A2(_1260_),
    .B(_1261_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2959_ (.A1(_0679_),
    .A2(_1242_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2960_ (.A1(_0679_),
    .A2(_1242_),
    .A3(_1268_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2961_ (.A1(_1268_),
    .A2(_1269_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2962_ (.A1(_1267_),
    .A2(_1268_),
    .A3(_1269_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2963_ (.A1(_1266_),
    .A2(_1272_),
    .B(_1265_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2964_ (.A1(_1219_),
    .A2(_1247_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2965_ (.A1(_1267_),
    .A2(_1271_),
    .B(_1270_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2966_ (.A1(_1273_),
    .A2(_1274_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2967_ (.A1(_1275_),
    .A2(_1276_),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2968_ (.A1(_1273_),
    .A2(_1274_),
    .B(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2969_ (.A1(_1253_),
    .A2(_1254_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2970_ (.A1(_1278_),
    .A2(_1279_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2971_ (.A1(_1148_),
    .A2(_1262_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2972_ (.A1(_0719_),
    .A2(_0720_),
    .A3(_1122_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2973_ (.A1(_0552_),
    .A2(_1122_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2974_ (.A1(_1259_),
    .A2(_1282_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2975_ (.A1(_0719_),
    .A2(_0720_),
    .A3(_0989_),
    .B(_1283_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2976_ (.A1(_0719_),
    .A2(_0720_),
    .A3(_0989_),
    .A4(_1283_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2977_ (.A1(_0846_),
    .A2(_1050_),
    .A3(_1051_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2978_ (.A1(_1285_),
    .A2(_1286_),
    .B(_1287_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2979_ (.A1(_0926_),
    .A2(_1238_),
    .A3(_1241_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2980_ (.A1(_1284_),
    .A2(_1288_),
    .B(_1289_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2981_ (.A1(_1284_),
    .A2(_1288_),
    .A3(_1289_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2982_ (.A1(_1290_),
    .A2(_1291_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2983_ (.A1(_0907_),
    .A2(_1194_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2984_ (.A1(_1290_),
    .A2(_1291_),
    .A3(_1293_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2985_ (.A1(_1292_),
    .A2(_1293_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2986_ (.A1(_1290_),
    .A2(_1291_),
    .B(_1293_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2987_ (.A1(_1281_),
    .A2(_1294_),
    .A3(_1296_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2988_ (.A1(_1266_),
    .A2(_1272_),
    .Z(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2989_ (.A1(_1297_),
    .A2(_1298_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2990_ (.A1(_1290_),
    .A2(_1295_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2991_ (.A1(_1297_),
    .A2(_1298_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2992_ (.A1(_1300_),
    .A2(_1301_),
    .B(_1299_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2993_ (.A1(_1275_),
    .A2(_1276_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2994_ (.A1(_1277_),
    .A2(_1302_),
    .A3(_1303_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2995_ (.A1(_0748_),
    .A2(_1194_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2996_ (.A1(_1049_),
    .A2(_1052_),
    .A3(_1122_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2997_ (.A1(_0989_),
    .A2(_1049_),
    .A3(_1052_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2998_ (.A1(_1282_),
    .A2(_1307_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2999_ (.A1(_0907_),
    .A2(_1238_),
    .A3(_1241_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3000_ (.A1(_1308_),
    .A2(_1309_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3001_ (.A1(_1308_),
    .A2(_1309_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3002_ (.A1(_1305_),
    .A2(_1308_),
    .A3(_1309_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3003_ (.A1(_1285_),
    .A2(_1286_),
    .A3(_1287_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3004_ (.A1(_1288_),
    .A2(_1313_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3005_ (.A1(_1312_),
    .A2(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3006_ (.A1(_1281_),
    .A2(_1292_),
    .A3(_1293_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3007_ (.A1(_1315_),
    .A2(_1316_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3008_ (.A1(_1305_),
    .A2(_1311_),
    .B(_1310_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3009_ (.A1(_1315_),
    .A2(_1316_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3010_ (.A1(_1318_),
    .A2(_1319_),
    .B(_1317_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3011_ (.A1(_1300_),
    .A2(_1301_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3012_ (.A1(_1320_),
    .A2(_1321_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3013_ (.A1(_1282_),
    .A2(_1307_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3014_ (.A1(_1282_),
    .A2(_1307_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3015_ (.A1(_0846_),
    .A2(_1239_),
    .A3(_1240_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3016_ (.A1(_0747_),
    .A2(_1239_),
    .A3(_1240_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3017_ (.A1(_0847_),
    .A2(_1192_),
    .A3(_1193_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3018_ (.A1(_1326_),
    .A2(_1327_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3019_ (.A1(_1326_),
    .A2(_1327_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3020_ (.A1(_1308_),
    .A2(_1323_),
    .A3(_1329_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3021_ (.A1(_1312_),
    .A2(_1314_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3022_ (.A1(_1312_),
    .A2(_1314_),
    .A3(_1330_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3023_ (.A1(_1328_),
    .A2(_1330_),
    .B(_1331_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3024_ (.A1(_1315_),
    .A2(_1316_),
    .A3(_1318_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3025_ (.A1(_1333_),
    .A2(_1334_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3026_ (.A1(_1333_),
    .A2(_1334_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3027_ (.A1(_1324_),
    .A2(_1329_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3028_ (.A1(_0988_),
    .A2(_1239_),
    .A3(_1240_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3029_ (.A1(_0989_),
    .A2(_1192_),
    .A3(_1193_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3030_ (.A1(_1327_),
    .A2(_1338_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _3031_ (.A1(_0989_),
    .A2(_1192_),
    .A3(_1193_),
    .B1(_1238_),
    .B2(_1241_),
    .B3(_0847_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3032_ (.A1(_1327_),
    .A2(_1338_),
    .B(_1341_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3033_ (.A1(_1054_),
    .A2(_1122_),
    .A3(_1342_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3034_ (.A1(_1327_),
    .A2(_1338_),
    .B(_1341_),
    .C(_1306_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3035_ (.A1(_1324_),
    .A2(_1329_),
    .A3(_1344_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3036_ (.A1(_1340_),
    .A2(_1343_),
    .B(_1337_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3037_ (.I(_1346_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3038_ (.A1(_1328_),
    .A2(_1332_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3039_ (.A1(_1347_),
    .A2(_1348_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3040_ (.A1(_1347_),
    .A2(_1348_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3041_ (.A1(_1340_),
    .A2(_1345_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3042_ (.A1(_1121_),
    .A2(_1242_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3043_ (.A1(_1122_),
    .A2(_1192_),
    .A3(_1193_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3044_ (.A1(_1122_),
    .A2(_1194_),
    .A3(_1338_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3045_ (.A1(_1306_),
    .A2(_1325_),
    .A3(_1339_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3046_ (.A1(_1122_),
    .A2(_1194_),
    .A3(_1338_),
    .A4(_1355_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3047_ (.A1(_1351_),
    .A2(_1356_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3048_ (.I(_1357_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3049_ (.A1(_1347_),
    .A2(_1348_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3050_ (.A1(_1347_),
    .A2(_1348_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3051_ (.A1(_1357_),
    .A2(_1360_),
    .B(_1349_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3052_ (.A1(_1358_),
    .A2(_1359_),
    .B(_1350_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3053_ (.A1(_1333_),
    .A2(_1334_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3054_ (.A1(_1333_),
    .A2(_1334_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3055_ (.A1(_1362_),
    .A2(_1364_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3056_ (.A1(_1362_),
    .A2(_1364_),
    .B(_1335_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3057_ (.A1(_1361_),
    .A2(_1363_),
    .B(_1336_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3058_ (.A1(_1320_),
    .A2(_1321_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3059_ (.A1(_1367_),
    .A2(_1368_),
    .B(_1322_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3060_ (.A1(_1275_),
    .A2(_1276_),
    .A3(_1302_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3061_ (.A1(_1369_),
    .A2(_1370_),
    .B(_1304_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3062_ (.A1(_1278_),
    .A2(_1279_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3063_ (.A1(_1371_),
    .A2(_1372_),
    .B(_1280_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3064_ (.A1(_1255_),
    .A2(_1256_),
    .B1(_1371_),
    .B2(_1372_),
    .C(_1280_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3065_ (.A1(_1257_),
    .A2(_1374_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3066_ (.A1(_1207_),
    .A2(_1257_),
    .A3(_1374_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3067_ (.A1(_1207_),
    .A2(_1257_),
    .A3(_1374_),
    .B(_1206_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3068_ (.A1(_1146_),
    .A2(_1377_),
    .B(_1147_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3069_ (.A1(_1089_),
    .A2(_1378_),
    .B(_1088_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3070_ (.A1(_1083_),
    .A2(_1086_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3071_ (.A1(_0940_),
    .A2(_1072_),
    .B(_1076_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3072_ (.A1(_0598_),
    .A2(_0824_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3073_ (.A1(_1073_),
    .A2(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3074_ (.A1(_1381_),
    .A2(_1383_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3075_ (.A1(_1071_),
    .A2(_1078_),
    .A3(_1384_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3076_ (.A1(_1079_),
    .A2(_1384_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3077_ (.A1(_1380_),
    .A2(_1386_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3078_ (.A1(_1086_),
    .A2(_1386_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3079_ (.A1(_1379_),
    .A2(_1387_),
    .B(_1388_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3080_ (.A1(_1079_),
    .A2(_1080_),
    .A3(_1082_),
    .A4(_1384_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3081_ (.A1(_0598_),
    .A2(_0775_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3082_ (.A1(_0679_),
    .A2(_0824_),
    .B(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3083_ (.A1(_1381_),
    .A2(_1383_),
    .B(_1385_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3084_ (.A1(_1392_),
    .A2(_1393_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3085_ (.A1(_1390_),
    .A2(_1394_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3086_ (.A1(_1390_),
    .A2(_1394_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3087_ (.A1(_1395_),
    .A2(_1396_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3088_ (.A1(_1389_),
    .A2(_1397_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3089_ (.A1(_0529_),
    .A2(_1398_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3090_ (.A1(_0529_),
    .A2(_1389_),
    .A3(_1397_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3091_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .I1(Tile_X0Y0_S2MID[1]),
    .I2(Tile_X0Y0_E2MID[1]),
    .I3(Tile_X0Y0_W2MID[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q ),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3092_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3093_ (.A1(_0124_),
    .A2(_1402_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3094_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3095_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ),
    .A2(_1404_),
    .B(_0125_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3096_ (.I0(Tile_X0Y0_S1END[0]),
    .I1(Tile_X0Y0_S1END[2]),
    .I2(Tile_X0Y0_S2END[6]),
    .I3(Tile_X0Y0_W1END[2]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3097_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ),
    .A2(_1406_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3098_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .I1(Tile_X0Y0_E1END[2]),
    .I2(Tile_X0Y1_N2MID[6]),
    .I3(Tile_X0Y0_E2END[6]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3099_ (.A1(_0124_),
    .A2(_1408_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3100_ (.A1(_1403_),
    .A2(_1405_),
    .B1(_1407_),
    .B2(_1409_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3101_ (.I0(Tile_X0Y1_NN4END[6]),
    .I1(Tile_X0Y0_E2END[1]),
    .I2(Tile_X0Y0_S2END[1]),
    .I3(Tile_X0Y0_W2END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q ),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3102_ (.I0(Tile_X0Y0_E2MID[0]),
    .I1(Tile_X0Y0_W2MID[0]),
    .I2(Tile_X0Y0_S2MID[0]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q ),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3103_ (.I0(Tile_X0Y0_EE4END[3]),
    .I1(Tile_X0Y0_WW4END[1]),
    .I2(Tile_X0Y0_S4END[0]),
    .I3(_0561_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q ),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3104_ (.I0(_1411_),
    .I1(_1410_),
    .I2(_1401_),
    .I3(_1412_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3105_ (.A1(_0162_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3106_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[13] ),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3107_ (.A1(_0163_),
    .A2(_1414_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3108_ (.A1(_0163_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[13] ),
    .B1(_1413_),
    .B2(_1415_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3109_ (.A1(_1379_),
    .A2(_1387_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3110_ (.A1(_1416_),
    .A2(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3111_ (.I0(Tile_X0Y1_N2MID[5]),
    .I1(Tile_X0Y0_SS4END[1]),
    .I2(Tile_X0Y0_E2END[5]),
    .I3(Tile_X0Y0_W2END[5]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q ),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3112_ (.I0(_0672_),
    .I1(_0104_),
    .I2(_0039_),
    .I3(_0454_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q ),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3113_ (.I(_1420_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3114_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .I1(Tile_X0Y0_S2MID[5]),
    .I2(Tile_X0Y0_E2MID[5]),
    .I3(Tile_X0Y0_W2MID[5]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q ),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3115_ (.I0(_1421_),
    .I1(_1422_),
    .I2(_1419_),
    .I3(_0653_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3116_ (.A1(_0162_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3117_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[12] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3118_ (.A1(_0161_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .B1(_1423_),
    .B2(_1424_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3119_ (.A1(_1089_),
    .A2(_1378_),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3120_ (.A1(_1425_),
    .A2(_1426_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3121_ (.A1(_0163_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[11] ),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3122_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .I1(Tile_X0Y0_E2MID[3]),
    .I2(Tile_X0Y0_S2MID[3]),
    .I3(Tile_X0Y0_W2MID[3]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q ),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3123_ (.I(_1429_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3124_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3125_ (.A1(_0122_),
    .A2(_1431_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3126_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3127_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ),
    .A2(_1433_),
    .B(_0123_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3128_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .I1(Tile_X0Y0_E1END[2]),
    .I2(Tile_X0Y1_N2MID[6]),
    .I3(Tile_X0Y0_E2END[6]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ),
    .Z(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3129_ (.A1(_0122_),
    .A2(_1435_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3130_ (.I0(Tile_X0Y0_S1END[0]),
    .I1(Tile_X0Y0_S1END[2]),
    .I2(Tile_X0Y0_S2END[6]),
    .I3(Tile_X0Y0_W1END[2]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3131_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ),
    .A2(_1437_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3132_ (.A1(_1432_),
    .A2(_1434_),
    .B1(_1436_),
    .B2(_1438_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3133_ (.A1(Tile_X0Y1_N2MID[3]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q ),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3134_ (.A1(_0057_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q ),
    .C(_1439_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3135_ (.I0(Tile_X0Y0_S2END[3]),
    .I1(Tile_X0Y0_WW4END[1]),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q ),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3136_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q ),
    .A2(_1441_),
    .B(_1440_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3137_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .I1(Tile_X0Y0_E2MID[2]),
    .I2(Tile_X0Y0_S2MID[2]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q ),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3138_ (.I0(_1443_),
    .I1(_1429_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3139_ (.I0(Tile_X0Y1_NN4END[6]),
    .I1(Tile_X0Y0_S4END[2]),
    .I2(Tile_X0Y0_E2END[2]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q ),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3140_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ),
    .A2(_1445_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3141_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ),
    .A2(_1442_),
    .B(_1446_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q ),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3142_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q ),
    .A2(_1444_),
    .B(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3143_ (.I(_1448_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3144_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(_1448_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3145_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[11] ),
    .B(_1449_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3146_ (.A1(_1428_),
    .A2(_1450_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3147_ (.A1(_1090_),
    .A2(_1145_),
    .A3(_1377_),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3148_ (.A1(_1451_),
    .A2(_1452_),
    .Z(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3149_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3150_ (.A1(_0059_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q ),
    .C(_1454_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3151_ (.A1(Tile_X0Y1_N4END[7]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3152_ (.A1(_0057_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ),
    .B(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3153_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q ),
    .A2(_1457_),
    .B(_1455_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3154_ (.I0(Tile_X0Y1_N2MID[7]),
    .I1(Tile_X0Y0_EE4END[2]),
    .I2(Tile_X0Y0_S2END[7]),
    .I3(Tile_X0Y0_W2END[7]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q ),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3155_ (.I(_1459_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3156_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q ),
    .A2(_1458_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3157_ (.A1(_0121_),
    .A2(_1459_),
    .B(_1461_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3158_ (.A1(Tile_X0Y0_E2MID[6]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q ),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3159_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ),
    .A2(_0421_),
    .B(_1463_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3160_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3161_ (.A1(_0119_),
    .A2(_1465_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3162_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .Z(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3163_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ),
    .A2(_1467_),
    .B(_0120_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3164_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .I1(Tile_X0Y0_E1END[2]),
    .I2(Tile_X0Y1_N2MID[6]),
    .I3(Tile_X0Y0_E2END[6]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .Z(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3165_ (.A1(_0119_),
    .A2(_1469_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3166_ (.I0(Tile_X0Y0_S1END[2]),
    .I1(Tile_X0Y0_S2END[6]),
    .I2(Tile_X0Y0_W1END[0]),
    .I3(Tile_X0Y0_W1END[2]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3167_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ),
    .A2(_1471_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3168_ (.A1(_1466_),
    .A2(_1468_),
    .B1(_1470_),
    .B2(_1472_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3169_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3170_ (.A1(_0097_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q ),
    .C(_1473_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3171_ (.A1(_0121_),
    .A2(_1464_),
    .A3(_1474_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3172_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ),
    .A2(_0630_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q ),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3173_ (.A1(_1475_),
    .A2(_1476_),
    .B(_1462_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3174_ (.A1(_0162_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3175_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[10] ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3176_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .A2(_0164_),
    .B1(_1477_),
    .B2(_1478_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3177_ (.A1(_1257_),
    .A2(_1374_),
    .B(_1207_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3178_ (.A1(_1376_),
    .A2(_1479_),
    .A3(_1480_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3179_ (.A1(_1207_),
    .A2(_1375_),
    .A3(_1479_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3180_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .Z(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3181_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3182_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_1483_),
    .Z(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3183_ (.A1(_0165_),
    .A2(_1484_),
    .B(_1485_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3184_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0351_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3185_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0488_),
    .B(_1487_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3186_ (.A1(Tile_X0Y1_WW4END[0]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3187_ (.A1(_0140_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .C(_1489_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3188_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_1488_),
    .A3(_1490_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3189_ (.I0(Tile_X0Y1_N1END[0]),
    .I1(Tile_X0Y1_E1END[0]),
    .I2(Tile_X0Y1_N2END[0]),
    .I3(Tile_X0Y1_E2END[0]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3190_ (.A1(_0165_),
    .A2(_1492_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q ),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3191_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q ),
    .A2(_1486_),
    .B1(_1491_),
    .B2(_1493_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3192_ (.I0(_0489_),
    .I1(_0351_),
    .I2(Tile_X0Y0_S2MID[6]),
    .I3(Tile_X0Y1_W1END[2]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .Z(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3193_ (.I0(Tile_X0Y1_N1END[2]),
    .I1(Tile_X0Y1_E1END[2]),
    .I2(Tile_X0Y1_N2END[6]),
    .I3(Tile_X0Y1_E2END[6]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3194_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .Z(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3195_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .Z(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3196_ (.I0(_1495_),
    .I1(_1497_),
    .I2(_1494_),
    .I3(_1496_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3197_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .A2(_0351_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3198_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .A2(_0488_),
    .B(_1498_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3199_ (.A1(Tile_X0Y1_W1END[2]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3200_ (.A1(_0083_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .C(_1500_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3201_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .A2(_1499_),
    .B(_1501_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3202_ (.I0(Tile_X0Y1_N1END[2]),
    .I1(Tile_X0Y1_E1END[2]),
    .I2(Tile_X0Y1_N2END[6]),
    .I3(Tile_X0Y1_E2END[6]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3203_ (.A1(_0170_),
    .A2(_1503_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3204_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .A2(_0207_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3205_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .B(_1505_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3206_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3207_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .A2(_1507_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3208_ (.A1(_0169_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .B(_1508_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3209_ (.A1(_0169_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3210_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3211_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .A2(_0212_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3212_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .B(_1512_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3213_ (.A1(_1510_),
    .A2(_1511_),
    .B1(_1513_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3214_ (.A1(_0170_),
    .A2(_1506_),
    .A3(_1509_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3215_ (.A1(_1514_),
    .A2(_1515_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3216_ (.A1(_1502_),
    .A2(_1504_),
    .B(_1516_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3217_ (.I0(_0489_),
    .I1(_0351_),
    .I2(Tile_X0Y0_S2MID[0]),
    .I3(Tile_X0Y1_W1END[0]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3218_ (.I0(Tile_X0Y1_N1END[0]),
    .I1(Tile_X0Y1_E1END[0]),
    .I2(Tile_X0Y1_N2END[0]),
    .I3(Tile_X0Y1_E2END[0]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3219_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3220_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3221_ (.I0(_1518_),
    .I1(_1519_),
    .I2(_1517_),
    .I3(_1520_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ),
    .Z(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3222_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3223_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .Z(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3224_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(_1523_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3225_ (.A1(_0166_),
    .A2(_1522_),
    .B(_0167_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3226_ (.I0(_0351_),
    .I1(Tile_X0Y0_S2MID[6]),
    .I2(Tile_X0Y1_W1END[0]),
    .I3(Tile_X0Y1_W1END[2]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3227_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(_1526_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3228_ (.I0(Tile_X0Y1_N1END[2]),
    .I1(Tile_X0Y1_E1END[2]),
    .I2(Tile_X0Y1_N2END[6]),
    .I3(Tile_X0Y1_E2END[6]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3229_ (.A1(_0166_),
    .A2(_1528_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3230_ (.A1(_1524_),
    .A2(_1525_),
    .B1(_1527_),
    .B2(_1529_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3231_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3232_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3233_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .A2(_1530_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3234_ (.A1(_0168_),
    .A2(_1531_),
    .B(_1532_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3235_ (.A1(Tile_X0Y0_S2MID[0]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3236_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .A2(_0488_),
    .B(_1534_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3237_ (.A1(Tile_X0Y1_W1END[2]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3238_ (.A1(_0060_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .C(_1536_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3239_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .A2(_1535_),
    .A3(_1537_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3240_ (.I0(Tile_X0Y1_N1END[0]),
    .I1(Tile_X0Y1_E1END[0]),
    .I2(Tile_X0Y1_N2END[0]),
    .I3(Tile_X0Y1_E2END[0]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .Z(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3241_ (.A1(_0168_),
    .A2(_1539_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3242_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .A2(_1533_),
    .B1(_1538_),
    .B2(_1540_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3243_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 ),
    .I3(_1521_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3244_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .Z(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3245_ (.I(_1542_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3246_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q ),
    .A2(_1543_),
    .ZN(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3247_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q ),
    .A2(_1541_),
    .B(_1544_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3248_ (.I(_1545_),
    .ZN(\Tile_X0Y1_DSP_bot.C9 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3249_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[9] ),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3250_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(_1545_),
    .B(_1546_),
    .C(_0163_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3251_ (.A1(_0163_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[9] ),
    .B(_1547_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3252_ (.I(_1548_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3253_ (.A1(_1255_),
    .A2(_1256_),
    .A3(_1373_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3254_ (.A1(_1549_),
    .A2(_1550_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3255_ (.A1(_0163_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[8] ),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3256_ (.A1(_0177_),
    .A2(_0693_),
    .B(_0171_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3257_ (.A1(_0177_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ),
    .B(_1553_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3258_ (.A1(_0172_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3259_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3260_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(_0212_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3261_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .B(_1557_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3262_ (.A1(_1555_),
    .A2(_1556_),
    .B1(_1558_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3263_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3264_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .A2(_1560_),
    .B(_1559_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3265_ (.I0(_0412_),
    .I1(_0657_),
    .I2(Tile_X0Y1_W1END[3]),
    .I3(Tile_X0Y0_S2MID[7]),
    .S0(_0172_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3266_ (.A1(Tile_X0Y1_N1END[3]),
    .A2(_0172_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3267_ (.A1(Tile_X0Y1_N2END[7]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3268_ (.A1(Tile_X0Y1_E2END[7]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3269_ (.A1(Tile_X0Y1_E1END[3]),
    .A2(_0172_),
    .B(_1565_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3270_ (.A1(_1563_),
    .A2(_1564_),
    .B1(_1566_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3271_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .A2(_1562_),
    .B(_1567_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3272_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ),
    .A2(_1561_),
    .B(_1568_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3273_ (.A1(_0177_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3274_ (.I0(_0657_),
    .I1(_0412_),
    .I2(Tile_X0Y0_S2MID[7]),
    .I3(Tile_X0Y1_W1END[3]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .Z(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3275_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .A2(_1570_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3276_ (.I0(Tile_X0Y1_N1END[3]),
    .I1(Tile_X0Y1_N2END[7]),
    .I2(Tile_X0Y1_E1END[3]),
    .I3(Tile_X0Y1_E2END[7]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3277_ (.A1(_0175_),
    .A2(_1572_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3278_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .Z(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3279_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3280_ (.A1(_0175_),
    .A2(_1575_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3281_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .A2(_1574_),
    .B(_0176_),
    .ZN(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3282_ (.A1(_1571_),
    .A2(_1573_),
    .B1(_1576_),
    .B2(_1577_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3283_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 ),
    .ZN(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3284_ (.A1(_0177_),
    .A2(_1578_),
    .B(_1569_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3285_ (.A1(_0171_),
    .A2(_1579_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3286_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(_0672_),
    .B(_0171_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3287_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ),
    .B(_1581_),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3288_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3289_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3290_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(_1584_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3291_ (.A1(_0173_),
    .A2(_1583_),
    .B(_0174_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3292_ (.I0(_0412_),
    .I1(Tile_X0Y1_W1END[1]),
    .I2(Tile_X0Y0_S2MID[7]),
    .I3(Tile_X0Y1_W1END[3]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3293_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(_1587_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3294_ (.I0(Tile_X0Y1_N1END[3]),
    .I1(Tile_X0Y1_N2END[7]),
    .I2(Tile_X0Y1_E1END[3]),
    .I3(Tile_X0Y1_E2END[7]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3295_ (.A1(_0173_),
    .A2(_1589_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3296_ (.A1(_1585_),
    .A2(_1586_),
    .B1(_1588_),
    .B2(_1590_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3297_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(_0421_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3298_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ),
    .B(_1591_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3299_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ),
    .A2(_1582_),
    .A3(_1592_),
    .B1(_1554_),
    .B2(_1580_),
    .ZN(\Tile_X0Y1_DSP_bot.C8 ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3300_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[8] ),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3301_ (.A1(_0162_),
    .A2(\Tile_X0Y1_DSP_bot.C8 ),
    .B(_1593_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .ZN(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3302_ (.A1(_1552_),
    .A2(_1594_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3303_ (.A1(_1371_),
    .A2(_1372_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3304_ (.A1(_1595_),
    .A2(_1596_),
    .Z(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3305_ (.A1(_0163_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[7] ),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3306_ (.A1(Tile_X0Y1_NN4END[0]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3307_ (.A1(_0022_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .C(_1599_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3308_ (.A1(Tile_X0Y1_W2END[0]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3309_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .A2(_0693_),
    .B(_1601_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3310_ (.A1(_1600_),
    .A2(_1602_),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3311_ (.I(_1603_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3312_ (.I0(Tile_X0Y1_N2END[1]),
    .I1(Tile_X0Y1_EE4END[3]),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q ),
    .Z(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3313_ (.A1(Tile_X0Y1_W2END[1]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q ),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3314_ (.A1(_0025_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q ),
    .C(_1606_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3315_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q ),
    .A2(_1605_),
    .B(_1607_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3316_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(_1608_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3317_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(_1604_),
    .B(_1609_),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3318_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .A2(_1578_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3319_ (.A1(Tile_X0Y1_W2MID[0]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .B(_1611_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3320_ (.A1(Tile_X0Y1_E2MID[0]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3321_ (.A1(_0046_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .B(_1613_),
    .ZN(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3322_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .A2(_1612_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3323_ (.I0(Tile_X0Y1_N2MID[1]),
    .I1(Tile_X0Y1_E2MID[1]),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .I3(Tile_X0Y1_W2MID[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q ),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3324_ (.A1(_1614_),
    .A2(_1615_),
    .B1(_1616_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3325_ (.A1(_1610_),
    .A2(_1617_),
    .ZN(\Tile_X0Y1_DSP_bot.C7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3326_ (.I0(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[7] ),
    .I1(\Tile_X0Y1_DSP_bot.C7 ),
    .S(_0162_),
    .Z(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3327_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .A2(_1618_),
    .B(_1598_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3328_ (.I(_1619_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3329_ (.A1(_1369_),
    .A2(_1370_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3330_ (.A1(_1620_),
    .A2(_1621_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3331_ (.I0(Tile_X0Y1_E6END[1]),
    .I1(Tile_X0Y0_S4END[5]),
    .I2(Tile_X0Y1_WW4END[3]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .Z(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3332_ (.I(_1623_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3333_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_1624_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3334_ (.I0(Tile_X0Y1_NN4END[1]),
    .I1(Tile_X0Y1_E2END[5]),
    .I2(Tile_X0Y0_S2MID[5]),
    .I3(Tile_X0Y1_W2END[5]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q ),
    .Z(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3335_ (.I(_1626_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3336_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_1626_),
    .B(_1625_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q ),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3337_ (.I0(Tile_X0Y1_E2MID[4]),
    .I1(Tile_X0Y1_W2MID[4]),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q ),
    .Z(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3338_ (.I0(Tile_X0Y1_N2MID[5]),
    .I1(Tile_X0Y1_E2MID[5]),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3339_ (.A1(Tile_X0Y1_W2MID[5]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3340_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .A2(_0454_),
    .B(_1631_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q ),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3341_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q ),
    .A2(_1630_),
    .B(_1632_),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3342_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_1633_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q ),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3343_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_1629_),
    .B(_1634_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3344_ (.A1(_1628_),
    .A2(_1635_),
    .ZN(\Tile_X0Y1_DSP_bot.C6 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3345_ (.A1(_1628_),
    .A2(_1635_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3346_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[6] ),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3347_ (.A1(_0163_),
    .A2(_1637_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3348_ (.A1(_0163_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[6] ),
    .B1(_1636_),
    .B2(_1638_),
    .ZN(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3349_ (.A1(_1366_),
    .A2(_1368_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3350_ (.A1(_1639_),
    .A2(_1640_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3351_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3352_ (.A1(_0023_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .C(_1642_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3353_ (.I0(Tile_X0Y1_N4END[2]),
    .I1(Tile_X0Y0_SS4END[6]),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3354_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_1644_),
    .B(_1643_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3355_ (.I0(Tile_X0Y1_N2END[3]),
    .I1(Tile_X0Y1_E2END[3]),
    .I2(Tile_X0Y0_SS4END[4]),
    .I3(Tile_X0Y1_W2END[3]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q ),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3356_ (.I(_1646_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3357_ (.A1(_0178_),
    .A2(_1646_),
    .B(_0179_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3358_ (.I0(Tile_X0Y1_N2MID[2]),
    .I1(Tile_X0Y1_W2MID[2]),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .Z(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3359_ (.A1(_0178_),
    .A2(_1649_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3360_ (.I0(Tile_X0Y1_N2MID[3]),
    .I1(Tile_X0Y1_E2MID[3]),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .I3(Tile_X0Y1_W2MID[3]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q ),
    .Z(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3361_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .A2(_1651_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q ),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3362_ (.A1(_1645_),
    .A2(_1648_),
    .B1(_1650_),
    .B2(_1652_),
    .ZN(\Tile_X0Y1_DSP_bot.C5 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3363_ (.A1(_0162_),
    .A2(\Tile_X0Y1_DSP_bot.C5 ),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3364_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[5] ),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3365_ (.A1(_0163_),
    .A2(_1653_),
    .A3(_1654_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3366_ (.A1(_0163_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[5] ),
    .B(_1655_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3367_ (.A1(_1362_),
    .A2(_1364_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3368_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .A2(_0421_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3369_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .B(_1658_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3370_ (.A1(Tile_X0Y1_N2MID[6]),
    .A2(_0180_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3371_ (.A1(Tile_X0Y1_E2MID[6]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3372_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .A2(_1659_),
    .B1(_1660_),
    .B2(_1661_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3373_ (.A1(_0048_),
    .A2(_0181_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q ),
    .ZN(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3374_ (.A1(_0181_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .B(_1663_),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3375_ (.A1(Tile_X0Y1_N2MID[7]),
    .A2(_0181_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3376_ (.A1(Tile_X0Y1_E2MID[7]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q ),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3377_ (.A1(_1665_),
    .A2(_1666_),
    .B(_0182_),
    .C(_1664_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3378_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .A2(_0672_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3379_ (.A1(Tile_X0Y0_S4END[7]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .B(_1668_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3380_ (.A1(_0042_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3381_ (.A1(Tile_X0Y1_EE4END[0]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .C(_1670_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3382_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(_1669_),
    .B(_1671_),
    .C(_0182_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3383_ (.I0(Tile_X0Y1_N2END[7]),
    .I1(Tile_X0Y1_E2END[7]),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q ),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3384_ (.A1(Tile_X0Y1_WW4END[0]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q ),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3385_ (.A1(_0063_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q ),
    .C(_1674_),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3386_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q ),
    .A2(_1673_),
    .B(_1675_),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3387_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ),
    .A2(_1676_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q ),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3388_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q ),
    .A2(_1662_),
    .A3(_1667_),
    .B1(_1672_),
    .B2(_1677_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3389_ (.I(_1678_),
    .ZN(\Tile_X0Y1_DSP_bot.C4 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3390_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[4] ),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3391_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(_1678_),
    .B(_1679_),
    .C(_0163_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3392_ (.A1(_0163_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[4] ),
    .B(_1680_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3393_ (.A1(_1346_),
    .A2(_1348_),
    .A3(_1357_),
    .Z(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3394_ (.A1(_1681_),
    .A2(_1682_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3395_ (.A1(_1340_),
    .A2(_1345_),
    .A3(_1356_),
    .Z(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3396_ (.I0(Tile_X0Y1_EE4END[3]),
    .I1(Tile_X0Y1_WW4END[1]),
    .I2(Tile_X0Y0_S4END[4]),
    .I3(_0242_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q ),
    .Z(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3397_ (.I0(Tile_X0Y1_NN4END[2]),
    .I1(Tile_X0Y1_E2END[1]),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q ),
    .Z(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3398_ (.A1(Tile_X0Y1_W2END[1]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q ),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3399_ (.A1(_0025_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q ),
    .C(_1687_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3400_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q ),
    .A2(_1686_),
    .B(_1688_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3401_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .A2(_1689_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3402_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .A2(_1685_),
    .B(_1690_),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3403_ (.I0(Tile_X0Y1_E2MID[0]),
    .I1(Tile_X0Y1_W2MID[0]),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q ),
    .Z(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3404_ (.A1(_0184_),
    .A2(_1692_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3405_ (.I0(Tile_X0Y1_N2MID[1]),
    .I1(Tile_X0Y1_E2MID[1]),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .I3(Tile_X0Y1_W2MID[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q ),
    .Z(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3406_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .A2(_1694_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q ),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3407_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q ),
    .A2(_1691_),
    .B1(_1693_),
    .B2(_1695_),
    .ZN(\Tile_X0Y1_DSP_bot.C3 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3408_ (.A1(_0162_),
    .A2(\Tile_X0Y1_DSP_bot.C3 ),
    .ZN(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3409_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[3] ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3410_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .A2(_0183_),
    .B1(_1696_),
    .B2(_1697_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3411_ (.A1(_1684_),
    .A2(_1698_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3412_ (.A1(_1354_),
    .A2(_1355_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3413_ (.I0(Tile_X0Y1_N2END[5]),
    .I1(Tile_X0Y1_E2END[5]),
    .I2(Tile_X0Y0_SS4END[5]),
    .I3(Tile_X0Y1_W2END[5]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q ),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3414_ (.A1(_0186_),
    .A2(_1701_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3415_ (.A1(_0186_),
    .A2(_0287_),
    .B(_1702_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q ),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3416_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3417_ (.A1(_0027_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .B(_0185_),
    .C(_1704_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3418_ (.I0(Tile_X0Y1_W2MID[4]),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3419_ (.A1(_0185_),
    .A2(_1706_),
    .B(_1705_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3420_ (.I(_1707_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3421_ (.A1(Tile_X0Y1_W2MID[5]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q ),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3422_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q ),
    .A2(_0454_),
    .B(_1709_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q ),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3423_ (.I0(Tile_X0Y1_N2MID[5]),
    .I1(Tile_X0Y1_E2MID[5]),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q ),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3424_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q ),
    .A2(_1711_),
    .B(_1710_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3425_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ),
    .A2(_1707_),
    .B(_1712_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3426_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q ),
    .A2(_1713_),
    .B(_1703_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3427_ (.I(_1714_),
    .ZN(\Tile_X0Y1_DSP_bot.C2 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3428_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[2] ),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3429_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(_1714_),
    .B(_1715_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3430_ (.I0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[2] ),
    .I1(_1716_),
    .S(_0163_),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3431_ (.A1(_1700_),
    .A2(_1717_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3432_ (.A1(_1338_),
    .A2(_1353_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3433_ (.A1(_0163_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[1] ),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3434_ (.I0(Tile_X0Y1_NN4END[2]),
    .I1(Tile_X0Y0_S4END[6]),
    .I2(Tile_X0Y1_E2END[2]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q ),
    .Z(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3435_ (.A1(Tile_X0Y1_N2END[3]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q ),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3436_ (.A1(_0043_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q ),
    .C(_1722_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3437_ (.I0(Tile_X0Y0_S2MID[3]),
    .I1(Tile_X0Y1_WW4END[1]),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q ),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3438_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q ),
    .A2(_1724_),
    .B(_1723_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3439_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_1725_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3440_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_1721_),
    .B(_1726_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3441_ (.I0(Tile_X0Y1_N2MID[2]),
    .I1(Tile_X0Y1_E2MID[2]),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3442_ (.A1(_0187_),
    .A2(_1728_),
    .ZN(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3443_ (.I0(Tile_X0Y1_N2MID[3]),
    .I1(Tile_X0Y1_E2MID[3]),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .I3(Tile_X0Y1_W2MID[3]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q ),
    .Z(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3444_ (.I(_1730_),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3445_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_1730_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3446_ (.A1(_1729_),
    .A2(_1732_),
    .B(_1727_),
    .ZN(\Tile_X0Y1_DSP_bot.C1 ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3447_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[1] ),
    .Z(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3448_ (.A1(_0162_),
    .A2(\Tile_X0Y1_DSP_bot.C1 ),
    .B(_1733_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3449_ (.A1(_1720_),
    .A2(_1734_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3450_ (.A1(_0163_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[0] ),
    .Z(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3451_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3452_ (.A1(_0044_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q ),
    .C(_1737_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3453_ (.I0(Tile_X0Y1_N4END[3]),
    .I1(Tile_X0Y1_E2END[3]),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q ),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3454_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q ),
    .A2(_1739_),
    .B(_1738_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3455_ (.I0(Tile_X0Y1_N2END[7]),
    .I1(Tile_X0Y1_EE4END[2]),
    .I2(Tile_X0Y0_S2MID[7]),
    .I3(Tile_X0Y1_W2END[7]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q ),
    .Z(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3456_ (.I(_1741_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3457_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .A2(_1742_),
    .B(_1740_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q ),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3458_ (.I0(Tile_X0Y1_N2MID[6]),
    .I1(Tile_X0Y1_W2MID[6]),
    .I2(Tile_X0Y1_E2MID[6]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3459_ (.I0(_1744_),
    .I1(_0272_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3460_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q ),
    .A2(_1745_),
    .B(_1743_),
    .ZN(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3461_ (.I(_1746_),
    .ZN(\Tile_X0Y1_DSP_bot.C0 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3462_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[0] ),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3463_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(_1746_),
    .B(_1747_),
    .C(_0163_),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3464_ (.A1(_1736_),
    .A2(_1748_),
    .ZN(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3465_ (.A1(_1121_),
    .A2(_1242_),
    .A3(_1736_),
    .A4(_1748_),
    .ZN(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3466_ (.A1(_1338_),
    .A2(_1353_),
    .A3(_1735_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3467_ (.A1(_1719_),
    .A2(_1720_),
    .A3(_1734_),
    .B1(_1750_),
    .B2(_1751_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3468_ (.A1(_1354_),
    .A2(_1355_),
    .A3(_1717_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3469_ (.A1(_1752_),
    .A2(_1753_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3470_ (.A1(_1718_),
    .A2(_1754_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3471_ (.A1(_1684_),
    .A2(_1698_),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3472_ (.A1(_1755_),
    .A2(_1756_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3473_ (.A1(_1699_),
    .A2(_1757_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3474_ (.A1(_1681_),
    .A2(_1682_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3475_ (.A1(_1758_),
    .A2(_1759_),
    .B(_1683_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3476_ (.A1(_1362_),
    .A2(_1364_),
    .A3(_1656_),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3477_ (.A1(_1365_),
    .A2(_1656_),
    .A3(_1657_),
    .B1(_1760_),
    .B2(_1761_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3478_ (.A1(_1366_),
    .A2(_1368_),
    .A3(_1639_),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3479_ (.A1(_1762_),
    .A2(_1763_),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3480_ (.A1(_1369_),
    .A2(_1370_),
    .A3(_1620_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3481_ (.A1(_1641_),
    .A2(_1764_),
    .B(_1765_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3482_ (.A1(_1371_),
    .A2(_1372_),
    .A3(_1595_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3483_ (.A1(_1622_),
    .A2(_1766_),
    .B(_1767_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3484_ (.A1(_1597_),
    .A2(_1768_),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3485_ (.A1(_1549_),
    .A2(_1550_),
    .B(_1597_),
    .C(_1768_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3486_ (.A1(_1551_),
    .A2(_1770_),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3487_ (.A1(_1482_),
    .A2(_1551_),
    .A3(_1770_),
    .B(_1481_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3488_ (.A1(_1451_),
    .A2(_1452_),
    .Z(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3489_ (.A1(_1772_),
    .A2(_1773_),
    .B(_1453_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3490_ (.A1(_1425_),
    .A2(_1426_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3491_ (.A1(_1774_),
    .A2(_1775_),
    .Z(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3492_ (.A1(_1427_),
    .A2(_1776_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3493_ (.A1(_1416_),
    .A2(_1417_),
    .B1(_1774_),
    .B2(_1775_),
    .C(_1427_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3494_ (.A1(_1400_),
    .A2(_1418_),
    .A3(_1778_),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3495_ (.A1(_1418_),
    .A2(_1778_),
    .B(_1400_),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3496_ (.A1(_1779_),
    .A2(_1780_),
    .Z(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3497_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[14] ),
    .ZN(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3498_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1781_),
    .B(_1782_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3499_ (.A1(_1752_),
    .A2(_1753_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3500_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[2] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3501_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1783_),
    .B(_1784_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3502_ (.A1(_1352_),
    .A2(_1749_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3503_ (.A1(_1750_),
    .A2(_1785_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3504_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[0] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3505_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1786_),
    .B(_1787_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3506_ (.A1(_1758_),
    .A2(_1759_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3507_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[4] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3508_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1788_),
    .B(_1789_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3509_ (.A1(_1755_),
    .A2(_1756_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3510_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[3] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3511_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1790_),
    .B(_1791_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3512_ (.A1(_1760_),
    .A2(_1761_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3513_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[5] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3514_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1792_),
    .B(_1793_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3515_ (.A1(_1762_),
    .A2(_1763_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3516_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[6] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3517_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1794_),
    .B(_1795_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3518_ (.A1(_1641_),
    .A2(_1764_),
    .A3(_1765_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3519_ (.A1(_1766_),
    .A2(_1796_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3520_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[7] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3521_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1797_),
    .B(_1798_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3522_ (.A1(_1549_),
    .A2(_1550_),
    .A3(_1769_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3523_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[9] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3524_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1799_),
    .B(_1800_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3525_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ),
    .I2(_1651_),
    .I3(_1604_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3526_ (.A1(_1482_),
    .A2(_1771_),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3527_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[10] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3528_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1801_),
    .B(_1802_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3529_ (.A1(_1772_),
    .A2(_1773_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3530_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[11] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3531_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1803_),
    .B(_1804_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3532_ (.A1(_1774_),
    .A2(_1775_),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3533_ (.A1(_1776_),
    .A2(_1805_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3534_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[12] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3535_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1806_),
    .B(_1807_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3536_ (.A1(_1399_),
    .A2(_1779_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3537_ (.A1(_1072_),
    .A2(_1393_),
    .B(_1391_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3538_ (.A1(_1395_),
    .A2(_1809_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3539_ (.A1(_1389_),
    .A2(_1395_),
    .A3(_1396_),
    .B(_1810_),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3540_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3541_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .Z(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3542_ (.I0(_0456_),
    .I1(Tile_X0Y0_E1END[3]),
    .I2(Tile_X0Y1_N2MID[7]),
    .I3(Tile_X0Y0_E2END[7]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .Z(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3543_ (.I0(Tile_X0Y0_S1END[1]),
    .I1(Tile_X0Y0_S2END[7]),
    .I2(Tile_X0Y0_S1END[3]),
    .I3(Tile_X0Y0_W1END[3]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3544_ (.I0(_1814_),
    .I1(_1815_),
    .I2(_1812_),
    .I3(_1813_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3545_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .I1(Tile_X0Y0_W2MID[2]),
    .I2(Tile_X0Y0_S2MID[2]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q ),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3546_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(_0346_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3547_ (.A1(_0126_),
    .A2(_1816_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q ),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3548_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3549_ (.A1(_0035_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q ),
    .C(_1819_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3550_ (.I0(Tile_X0Y1_N4END[6]),
    .I1(Tile_X0Y0_SS4END[2]),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3551_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_1821_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3552_ (.I(_1822_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3553_ (.I0(Tile_X0Y1_N2MID[3]),
    .I1(Tile_X0Y0_E2END[3]),
    .I2(Tile_X0Y0_SS4END[0]),
    .I3(Tile_X0Y0_W2END[3]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q ),
    .Z(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3554_ (.I(_1824_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3555_ (.A1(_1820_),
    .A2(_1823_),
    .B1(_1824_),
    .B2(_0126_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3556_ (.A1(_1817_),
    .A2(_1818_),
    .B1(_1826_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q ),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3557_ (.A1(_0162_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3558_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[15] ),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3559_ (.A1(_0163_),
    .A2(_1827_),
    .A3(_1828_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3560_ (.A1(_0163_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[15] ),
    .B(_1829_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3561_ (.I(_1830_),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3562_ (.A1(_1811_),
    .A2(_1831_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3563_ (.A1(_1811_),
    .A2(_1831_),
    .Z(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3564_ (.A1(_1808_),
    .A2(_1811_),
    .A3(_1831_),
    .Z(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3565_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[15] ),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3566_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1834_),
    .B(_1835_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3567_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ),
    .A2(_1811_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3568_ (.A1(_0163_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[16] ),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3569_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3570_ (.A1(_0080_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q ),
    .C(_1838_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3571_ (.A1(Tile_X0Y0_S4END[1]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q ),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3572_ (.A1(_0058_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ),
    .B(_1840_),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3573_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ),
    .A2(_1839_),
    .A3(_1841_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3574_ (.I0(Tile_X0Y1_NN4END[5]),
    .I1(Tile_X0Y0_S2END[5]),
    .I2(Tile_X0Y0_E2END[5]),
    .I3(Tile_X0Y0_W2END[5]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q ),
    .Z(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3575_ (.I(_1843_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3576_ (.A1(_0128_),
    .A2(_1843_),
    .B(_0129_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3577_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .I1(Tile_X0Y0_S2MID[5]),
    .I2(Tile_X0Y0_E2MID[5]),
    .I3(Tile_X0Y0_W2MID[5]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ),
    .Z(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3578_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ),
    .A2(_1846_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3579_ (.I0(Tile_X0Y0_E2MID[4]),
    .I1(Tile_X0Y0_W2MID[4]),
    .I2(Tile_X0Y0_S2MID[4]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q ),
    .Z(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3580_ (.I(_1848_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3581_ (.A1(_0128_),
    .A2(_1848_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q ),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3582_ (.A1(_1842_),
    .A2(_1845_),
    .B1(_1847_),
    .B2(_1850_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3583_ (.I0(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[16] ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ),
    .S(_0162_),
    .Z(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3584_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .A2(_1851_),
    .B(_1837_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3585_ (.A1(_1836_),
    .A2(_1852_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3586_ (.A1(_1836_),
    .A2(_1852_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3587_ (.A1(_1399_),
    .A2(_1779_),
    .A3(_1833_),
    .B(_1832_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3588_ (.A1(_1854_),
    .A2(_1855_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3589_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[16] ),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3590_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1856_),
    .B(_1857_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3591_ (.A1(_1854_),
    .A2(_1855_),
    .B(_1853_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3592_ (.A1(_0163_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[17] ),
    .Z(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3593_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .Z(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3594_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .Z(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3595_ (.I0(_0456_),
    .I1(Tile_X0Y0_E1END[3]),
    .I2(Tile_X0Y1_N2MID[7]),
    .I3(Tile_X0Y0_E2END[7]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .Z(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3596_ (.I0(Tile_X0Y0_S1END[1]),
    .I1(Tile_X0Y0_S2END[7]),
    .I2(Tile_X0Y0_S1END[3]),
    .I3(Tile_X0Y0_W1END[3]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .Z(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3597_ (.I0(_1862_),
    .I1(_1863_),
    .I2(_1860_),
    .I3(_1861_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3598_ (.A1(Tile_X0Y0_W2MID[0]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q ),
    .Z(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3599_ (.A1(_0130_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ),
    .B(_1864_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3600_ (.A1(_0130_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3601_ (.A1(Tile_X0Y0_E2MID[0]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q ),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3602_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q ),
    .A2(_1865_),
    .B1(_1866_),
    .B2(_1867_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3603_ (.A1(Tile_X0Y0_E2MID[1]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q ),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3604_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ),
    .A2(_0428_),
    .A3(_0435_),
    .B(_1869_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3605_ (.A1(Tile_X0Y0_W2MID[1]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3606_ (.A1(_0025_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q ),
    .C(_1871_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3607_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(_1870_),
    .A3(_1872_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3608_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q ),
    .A2(_1868_),
    .A3(_1873_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3609_ (.A1(Tile_X0Y0_EE4END[3]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q ),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3610_ (.A1(_0033_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q ),
    .B(_1875_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3611_ (.A1(Tile_X0Y0_W2END[1]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q ),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3612_ (.A1(_0066_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q ),
    .C(_1877_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3613_ (.A1(_1876_),
    .A2(_1878_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3614_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(_1879_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q ),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3615_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(_0321_),
    .B(_1880_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3616_ (.A1(_1874_),
    .A2(_1881_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3617_ (.I0(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[17] ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ),
    .S(_0162_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3618_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .A2(_1882_),
    .B(_1859_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3619_ (.A1(_1836_),
    .A2(_1883_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3620_ (.A1(_1836_),
    .A2(_1858_),
    .A3(_1883_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3621_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[17] ),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3622_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1885_),
    .B(_1886_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3623_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3624_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(_0454_),
    .B(_1887_),
    .C(_0191_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3625_ (.A1(_0192_),
    .A2(_0255_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3626_ (.A1(Tile_X0Y1_N2MID[0]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .ZN(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3627_ (.A1(Tile_X0Y0_E1END[0]),
    .A2(_0192_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3628_ (.A1(Tile_X0Y0_E2END[0]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .B(_0193_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3629_ (.A1(_1889_),
    .A2(_1890_),
    .B1(_1891_),
    .B2(_1892_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3630_ (.I0(Tile_X0Y0_S1END[0]),
    .I1(Tile_X0Y0_S2END[0]),
    .I2(Tile_X0Y0_S1END[2]),
    .I3(Tile_X0Y0_W1END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .Z(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3631_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ),
    .A2(_1894_),
    .B(_1893_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3632_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3633_ (.I(_1896_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3634_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3635_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ),
    .A2(_1898_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3636_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ),
    .A2(_1897_),
    .B(_1899_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3637_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(_1900_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3638_ (.A1(_0190_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3639_ (.A1(_1895_),
    .A2(_1901_),
    .B(_1902_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3640_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ),
    .A2(_1888_),
    .A3(_1903_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3641_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3642_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .Z(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3643_ (.I0(_0255_),
    .I1(Tile_X0Y1_N2MID[0]),
    .I2(Tile_X0Y0_E1END[0]),
    .I3(Tile_X0Y0_EE4END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .Z(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3644_ (.I0(Tile_X0Y0_S1END[0]),
    .I1(Tile_X0Y0_S2END[0]),
    .I2(Tile_X0Y0_W1END[0]),
    .I3(Tile_X0Y0_W1END[2]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3645_ (.I0(_1907_),
    .I1(_1908_),
    .I2(_1905_),
    .I3(_1906_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3646_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ),
    .Z(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3647_ (.A1(_0190_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ),
    .B(_1909_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3648_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .Z(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3649_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .Z(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3650_ (.I0(_0255_),
    .I1(Tile_X0Y1_N2MID[0]),
    .I2(Tile_X0Y0_E1END[0]),
    .I3(Tile_X0Y0_E2END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3651_ (.I0(Tile_X0Y0_S1END[0]),
    .I1(Tile_X0Y0_S1END[2]),
    .I2(Tile_X0Y0_SS4END[0]),
    .I3(Tile_X0Y0_WW4END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3652_ (.I0(_1913_),
    .I1(_1914_),
    .I2(_1911_),
    .I3(_1912_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3653_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3654_ (.A1(_0190_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ),
    .B(_1915_),
    .C(_0191_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3655_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ),
    .A2(_1910_),
    .A3(_1916_),
    .B(_1904_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3656_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[19] ),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3657_ (.A1(_0162_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3658_ (.A1(_1917_),
    .A2(_1918_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3659_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ),
    .B(_1919_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3660_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .A2(_0315_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3661_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ),
    .B(_1921_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3662_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .ZN(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3663_ (.A1(_0189_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3664_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ),
    .A2(_1922_),
    .B1(_1923_),
    .B2(_1924_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3665_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ),
    .S0(_0189_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ),
    .Z(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3666_ (.I0(_1926_),
    .I1(_1925_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3667_ (.A1(_0162_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3668_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[18] ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3669_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .A2(_0188_),
    .B1(_1927_),
    .B2(_1928_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3670_ (.I(_1929_),
    .ZN(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3671_ (.A1(_1854_),
    .A2(_1855_),
    .B1(_1883_),
    .B2(_1836_),
    .C(_1853_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3672_ (.A1(_1884_),
    .A2(_1931_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3673_ (.A1(_1884_),
    .A2(_1929_),
    .A3(_1931_),
    .Z(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3674_ (.A1(_1836_),
    .A2(_1931_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3675_ (.A1(_1836_),
    .A2(_1930_),
    .B1(_1933_),
    .B2(_1934_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3676_ (.A1(_1920_),
    .A2(_1935_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3677_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3678_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1936_),
    .B(_1937_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3679_ (.A1(_1416_),
    .A2(_1417_),
    .A3(_1777_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3680_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[13] ),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3681_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1938_),
    .B(_1939_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3682_ (.A1(_1836_),
    .A2(_1930_),
    .A3(_1932_),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3683_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[18] ),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3684_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1940_),
    .B(_1941_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3685_ (.A1(_1750_),
    .A2(_1751_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3686_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[1] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3687_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1942_),
    .B(_1943_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3688_ (.A1(_1622_),
    .A2(_1766_),
    .A3(_1767_),
    .Z(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3689_ (.A1(_1768_),
    .A2(_1944_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3690_ (.I(_1945_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3691_ (.A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[8] ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3692_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .A2(_1946_),
    .B(_1947_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3693_ (.I0(_0456_),
    .I1(Tile_X0Y0_E2END[1]),
    .I2(Tile_X0Y1_N2MID[1]),
    .I3(Tile_X0Y0_E6END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .Z(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3694_ (.I0(Tile_X0Y0_S2END[1]),
    .I1(Tile_X0Y0_S4END[1]),
    .I2(Tile_X0Y0_W2END[1]),
    .I3(Tile_X0Y0_W6END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .Z(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3695_ (.A1(_0067_),
    .A2(_1949_),
    .Z(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3696_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ),
    .A2(_1948_),
    .B(_1950_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3697_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .Z(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3698_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ),
    .A2(_1952_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3699_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .Z(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3700_ (.A1(_0067_),
    .A2(_1954_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3701_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ),
    .A2(_1951_),
    .B1(_1953_),
    .B2(_1955_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3702_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I1(_0630_),
    .I2(_1956_),
    .I3(_0653_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3703_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I1(_0346_),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ),
    .I3(_0321_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3704_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I1(_0374_),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ),
    .I3(_0407_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3705_ (.I0(Tile_X0Y1_N2MID[2]),
    .I1(Tile_X0Y1_N4END[5]),
    .I2(Tile_X0Y0_E6END[1]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3706_ (.I0(Tile_X0Y1_N2MID[3]),
    .I1(Tile_X0Y1_N4END[6]),
    .I2(Tile_X0Y0_E6END[0]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3707_ (.I0(Tile_X0Y1_N2MID[0]),
    .I1(Tile_X0Y1_N4END[7]),
    .I2(Tile_X0Y0_W6END[1]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3708_ (.I0(Tile_X0Y1_N2MID[1]),
    .I1(Tile_X0Y0_W6END[0]),
    .I2(Tile_X0Y1_N4END[4]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3709_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I1(_0482_),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .I3(_0468_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3710_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .Z(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3711_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .A2(_0210_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3712_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .B(_1958_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3713_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .A2(_0214_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3714_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .B(_1960_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3715_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ),
    .A2(_1959_),
    .A3(_1961_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3716_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ),
    .A2(_1957_),
    .B(_1962_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3717_ (.I0(Tile_X0Y0_E6END[1]),
    .I1(Tile_X0Y0_W2END[1]),
    .I2(Tile_X0Y0_SS4END[1]),
    .I3(Tile_X0Y0_W6END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .Z(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3718_ (.I(_1964_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3719_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ),
    .A2(_1965_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3720_ (.I0(Tile_X0Y1_N2MID[1]),
    .I1(Tile_X0Y1_N4END[5]),
    .I2(Tile_X0Y0_E1END[3]),
    .I3(Tile_X0Y0_E2END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .Z(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3721_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ),
    .A2(_1967_),
    .B(_1966_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3722_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ),
    .A2(_1968_),
    .B(_1963_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3723_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I1(_0630_),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ),
    .I3(_0653_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3724_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I1(_0346_),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ),
    .I3(_0321_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3725_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ),
    .A2(_0408_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3726_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ),
    .B(_1969_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q ),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3727_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ),
    .A2(_0210_),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3728_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ),
    .A2(_0374_),
    .B(_1971_),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3729_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q ),
    .A2(_1972_),
    .B(_1970_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3730_ (.I0(Tile_X0Y0_E6END[1]),
    .I1(Tile_X0Y0_S4END[1]),
    .I2(Tile_X0Y0_S2END[2]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3731_ (.I0(Tile_X0Y0_E6END[0]),
    .I1(Tile_X0Y0_S4END[2]),
    .I2(Tile_X0Y0_S2END[3]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3732_ (.I0(Tile_X0Y0_S2END[0]),
    .I1(Tile_X0Y0_W6END[1]),
    .I2(Tile_X0Y0_S4END[3]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3733_ (.I0(Tile_X0Y0_S2END[1]),
    .I1(Tile_X0Y0_S4END[0]),
    .I2(Tile_X0Y0_W6END[0]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3734_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I1(_0482_),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .I3(_0468_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3735_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I1(_0630_),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .I3(_0653_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3736_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .I2(_0346_),
    .I3(_0321_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3737_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(_0374_),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .I3(_0407_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3738_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_0916_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3739_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .B(_1973_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3740_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_1825_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3741_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_0875_),
    .B(_1975_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3742_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ),
    .A2(_1974_),
    .B(_1976_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3743_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .I1(Tile_X0Y0_E1END[2]),
    .I2(Tile_X0Y0_W1END[2]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ),
    .Z(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3744_ (.I0(_1978_),
    .I1(_1977_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3745_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3746_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .A2(_0673_),
    .B(_1979_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3747_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .A2(_1442_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3748_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .A2(_0815_),
    .B(_1981_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3749_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q ),
    .A2(_1982_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3750_ (.I0(_0456_),
    .I1(Tile_X0Y0_W1END[3]),
    .I2(Tile_X0Y0_E1END[3]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .Z(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3751_ (.A1(_1980_),
    .A2(_1983_),
    .B1(_1984_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q ),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3752_ (.I(_1985_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3753_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(_0880_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3754_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(_0346_),
    .B(_1986_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ),
    .ZN(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3755_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(_1430_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3756_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .B(_1988_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3757_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ),
    .A2(_1989_),
    .B(_1987_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3758_ (.I0(_0255_),
    .I1(Tile_X0Y0_W1END[0]),
    .I2(Tile_X0Y0_E1END[0]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .Z(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3759_ (.I0(_1991_),
    .I1(_1990_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3760_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3761_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ),
    .A2(_1420_),
    .B(_1992_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3762_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ),
    .A2(_0922_),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3763_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ),
    .A2(_1848_),
    .B(_1994_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3764_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q ),
    .A2(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3765_ (.I0(_0306_),
    .I1(Tile_X0Y0_W1END[1]),
    .I2(Tile_X0Y0_E1END[1]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ),
    .Z(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3766_ (.A1(_1993_),
    .A2(_1996_),
    .B1(_1997_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q ),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3767_ (.I(_1998_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3768_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ),
    .A2(_0916_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3769_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .B(_1999_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3770_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ),
    .A2(_0525_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3771_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ),
    .A2(_0875_),
    .B(_2001_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3772_ (.A1(_2000_),
    .A2(_2002_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3773_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .I1(Tile_X0Y0_S1END[2]),
    .I2(Tile_X0Y0_E1END[2]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ),
    .Z(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3774_ (.I0(_2004_),
    .I1(_2003_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3775_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3776_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .A2(_0673_),
    .B(_2005_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3777_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .A2(_1460_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3778_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .A2(_0815_),
    .B(_2007_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3779_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q ),
    .A2(_2008_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3780_ (.I0(_0456_),
    .I1(Tile_X0Y0_E1END[3]),
    .I2(Tile_X0Y0_S1END[3]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ),
    .Z(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3781_ (.A1(_2006_),
    .A2(_2009_),
    .B1(_2010_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q ),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3782_ (.I(_2011_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3783_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .I1(_0346_),
    .I2(_1429_),
    .I3(_0538_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3784_ (.I0(_0255_),
    .I1(Tile_X0Y0_S1END[0]),
    .I2(Tile_X0Y0_E1END[0]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ),
    .Z(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3785_ (.I0(_2013_),
    .I1(_2012_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3786_ (.I0(_0306_),
    .I1(Tile_X0Y0_S1END[1]),
    .I2(Tile_X0Y0_E1END[1]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ),
    .Z(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3787_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .I1(_1421_),
    .I2(_1848_),
    .I3(_0884_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ),
    .Z(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3788_ (.I0(_2014_),
    .I1(_2015_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3789_ (.I0(Tile_X0Y0_E1END[3]),
    .I1(Tile_X0Y0_W1END[3]),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .Z(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3790_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_2016_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3791_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .Z(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3792_ (.A1(_0194_),
    .A2(_2018_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3793_ (.I0(_0915_),
    .I1(_1429_),
    .I2(_0875_),
    .I3(_0346_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3794_ (.A1(_0194_),
    .A2(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3795_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .Z(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3796_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_2022_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3797_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ),
    .A2(_2017_),
    .A3(_2019_),
    .B1(_2021_),
    .B2(_2023_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3798_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .A2(_0674_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3799_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .A2(_0816_),
    .B(_2024_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3800_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .A2(_1849_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3801_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .A2(_1421_),
    .B(_2026_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3802_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_2027_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3803_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .Z(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3804_ (.A1(_2025_),
    .A2(_2028_),
    .B1(_2029_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q ),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3805_ (.I0(Tile_X0Y0_E1END[2]),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I2(Tile_X0Y0_W1END[2]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .Z(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3806_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .Z(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3807_ (.I(_2032_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3808_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_2033_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q ),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3809_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_2031_),
    .B(_2034_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3810_ (.A1(_2030_),
    .A2(_2035_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3811_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ),
    .A2(_0916_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3812_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .B(_2036_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3813_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ),
    .A2(_1879_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3814_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ),
    .A2(_0875_),
    .B(_2038_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3815_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ),
    .A2(_2037_),
    .B(_2039_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3816_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .I1(Tile_X0Y0_E1END[2]),
    .I2(Tile_X0Y0_W1END[2]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3817_ (.I0(_2041_),
    .I1(_2040_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3818_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I1(_0674_),
    .I2(_0815_),
    .I3(_1410_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ),
    .Z(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3819_ (.I0(_0456_),
    .I1(Tile_X0Y0_W1END[3]),
    .I2(Tile_X0Y0_E1END[3]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ),
    .Z(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3820_ (.I0(_2043_),
    .I1(_2042_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3821_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .A2(_1430_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3822_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .B(_2044_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3823_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .A2(_0771_),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3824_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .A2(_0346_),
    .B(_2046_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3825_ (.A1(_2045_),
    .A2(_2047_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3826_ (.I0(_0255_),
    .I1(Tile_X0Y0_W1END[0]),
    .I2(Tile_X0Y0_E1END[0]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .Z(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3827_ (.I0(_2049_),
    .I1(_2048_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3828_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3829_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ),
    .A2(_1420_),
    .B(_2050_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3830_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ),
    .A2(_0594_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3831_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ),
    .A2(_1848_),
    .B(_2052_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ),
    .ZN(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3832_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q ),
    .A2(_2053_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3833_ (.I0(_0306_),
    .I1(Tile_X0Y0_W1END[1]),
    .I2(Tile_X0Y0_E1END[1]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ),
    .Z(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3834_ (.A1(_2051_),
    .A2(_2054_),
    .B1(_2055_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q ),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3835_ (.I(_2056_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3836_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ),
    .A2(_0916_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3837_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .B(_2057_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3838_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ),
    .A2(_1844_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3839_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ),
    .A2(_0875_),
    .B(_2059_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3840_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ),
    .A2(_2058_),
    .B(_2060_),
    .ZN(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3841_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .I1(Tile_X0Y0_S1END[2]),
    .I2(Tile_X0Y0_W1END[2]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3842_ (.I0(_2062_),
    .I1(_2061_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3843_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I1(_0674_),
    .I2(_0815_),
    .I3(_1419_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ),
    .Z(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3844_ (.I0(_0456_),
    .I1(Tile_X0Y0_W1END[3]),
    .I2(Tile_X0Y0_S1END[3]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3845_ (.I0(_2064_),
    .I1(_2063_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3846_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(_1430_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3847_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .B(_2065_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3848_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(_0795_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3849_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(_0346_),
    .B(_2067_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3850_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ),
    .A2(_2066_),
    .B(_2068_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3851_ (.I0(_0255_),
    .I1(Tile_X0Y0_W1END[0]),
    .I2(Tile_X0Y0_S1END[0]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .Z(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3852_ (.I0(_2070_),
    .I1(_2069_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3853_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3854_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ),
    .A2(_1420_),
    .B(_2071_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3855_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ),
    .A2(_0607_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3856_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ),
    .A2(_1848_),
    .B(_2073_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3857_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q ),
    .A2(_2074_),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3858_ (.I0(_0306_),
    .I1(Tile_X0Y0_W1END[1]),
    .I2(Tile_X0Y0_S1END[1]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3859_ (.A1(_2072_),
    .A2(_2075_),
    .B1(_2076_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q ),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3860_ (.I(_2077_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3861_ (.I0(Tile_X0Y0_E1END[3]),
    .I1(Tile_X0Y0_W1END[3]),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .Z(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3862_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_2078_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3863_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .Z(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3864_ (.A1(_0195_),
    .A2(_2080_),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3865_ (.I0(_0915_),
    .I1(_1429_),
    .I2(_0875_),
    .I3(_0346_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3866_ (.A1(_0195_),
    .A2(_2082_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3867_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3868_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_2084_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3869_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ),
    .A2(_2079_),
    .A3(_2081_),
    .B1(_2083_),
    .B2(_2085_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3870_ (.I0(Tile_X0Y0_E1END[2]),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I2(Tile_X0Y0_W1END[2]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .Z(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3871_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3872_ (.I(_2087_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3873_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_2088_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q ),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3874_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_2086_),
    .B(_2089_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3875_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .A2(_0816_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3876_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .A2(_0674_),
    .B(_2091_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3877_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .A2(_1849_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3878_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .A2(_1421_),
    .B(_2093_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3879_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .A2(_2092_),
    .B(_2094_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3880_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3881_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_2096_),
    .B(_2095_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q ),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3882_ (.A1(_2090_),
    .A2(_2097_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3883_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I1(_0482_),
    .I2(_0561_),
    .I3(_0468_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3884_ (.I0(Tile_X0Y1_N2END[2]),
    .I1(Tile_X0Y1_E6END[1]),
    .I2(Tile_X0Y1_N4END[1]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q ),
    .Z(\Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3885_ (.I0(Tile_X0Y1_N2END[3]),
    .I1(Tile_X0Y1_E6END[0]),
    .I2(Tile_X0Y1_N4END[2]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q ),
    .Z(\Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3886_ (.I0(Tile_X0Y1_N2END[0]),
    .I1(Tile_X0Y1_N4END[3]),
    .I2(Tile_X0Y1_W6END[1]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q ),
    .Z(\Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3887_ (.I0(Tile_X0Y1_N2END[1]),
    .I1(Tile_X0Y1_N4END[0]),
    .I2(Tile_X0Y1_W6END[0]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q ),
    .Z(\Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3888_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I1(_0254_),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .I3(_0231_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3889_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I1(_0272_),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .I3(_0286_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3890_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .I2(_1651_),
    .I3(_1604_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3891_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I1(_0455_),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .I3(_0436_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3892_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I1(_0254_),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .I3(_0231_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3893_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .Z(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3894_ (.A1(_0197_),
    .A2(_2098_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3895_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3896_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .A2(_2100_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3897_ (.I0(Tile_X0Y1_E6END[1]),
    .I1(Tile_X0Y1_W2END[1]),
    .I2(Tile_X0Y0_S2MID[1]),
    .I3(Tile_X0Y1_W6END[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3898_ (.A1(_0197_),
    .A2(_2102_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3899_ (.I0(Tile_X0Y1_N1END[3]),
    .I1(Tile_X0Y1_N4END[1]),
    .I2(Tile_X0Y1_N2END[1]),
    .I3(Tile_X0Y1_EE4END[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .Z(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3900_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .A2(_2104_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3901_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_2103_),
    .A3(_2105_),
    .B1(_2099_),
    .B2(_2101_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3902_ (.A1(_0196_),
    .A2(_0286_),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3903_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q ),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3904_ (.A1(_0196_),
    .A2(_0272_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3905_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3906_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q ),
    .A2(_2108_),
    .A3(_2109_),
    .B1(_2106_),
    .B2(_2107_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3907_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ),
    .I2(_1651_),
    .I3(_1604_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3908_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ),
    .I2(_0455_),
    .I3(_0436_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3909_ (.I0(Tile_X0Y1_E6END[1]),
    .I1(Tile_X0Y0_S4END[5]),
    .I2(Tile_X0Y0_S2MID[2]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3910_ (.I0(Tile_X0Y1_E6END[0]),
    .I1(Tile_X0Y0_S2MID[3]),
    .I2(Tile_X0Y0_S4END[6]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3911_ (.I0(Tile_X0Y0_S2MID[0]),
    .I1(Tile_X0Y0_S4END[7]),
    .I2(Tile_X0Y1_W6END[1]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3912_ (.I0(Tile_X0Y0_S2MID[1]),
    .I1(Tile_X0Y0_S4END[4]),
    .I2(Tile_X0Y1_W6END[0]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3913_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(_0254_),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .I3(_0231_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3914_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .Z(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3915_ (.I(_2110_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3916_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(_2111_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3917_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .Z(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3918_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(_2113_),
    .B(_2112_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3919_ (.I0(Tile_X0Y0_S2MID[1]),
    .I1(Tile_X0Y0_S4END[5]),
    .I2(Tile_X0Y1_W2END[1]),
    .I3(Tile_X0Y1_W6END[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .Z(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3920_ (.I(_2115_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3921_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(_2116_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3922_ (.I0(Tile_X0Y1_NN4END[1]),
    .I1(Tile_X0Y1_E1END[3]),
    .I2(Tile_X0Y1_E2END[1]),
    .I3(Tile_X0Y1_E6END[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3923_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(_2118_),
    .B(_2117_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3924_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ),
    .A2(_2119_),
    .B(_2114_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3925_ (.A1(_0198_),
    .A2(_0286_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3926_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q ),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3927_ (.A1(_0198_),
    .A2(_0272_),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3928_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .ZN(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3929_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q ),
    .A2(_2122_),
    .A3(_2123_),
    .B1(_2120_),
    .B2(_2121_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3930_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ),
    .I2(_1651_),
    .I3(_1604_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3931_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(_0455_),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .I3(_0436_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3932_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ),
    .A2(_0956_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3933_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .B(_2124_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3934_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ),
    .A2(_1647_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3935_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ),
    .A2(_1188_),
    .B(_2126_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3936_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ),
    .A2(_2125_),
    .B(_2127_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3937_ (.I0(Tile_X0Y1_N1END[2]),
    .I1(Tile_X0Y1_E1END[2]),
    .I2(Tile_X0Y1_W1END[2]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3938_ (.I0(_2129_),
    .I1(_2128_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q ),
    .Z(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3939_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .A2(_1725_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3940_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .A2(_1026_),
    .B(_2130_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3941_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .A2(_0827_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3942_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .B(_2132_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3943_ (.A1(_2131_),
    .A2(_2133_),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3944_ (.I0(Tile_X0Y1_N1END[3]),
    .I1(Tile_X0Y1_E1END[3]),
    .I2(Tile_X0Y1_W1END[3]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ),
    .Z(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3945_ (.I0(_2135_),
    .I1(_2134_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q ),
    .Z(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3946_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .I1(_1651_),
    .I2(_1730_),
    .I3(_1164_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3947_ (.I0(Tile_X0Y1_N1END[0]),
    .I1(Tile_X0Y1_E1END[0]),
    .I2(Tile_X0Y1_W1END[0]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3948_ (.I0(_2137_),
    .I1(_2136_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q ),
    .Z(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3949_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .I1(_1629_),
    .I2(_1708_),
    .I3(_0978_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3950_ (.I0(Tile_X0Y1_N1END[1]),
    .I1(Tile_X0Y1_W1END[1]),
    .I2(Tile_X0Y1_E1END[1]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3951_ (.I0(_2139_),
    .I1(_2138_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q ),
    .Z(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3952_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .A2(_0956_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3953_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .B(_2140_),
    .ZN(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3954_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .A2(_1676_),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3955_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .A2(_1188_),
    .B(_2142_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3956_ (.A1(_2141_),
    .A2(_2143_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3957_ (.I0(Tile_X0Y1_N1END[2]),
    .I1(Tile_X0Y1_E1END[2]),
    .I2(_0351_),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3958_ (.I0(_2145_),
    .I1(_2144_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3959_ (.I0(Tile_X0Y1_N1END[3]),
    .I1(Tile_X0Y1_E1END[3]),
    .I2(_0412_),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ),
    .Z(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3960_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .A2(_1742_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3961_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .A2(_1026_),
    .B(_2147_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3962_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .A2(_0827_),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3963_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .B(_2149_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3964_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ),
    .A2(_2150_),
    .B(_2148_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q ),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3965_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q ),
    .A2(_2146_),
    .B(_2151_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3966_ (.I(_2152_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3967_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .A2(_0207_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3968_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .A2(_0489_),
    .B(_2153_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3969_ (.A1(Tile_X0Y1_N1END[0]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3970_ (.A1(_0021_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ),
    .C(_2155_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3971_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q ),
    .A2(_2156_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3972_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .I1(_1651_),
    .I2(_1730_),
    .I3(_1222_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .Z(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3973_ (.I(_2158_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3974_ (.A1(_2154_),
    .A2(_2157_),
    .B1(_2159_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q ),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3975_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .A2(_1094_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3976_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .A2(_1629_),
    .B(_2160_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3977_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .A2(_1707_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3978_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .B(_2162_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3979_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ),
    .A2(_2163_),
    .B(_2161_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q ),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3980_ (.I0(Tile_X0Y1_N1END[1]),
    .I1(Tile_X0Y1_E1END[1]),
    .I2(_0657_),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ),
    .Z(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3981_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q ),
    .A2(_2165_),
    .B(_2164_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3982_ (.I(_2166_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3983_ (.I0(Tile_X0Y1_E1END[3]),
    .I1(Tile_X0Y1_W1END[3]),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3984_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ),
    .A2(_2167_),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3985_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .Z(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3986_ (.A1(_0199_),
    .A2(_2169_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3987_ (.I0(_0955_),
    .I1(_1188_),
    .I2(_1730_),
    .I3(_1651_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .Z(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3988_ (.A1(_0199_),
    .A2(_2171_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3989_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .Z(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3990_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ),
    .A2(_2173_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q ),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3991_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q ),
    .A2(_2168_),
    .A3(_2170_),
    .B1(_2172_),
    .B2(_2174_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3992_ (.A1(_0200_),
    .A2(_1026_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3993_ (.A1(_0200_),
    .A2(_0827_),
    .B(_2175_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .ZN(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3994_ (.A1(_0200_),
    .A2(_1707_),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3995_ (.A1(_0200_),
    .A2(_1629_),
    .B(_2177_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3996_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_2178_),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3997_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .Z(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3998_ (.A1(_2176_),
    .A2(_2179_),
    .B1(_2180_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q ),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3999_ (.I0(Tile_X0Y1_E1END[2]),
    .I1(Tile_X0Y1_W1END[2]),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .Z(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4000_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .Z(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4001_ (.I(_2183_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4002_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_2184_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q ),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4003_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_2182_),
    .B(_2185_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4004_ (.A1(_2181_),
    .A2(_2186_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4005_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .A2(_0956_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4006_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .B(_2187_),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4007_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .A2(_1608_),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4008_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .A2(_1188_),
    .B(_2189_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4009_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ),
    .A2(_2188_),
    .B(_2190_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4010_ (.I0(Tile_X0Y1_N1END[2]),
    .I1(Tile_X0Y1_E1END[2]),
    .I2(Tile_X0Y1_W1END[2]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ),
    .Z(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4011_ (.I0(_2192_),
    .I1(_2191_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4012_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ),
    .A2(_1689_),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4013_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ),
    .A2(_1026_),
    .B(_2193_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4014_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ),
    .A2(_0827_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4015_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .B(_2195_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4016_ (.A1(_2194_),
    .A2(_2196_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4017_ (.I0(Tile_X0Y1_N1END[3]),
    .I1(Tile_X0Y1_E1END[3]),
    .I2(Tile_X0Y1_W1END[3]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ),
    .Z(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4018_ (.I0(_2198_),
    .I1(_2197_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4019_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ),
    .A2(_1731_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4020_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .B(_2199_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4021_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ),
    .A2(_0716_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4022_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ),
    .A2(_1651_),
    .B(_2201_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4023_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ),
    .A2(_2200_),
    .B(_2202_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4024_ (.I0(Tile_X0Y1_N1END[0]),
    .I1(Tile_X0Y1_E1END[0]),
    .I2(Tile_X0Y1_W1END[0]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ),
    .Z(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4025_ (.I0(_2204_),
    .I1(_2203_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4026_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ),
    .A2(_0743_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4027_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ),
    .A2(_1629_),
    .B(_2205_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4028_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ),
    .A2(_1707_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4029_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .B(_2207_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4030_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ),
    .A2(_2208_),
    .B(_2206_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4031_ (.I0(Tile_X0Y1_N1END[1]),
    .I1(Tile_X0Y1_W1END[1]),
    .I2(Tile_X0Y1_E1END[1]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4032_ (.I0(_2210_),
    .I1(_2209_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4033_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .A2(_1627_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4034_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .A2(_1188_),
    .B(_2211_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4035_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .A2(_0956_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4036_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .B(_2213_),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4037_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ),
    .A2(_2214_),
    .B(_2212_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4038_ (.I0(Tile_X0Y1_N1END[2]),
    .I1(Tile_X0Y1_W1END[2]),
    .I2(_0351_),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .Z(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4039_ (.I0(_2216_),
    .I1(_2215_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q ),
    .Z(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4040_ (.I0(_1026_),
    .I1(_1701_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ),
    .Z(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4041_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4042_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ),
    .A2(_0827_),
    .B(_2218_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4043_ (.I0(Tile_X0Y1_N1END[3]),
    .I1(Tile_X0Y1_W1END[3]),
    .I2(_0412_),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ),
    .Z(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4044_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ),
    .A2(_2217_),
    .B(_2219_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4045_ (.A1(_0201_),
    .A2(_2220_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4046_ (.A1(_0201_),
    .A2(_2221_),
    .B(_2222_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4047_ (.A1(Tile_X0Y1_N1END[0]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4048_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .A2(_0488_),
    .B(_2223_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4049_ (.I0(Tile_X0Y1_W1END[0]),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .Z(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4050_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ),
    .A2(_2225_),
    .B(_2224_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q ),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4051_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4052_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .A2(_1731_),
    .B(_2227_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4053_ (.I0(_1651_),
    .I1(_1045_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .Z(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4054_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ),
    .A2(_2229_),
    .B(_2228_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4055_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q ),
    .A2(_2230_),
    .B(_2226_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4056_ (.I0(Tile_X0Y1_N1END[1]),
    .I1(Tile_X0Y1_W1END[1]),
    .I2(_0657_),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .Z(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4057_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .A2(_0839_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4058_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .A2(_1629_),
    .B(_2232_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4059_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .A2(_1707_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4060_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .B(_2234_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4061_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(_2235_),
    .B(_2233_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q ),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4062_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q ),
    .A2(_2231_),
    .B(_2236_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4063_ (.I(_2237_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4064_ (.I0(Tile_X0Y1_E1END[3]),
    .I1(Tile_X0Y1_W1END[3]),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .Z(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4065_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ),
    .A2(_2238_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4066_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .Z(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4067_ (.A1(_0202_),
    .A2(_2240_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4068_ (.I0(_0955_),
    .I1(_1188_),
    .I2(_1730_),
    .I3(_1651_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .Z(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4069_ (.A1(_0202_),
    .A2(_2242_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4070_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4071_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ),
    .A2(_2244_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q ),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4072_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q ),
    .A2(_2239_),
    .A3(_2241_),
    .B1(_2243_),
    .B2(_2245_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4073_ (.I0(Tile_X0Y1_E1END[2]),
    .I1(Tile_X0Y1_W1END[2]),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .Z(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4074_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .Z(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4075_ (.I(_2247_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4076_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_2248_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q ),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4077_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_2246_),
    .B(_2249_),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4078_ (.A1(_0203_),
    .A2(_1026_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4079_ (.A1(_0203_),
    .A2(_0827_),
    .B(_2251_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4080_ (.A1(_0203_),
    .A2(_1707_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4081_ (.A1(_0203_),
    .A2(_1629_),
    .B(_2253_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4082_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_2254_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4083_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .Z(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4084_ (.A1(_2252_),
    .A2(_2255_),
    .B1(_2256_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q ),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4085_ (.A1(_2250_),
    .A2(_2257_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4086_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .A2(_0204_),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4087_ (.I0(Tile_X0Y1_N2MID[6]),
    .I1(Tile_X0Y1_E2MID[0]),
    .I2(Tile_X0Y1_E2MID[6]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4088_ (.I0(Tile_X0Y1_W2MID[0]),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .Z(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4089_ (.A1(_0205_),
    .A2(_2260_),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4090_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .A2(_2259_),
    .B(_2261_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4091_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(_0241_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4092_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .A2(_2258_),
    .B1(_2263_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4093_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .S1(_0204_),
    .Z(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4094_ (.A1(_0205_),
    .A2(_2265_),
    .B(_0206_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4095_ (.A1(_0206_),
    .A2(_2262_),
    .B1(_2264_),
    .B2(_2266_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4096_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1786_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4097_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1942_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4098_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1783_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4099_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1790_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4100_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1788_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4101_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1792_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4102_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1794_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4103_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1797_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4104_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1946_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4105_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1799_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4106_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1801_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4107_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1803_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4108_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1806_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4109_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1938_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4110_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1781_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4111_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1834_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4112_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1856_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4113_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1885_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4114_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1940_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4115_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A2(_1936_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4116_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4117_ (.I(Tile_X0Y1_E1END[0]),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4118_ (.I(Tile_X0Y1_E6END[0]),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4119_ (.I(Tile_X0Y1_W2END[2]),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4120_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4121_ (.I(Tile_X0Y0_S2MID[1]),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4122_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4123_ (.I(Tile_X0Y1_N2MID[4]),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4124_ (.I(Tile_X0Y0_E6END[0]),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4125_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4126_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q ),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4127_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4128_ (.I(Tile_X0Y1_E2MID[7]),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4129_ (.I(Tile_X0Y1_N2MID[1]),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4130_ (.I(Tile_X0Y1_E2MID[1]),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4131_ (.I(Tile_X0Y0_W2END[2]),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4132_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4133_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q ),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4134_ (.I(Tile_X0Y1_W2MID[1]),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4135_ (.I(Tile_X0Y0_S2MID[4]),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4136_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4137_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4138_ (.I(Tile_X0Y1_N4END[3]),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4139_ (.I(Tile_X0Y1_E2END[3]),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4140_ (.I(Tile_X0Y1_W2END[3]),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4141_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4142_ (.I(Tile_X0Y1_N2MID[0]),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4143_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4144_ (.I(Tile_X0Y1_W2MID[7]),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4145_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q ),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4146_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4147_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4148_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4149_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q ),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4150_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4151_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4152_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4153_ (.I(Tile_X0Y0_E2END[3]),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4154_ (.I(Tile_X0Y0_E6END[1]),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4155_ (.I(Tile_X0Y0_W2END[3]),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4156_ (.I(Tile_X0Y1_W1END[0]),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4157_ (.I(Tile_X0Y0_E2MID[7]),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4158_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4159_ (.I(Tile_X0Y0_S2MID[7]),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4160_ (.I(Tile_X0Y0_W2MID[7]),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4161_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4162_ (.I(Tile_X0Y0_S2END[1]),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4163_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4164_ (.I(Tile_X0Y0_SS4END[1]),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4165_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4166_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4167_ (.I(Tile_X0Y0_E2MID[3]),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4168_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4169_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4170_ (.I(Tile_X0Y0_W2MID[3]),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4171_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4172_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4173_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4174_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4175_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4176_ (.I(Tile_X0Y0_WW4END[3]),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4177_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4178_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q ),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4179_ (.I(Tile_X0Y0_S2MID[6]),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4180_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4181_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4182_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4183_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4184_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q ),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4185_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4186_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4187_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4188_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4189_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4190_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4191_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4192_ (.I(Tile_X0Y1_W1END[1]),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4193_ (.I(Tile_X0Y0_W2MID[6]),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4194_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4195_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4196_ (.I(Tile_X0Y0_EE4END[1]),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4197_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4198_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q ),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4199_ (.I(Tile_X0Y0_E2MID[4]),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4200_ (.I(Tile_X0Y0_W2MID[4]),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4201_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4202_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4203_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q ),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4204_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4205_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4206_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4207_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4208_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q ),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4209_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4210_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4211_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4212_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4213_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q ),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4214_ (.I(Tile_X0Y0_SS4END[0]),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4215_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4216_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4217_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4218_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4219_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4220_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4221_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4222_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4223_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4224_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4225_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q ),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4226_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q ),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4227_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4228_ (.I(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[4] ),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4229_ (.I(Tile_X0Y1_E2MID[0]),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4230_ (.I(Tile_X0Y0_S4END[6]),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4231_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4232_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4233_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4234_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4235_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4236_ (.I(Tile_X0Y0_SS4END[4]),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4237_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4238_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4239_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q ),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4240_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q ),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4241_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4242_ (.I(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[1] ),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4243_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4244_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4245_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q ),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4246_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4247_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4248_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q ),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4249_ (.I(Tile_X0Y0_SS4END[7]),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4250_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4251_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4252_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4253_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4254_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4255_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4256_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4257_ (.I(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[12] ),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4258_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4259_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4260_ (.I(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[10] ),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4261_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4262_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4263_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4264_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4265_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4266_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4267_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4268_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4269_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4270_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4271_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4272_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4273_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4274_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4275_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q ),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4276_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4277_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q ),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4278_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4279_ (.I(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[3] ),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4280_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4281_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q ),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4282_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4283_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4284_ (.I(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[18] ),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4285_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4286_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4287_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4288_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4289_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4290_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4291_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4292_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4293_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4294_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4295_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4296_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4297_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q ),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4298_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4299_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4300_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4301_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4302_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q ),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4303_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4304_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4305_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4306_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4307_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4308_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4309_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4310_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4311_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4312_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4313_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4314_ (.I0(_0216_),
    .I1(_0217_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4315_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4316_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ),
    .A2(_0219_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4317_ (.I0(_0208_),
    .I1(_0210_),
    .I2(_0211_),
    .I3(_0213_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4318_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ),
    .A2(_0221_),
    .B(_0220_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4319_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4320_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .A2(_0223_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4321_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4322_ (.A1(_0045_),
    .A2(_0225_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4323_ (.I0(Tile_X0Y1_E6END[1]),
    .I1(Tile_X0Y0_S2MID[3]),
    .I2(Tile_X0Y1_W2END[3]),
    .I3(Tile_X0Y1_W6END[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4324_ (.A1(_0045_),
    .A2(_0227_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4325_ (.I0(Tile_X0Y1_N1END[1]),
    .I1(Tile_X0Y1_N2END[3]),
    .I2(Tile_X0Y1_N4END[3]),
    .I3(Tile_X0Y1_E2END[3]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4326_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .A2(_0229_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4327_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ),
    .A2(_0228_),
    .A3(_0230_),
    .B1(_0224_),
    .B2(_0226_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4328_ (.I0(Tile_X0Y1_N4END[2]),
    .I1(Tile_X0Y1_E2END[2]),
    .I2(Tile_X0Y1_W2END[7]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q ),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4329_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4330_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4331_ (.A1(_0040_),
    .A2(_0233_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4332_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .A2(_0232_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4333_ (.A1(_0234_),
    .A2(_0235_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4334_ (.I0(Tile_X0Y1_N1END[2]),
    .I1(Tile_X0Y1_N2END[4]),
    .I2(Tile_X0Y1_E2END[4]),
    .I3(Tile_X0Y1_E6END[0]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4335_ (.I0(Tile_X0Y0_S2MID[4]),
    .I1(Tile_X0Y0_S4END[4]),
    .I2(Tile_X0Y1_W2END[4]),
    .I3(Tile_X0Y1_W6END[0]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4336_ (.I0(_0237_),
    .I1(_0238_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4337_ (.A1(_0041_),
    .A2(_0239_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4338_ (.A1(_0041_),
    .A2(_0239_),
    .B(_0236_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4339_ (.A1(_0234_),
    .A2(_0235_),
    .B(_0240_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4340_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4341_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ),
    .A2(_0243_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4342_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4343_ (.A1(_0036_),
    .A2(_0245_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4344_ (.A1(_0037_),
    .A2(_0244_),
    .A3(_0246_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4345_ (.I0(Tile_X0Y1_NN4END[6]),
    .I1(Tile_X0Y0_E1END[0]),
    .I2(Tile_X0Y0_EE4END[2]),
    .I3(Tile_X0Y0_E6END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4346_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ),
    .A2(_0248_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4347_ (.I0(Tile_X0Y0_S4END[2]),
    .I1(Tile_X0Y0_SS4END[2]),
    .I2(Tile_X0Y0_W2END[2]),
    .I3(Tile_X0Y0_W6END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4348_ (.A1(_0036_),
    .A2(_0250_),
    .B(_0037_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4349_ (.A1(_0249_),
    .A2(_0251_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4350_ (.A1(_0247_),
    .A2(_0252_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4351_ (.I(_0253_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4352_ (.I0(Tile_X0Y1_N2MID[1]),
    .I1(Tile_X0Y1_E2MID[1]),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .I3(Tile_X0Y1_W2MID[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q ),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4353_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I1(_0242_),
    .I2(_0254_),
    .I3(_0231_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4354_ (.A1(_0046_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4355_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ),
    .A2(_0255_),
    .B(_0256_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4356_ (.I0(Tile_X0Y0_E1END[0]),
    .I1(Tile_X0Y0_E2END[0]),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4357_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0258_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4358_ (.I0(Tile_X0Y0_S1END[0]),
    .I1(Tile_X0Y0_S2END[0]),
    .I2(Tile_X0Y0_W1END[0]),
    .I3(Tile_X0Y0_W1END[2]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4359_ (.A1(_0047_),
    .A2(_0260_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4360_ (.A1(_0257_),
    .A2(_0259_),
    .B(_0261_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4361_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4362_ (.A1(_0047_),
    .A2(_0263_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4363_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4364_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ),
    .A2(_0265_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4365_ (.A1(_0264_),
    .A2(_0266_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4366_ (.A1(_0262_),
    .A2(_0267_),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4367_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .A2(_0048_),
    .B(_0049_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4368_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .A2(_0262_),
    .A3(_0267_),
    .B(_0268_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4369_ (.A1(_0032_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4370_ (.A1(Tile_X0Y1_N2MID[7]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .B(_0049_),
    .C(_0270_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4371_ (.A1(_0269_),
    .A2(_0271_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4372_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ),
    .A2(_0269_),
    .A3(_0271_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4373_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ),
    .A2(_0269_),
    .A3(_0271_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4374_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4375_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ),
    .A2(_0275_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4376_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ),
    .A2(_0275_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4377_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4378_ (.A1(_0054_),
    .A2(_0278_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4379_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4380_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .A2(_0280_),
    .B(_0055_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4381_ (.I0(Tile_X0Y1_N2END[4]),
    .I1(Tile_X0Y1_E2END[4]),
    .I2(Tile_X0Y1_E1END[2]),
    .I3(Tile_X0Y1_E6END[0]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4382_ (.A1(_0054_),
    .A2(_0282_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4383_ (.I0(Tile_X0Y0_S2MID[4]),
    .I1(Tile_X0Y0_S4END[4]),
    .I2(Tile_X0Y1_W2END[4]),
    .I3(Tile_X0Y1_WW4END[2]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4384_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .A2(_0284_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4385_ (.A1(_0279_),
    .A2(_0281_),
    .B1(_0283_),
    .B2(_0285_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4386_ (.I0(Tile_X0Y1_N4END[1]),
    .I1(Tile_X0Y0_SS4END[5]),
    .I2(Tile_X0Y1_W2END[4]),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q ),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4387_ (.I(_0286_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4388_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ),
    .A2(_0287_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4389_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4390_ (.A1(_0051_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4391_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4392_ (.A1(_0051_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4393_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .B(_0052_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4394_ (.A1(_0290_),
    .A2(_0291_),
    .B1(_0292_),
    .B2(_0293_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4395_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .A2(_0289_),
    .B(_0294_),
    .C(_0053_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4396_ (.I0(Tile_X0Y0_S2MID[1]),
    .I1(Tile_X0Y0_S4END[5]),
    .I2(Tile_X0Y1_W2END[1]),
    .I3(Tile_X0Y1_W6END[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4397_ (.A1(Tile_X0Y1_N1END[3]),
    .A2(_0051_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4398_ (.A1(Tile_X0Y1_N2END[1]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4399_ (.A1(Tile_X0Y1_E6END[1]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4400_ (.A1(_0051_),
    .A2(Tile_X0Y1_E2END[1]),
    .B(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4401_ (.A1(_0297_),
    .A2(_0298_),
    .B1(_0300_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4402_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .A2(_0296_),
    .B(_0301_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q ),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4403_ (.A1(_0295_),
    .A2(_0302_),
    .B(_0050_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4404_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ),
    .A2(_0288_),
    .A3(_0303_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4405_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ),
    .A2(_0288_),
    .A3(_0303_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4406_ (.A1(_0273_),
    .A2(_0277_),
    .B(_0305_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4407_ (.A1(_0274_),
    .A2(_0276_),
    .B(_0304_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4408_ (.A1(Tile_X0Y1_N2MID[5]),
    .A2(_0076_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4409_ (.I0(Tile_X0Y0_E1END[1]),
    .I1(Tile_X0Y0_E2END[5]),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4410_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .A2(_0309_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4411_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .A2(_0307_),
    .A3(_0308_),
    .B(_0310_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4412_ (.I0(Tile_X0Y0_S1END[1]),
    .I1(Tile_X0Y0_S2END[5]),
    .I2(Tile_X0Y0_S1END[3]),
    .I3(Tile_X0Y0_W1END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4413_ (.I(_0312_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4414_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ),
    .A2(_0313_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4415_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0222_),
    .B1(_0311_),
    .B2(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4416_ (.I(_0315_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4417_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0222_),
    .B1(_0311_),
    .B2(_0314_),
    .C(_0075_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4418_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ),
    .A2(Tile_X0Y0_W2END[0]),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4419_ (.A1(Tile_X0Y1_NN4END[4]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4420_ (.A1(Tile_X0Y0_E6END[0]),
    .A2(_0075_),
    .B(_0077_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4421_ (.A1(_0317_),
    .A2(_0318_),
    .B1(_0319_),
    .B2(_0320_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4422_ (.A1(_0317_),
    .A2(_0318_),
    .B1(_0319_),
    .B2(_0320_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4423_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4424_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4425_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .A2(_0208_),
    .B(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4426_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4427_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .A2(_0211_),
    .B(_0326_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4428_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ),
    .A2(_0325_),
    .A3(_0327_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4429_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ),
    .A2(_0328_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4430_ (.A1(_0081_),
    .A2(_0323_),
    .B(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4431_ (.I0(_0255_),
    .I1(Tile_X0Y1_N2MID[2]),
    .I2(Tile_X0Y1_N4END[6]),
    .I3(Tile_X0Y0_E2END[2]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4432_ (.A1(_0081_),
    .A2(_0331_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4433_ (.I0(Tile_X0Y0_E6END[0]),
    .I1(Tile_X0Y0_W2END[2]),
    .I2(Tile_X0Y0_S2END[2]),
    .I3(Tile_X0Y0_WW4END[3]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4434_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ),
    .A2(_0333_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4435_ (.A1(_0332_),
    .A2(_0334_),
    .B(_0330_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4436_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4437_ (.A1(_0082_),
    .A2(_0335_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4438_ (.A1(_0322_),
    .A2(_0336_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4439_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4440_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4441_ (.A1(_0072_),
    .A2(_0339_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4442_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .A2(_0338_),
    .B(_0073_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4443_ (.I0(Tile_X0Y1_E6END[0]),
    .I1(Tile_X0Y0_S2MID[4]),
    .I2(Tile_X0Y1_W2END[4]),
    .I3(Tile_X0Y1_W6END[0]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4444_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .A2(_0342_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4445_ (.I0(Tile_X0Y1_N2END[4]),
    .I1(Tile_X0Y1_E1END[2]),
    .I2(Tile_X0Y1_N4END[0]),
    .I3(Tile_X0Y1_E2END[4]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4446_ (.A1(_0072_),
    .A2(_0344_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4447_ (.A1(_0340_),
    .A2(_0341_),
    .B1(_0343_),
    .B2(_0345_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4448_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .I1(Tile_X0Y0_E2MID[3]),
    .I2(Tile_X0Y0_S2MID[3]),
    .I3(Tile_X0Y0_W2MID[3]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q ),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4449_ (.I(_0346_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4450_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ),
    .A2(_0347_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4451_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .B(_0348_),
    .C(_0082_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4452_ (.I(_0349_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4453_ (.A1(_0337_),
    .A2(_0349_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4454_ (.A1(_0322_),
    .A2(_0336_),
    .B(_0350_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4455_ (.A1(_0078_),
    .A2(Tile_X0Y0_S2MID[6]),
    .B(_0079_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4456_ (.A1(Tile_X0Y1_W1END[0]),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4457_ (.A1(Tile_X0Y1_W1END[2]),
    .A2(_0078_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4458_ (.A1(_0352_),
    .A2(_0353_),
    .B1(_0354_),
    .B2(_0355_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4459_ (.I0(Tile_X0Y1_N1END[2]),
    .I1(Tile_X0Y1_E1END[2]),
    .I2(Tile_X0Y1_N2END[6]),
    .I3(Tile_X0Y1_E2END[6]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4460_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .A2(_0357_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4461_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .A2(_0358_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4462_ (.A1(_0356_),
    .A2(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4463_ (.A1(_0078_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4464_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .B(_0079_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4465_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4466_ (.A1(_0078_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4467_ (.A1(_0361_),
    .A2(_0362_),
    .B1(_0363_),
    .B2(_0364_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4468_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4469_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .A2(_0366_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4470_ (.A1(_0084_),
    .A2(_0367_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4471_ (.A1(_0365_),
    .A2(_0368_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4472_ (.A1(_0360_),
    .A2(_0369_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4473_ (.A1(_0356_),
    .A2(_0359_),
    .B1(_0365_),
    .B2(_0368_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4474_ (.A1(Tile_X0Y0_E2MID[5]),
    .A2(_0085_),
    .B(_0086_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4475_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ),
    .A2(Tile_X0Y0_S2MID[5]),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4476_ (.A1(_0085_),
    .A2(Tile_X0Y0_W2MID[5]),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4477_ (.A1(_0370_),
    .A2(_0371_),
    .B1(_0372_),
    .B2(_0373_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4478_ (.A1(_0370_),
    .A2(_0371_),
    .B1(_0372_),
    .B2(_0373_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4479_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4480_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ),
    .A2(_0376_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4481_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4482_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4483_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .A2(_0210_),
    .B(_0379_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4484_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .A2(_0213_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4485_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .B(_0381_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4486_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ),
    .A2(_0382_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4487_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ),
    .A2(_0378_),
    .B1(_0380_),
    .B2(_0383_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4488_ (.I(_0384_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4489_ (.A1(_0274_),
    .A2(_0276_),
    .B(_0304_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4490_ (.A1(_0273_),
    .A2(_0277_),
    .B(_0305_),
    .C(_0056_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4491_ (.A1(Tile_X0Y1_N2MID[3]),
    .A2(_0056_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4492_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .A2(_0388_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4493_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .A2(Tile_X0Y1_N4END[7]),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4494_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .A2(_0057_),
    .B(_0390_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4495_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .A2(_0391_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4496_ (.A1(_0387_),
    .A2(_0389_),
    .B1(_0391_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4497_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .A2(_0386_),
    .A3(_0388_),
    .B(_0392_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4498_ (.I0(Tile_X0Y0_E6END[1]),
    .I1(Tile_X0Y0_S2END[3]),
    .I2(Tile_X0Y0_W2END[3]),
    .I3(Tile_X0Y0_W6END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4499_ (.I(_0395_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4500_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ),
    .A2(_0396_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4501_ (.I(_0397_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4502_ (.A1(_0393_),
    .A2(_0398_),
    .B(_0384_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4503_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4504_ (.A1(_0087_),
    .A2(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4505_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4506_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ),
    .A2(_0401_),
    .B(_0088_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4507_ (.I0(Tile_X0Y1_N2MID[2]),
    .I1(Tile_X0Y0_E1END[0]),
    .I2(Tile_X0Y1_N4END[6]),
    .I3(Tile_X0Y0_E2END[2]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4508_ (.A1(_0087_),
    .A2(_0403_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4509_ (.I0(Tile_X0Y0_E6END[0]),
    .I1(Tile_X0Y0_W2END[2]),
    .I2(Tile_X0Y0_S2END[2]),
    .I3(Tile_X0Y0_W6END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4510_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ),
    .A2(_0405_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q ),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4511_ (.A1(_0400_),
    .A2(_0402_),
    .B1(_0404_),
    .B2(_0406_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4512_ (.I0(Tile_X0Y1_NN4END[7]),
    .I1(Tile_X0Y0_WW4END[0]),
    .I2(Tile_X0Y0_S4END[3]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q ),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4513_ (.I(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4514_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4515_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ),
    .A2(_0408_),
    .B(_0409_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4516_ (.A1(_0375_),
    .A2(_0377_),
    .B(_0410_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4517_ (.I(_0411_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4518_ (.A1(_0375_),
    .A2(_0377_),
    .B(_0410_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4519_ (.A1(Tile_X0Y0_S2MID[7]),
    .A2(_0094_),
    .B(_0095_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4520_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .A2(Tile_X0Y1_W1END[1]),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4521_ (.A1(_0094_),
    .A2(Tile_X0Y1_W1END[3]),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4522_ (.A1(_0413_),
    .A2(_0414_),
    .B1(_0415_),
    .B2(_0416_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4523_ (.I0(Tile_X0Y1_N1END[3]),
    .I1(Tile_X0Y1_N2END[7]),
    .I2(Tile_X0Y1_E1END[3]),
    .I3(Tile_X0Y1_E2END[7]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4524_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .A2(_0418_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4525_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0419_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4526_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0218_),
    .B1(_0417_),
    .B2(_0420_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4527_ (.I(_0421_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4528_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4529_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4530_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4531_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4532_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .A2(_0425_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4533_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .A2(_0426_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4534_ (.A1(_0024_),
    .A2(_0424_),
    .B(_0427_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4535_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .A2(_0022_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4536_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .A2(Tile_X0Y0_S2MID[2]),
    .B(_0429_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4537_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .A2(_0023_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4538_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .A2(Tile_X0Y1_W6END[0]),
    .B(_0431_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4539_ (.A1(_0024_),
    .A2(_0430_),
    .A3(_0432_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4540_ (.I0(Tile_X0Y1_N2END[2]),
    .I1(Tile_X0Y1_N4END[2]),
    .I2(Tile_X0Y1_E1END[0]),
    .I3(Tile_X0Y1_E2END[2]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4541_ (.A1(_0024_),
    .A2(_0434_),
    .B(_0433_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4542_ (.A1(_0428_),
    .A2(_0435_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4543_ (.I0(Tile_X0Y1_NN4END[3]),
    .I1(Tile_X0Y1_WW4END[0]),
    .I2(Tile_X0Y0_S4END[7]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q ),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4544_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4545_ (.I(_0437_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4546_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4547_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .A2(_0439_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4548_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .A2(_0438_),
    .B(_0440_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4549_ (.I0(Tile_X0Y1_N1END[1]),
    .I1(Tile_X0Y1_N2END[3]),
    .I2(Tile_X0Y1_E2END[3]),
    .I3(Tile_X0Y1_E6END[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4550_ (.I0(Tile_X0Y0_S2MID[3]),
    .I1(Tile_X0Y1_W2END[3]),
    .I2(Tile_X0Y0_S4END[7]),
    .I3(Tile_X0Y1_W6END[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4551_ (.I0(_0442_),
    .I1(_0443_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4552_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ),
    .A2(_0444_),
    .B(_0441_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4553_ (.I(_0445_),
    .ZN(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4554_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4555_ (.I(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4556_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4557_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4558_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(_0447_),
    .B(_0449_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q ),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4559_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .I1(Tile_X0Y0_E1END[2]),
    .I2(Tile_X0Y1_N2MID[6]),
    .I3(Tile_X0Y0_E2END[6]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4560_ (.I0(Tile_X0Y0_S1END[2]),
    .I1(Tile_X0Y0_S2END[6]),
    .I2(Tile_X0Y0_W1END[0]),
    .I3(Tile_X0Y0_W1END[2]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4561_ (.I0(_0451_),
    .I1(_0452_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4562_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q ),
    .A2(_0453_),
    .B(_0450_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4563_ (.I(_0454_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4564_ (.I0(Tile_X0Y1_N2MID[5]),
    .I1(Tile_X0Y1_E2MID[5]),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .I3(Tile_X0Y1_W2MID[5]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q ),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4565_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ),
    .I2(_0455_),
    .I3(_0436_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q ),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4566_ (.I0(_0456_),
    .I1(Tile_X0Y0_E1END[3]),
    .I2(Tile_X0Y1_N2MID[7]),
    .I3(Tile_X0Y0_E2END[7]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4567_ (.I0(Tile_X0Y0_S1END[3]),
    .I1(Tile_X0Y0_W1END[1]),
    .I2(Tile_X0Y0_S2END[7]),
    .I3(Tile_X0Y0_W1END[3]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4568_ (.I0(_0457_),
    .I1(_0458_),
    .I2(_0422_),
    .I3(_0423_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4569_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .I1(Tile_X0Y0_E2MID[6]),
    .I2(Tile_X0Y0_S2MID[6]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q ),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4570_ (.A1(Tile_X0Y0_E2END[2]),
    .A2(_0031_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4571_ (.A1(Tile_X0Y1_N4END[6]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4572_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ),
    .A2(_0460_),
    .A3(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4573_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ),
    .A2(_0460_),
    .A3(_0461_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4574_ (.A1(_0394_),
    .A2(_0397_),
    .B(_0031_),
    .C(_0385_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4575_ (.A1(_0393_),
    .A2(_0398_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ),
    .C(_0384_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4576_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ),
    .A2(Tile_X0Y0_W2END[7]),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4577_ (.I(_0466_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4578_ (.A1(_0464_),
    .A2(_0466_),
    .B(_0463_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4579_ (.A1(_0465_),
    .A2(_0467_),
    .B(_0026_),
    .C(_0462_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4580_ (.A1(_0464_),
    .A2(_0466_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ),
    .C(_0463_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4581_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4582_ (.A1(_0029_),
    .A2(_0471_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4583_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4584_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ),
    .A2(_0473_),
    .B(_0030_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4585_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .I1(Tile_X0Y1_N4END[4]),
    .I2(Tile_X0Y1_N2MID[4]),
    .I3(Tile_X0Y0_E2END[4]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4586_ (.A1(_0029_),
    .A2(_0475_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4587_ (.I0(Tile_X0Y0_E6END[0]),
    .I1(Tile_X0Y0_S2END[4]),
    .I2(Tile_X0Y0_W2END[4]),
    .I3(Tile_X0Y0_W6END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4588_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ),
    .A2(_0477_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q ),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4589_ (.A1(_0472_),
    .A2(_0474_),
    .B1(_0476_),
    .B2(_0478_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4590_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4591_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ),
    .A2(_0479_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4592_ (.I(_0480_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4593_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .I1(Tile_X0Y0_S2MID[1]),
    .I2(Tile_X0Y0_E2MID[1]),
    .I3(Tile_X0Y0_W2MID[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q ),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4594_ (.I(_0482_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4595_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4596_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ),
    .A2(_0484_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4597_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ),
    .A2(_0483_),
    .B(_0484_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4598_ (.A1(_0026_),
    .A2(_0482_),
    .B(_0485_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4599_ (.A1(_0470_),
    .A2(_0480_),
    .B(_0486_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4600_ (.A1(_0469_),
    .A2(_0481_),
    .B(_0487_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4601_ (.A1(_0470_),
    .A2(_0480_),
    .B(_0486_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4602_ (.A1(_0469_),
    .A2(_0481_),
    .B(_0487_),
    .C(_0020_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4603_ (.A1(_0020_),
    .A2(Tile_X0Y0_S2MID[0]),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4604_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_0492_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4605_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_0492_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4606_ (.A1(_0020_),
    .A2(Tile_X0Y1_W1END[2]),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4607_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .A2(Tile_X0Y1_W1END[0]),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4608_ (.A1(_0495_),
    .A2(_0496_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4609_ (.A1(_0491_),
    .A2(_0493_),
    .B(_0497_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4610_ (.A1(_0490_),
    .A2(_0494_),
    .B1(_0495_),
    .B2(_0496_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4611_ (.I0(Tile_X0Y1_N1END[0]),
    .I1(Tile_X0Y1_E1END[0]),
    .I2(Tile_X0Y1_N2END[0]),
    .I3(Tile_X0Y1_EE4END[0]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4612_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .A2(_0500_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4613_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ),
    .A2(_0501_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4614_ (.I(_0502_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4615_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4616_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4617_ (.I(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4618_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .A2(_0506_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4619_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .A2(_0504_),
    .B(_0507_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4620_ (.I(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4621_ (.A1(_0498_),
    .A2(_0503_),
    .B(_0508_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4622_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ),
    .I1(Tile_X0Y0_S2MID[7]),
    .I2(Tile_X0Y0_E2MID[7]),
    .I3(Tile_X0Y0_W2MID[7]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q ),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4623_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4624_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4625_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .A2(_0208_),
    .B(_0512_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4626_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4627_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .A2(_0211_),
    .B(_0514_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4628_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(_0513_),
    .A3(_0515_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4629_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0516_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4630_ (.A1(_0110_),
    .A2(_0511_),
    .B(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4631_ (.I0(_0306_),
    .I1(Tile_X0Y0_E1END[1]),
    .I2(Tile_X0Y1_N2MID[5]),
    .I3(Tile_X0Y0_E2END[5]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4632_ (.I0(Tile_X0Y0_S1END[1]),
    .I1(Tile_X0Y0_W1END[1]),
    .I2(Tile_X0Y0_S2END[5]),
    .I3(Tile_X0Y0_W1END[3]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4633_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(_0520_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4634_ (.A1(_0110_),
    .A2(_0519_),
    .B(_0521_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4635_ (.A1(_0518_),
    .A2(_0522_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4636_ (.I0(Tile_X0Y1_N4END[7]),
    .I1(Tile_X0Y0_S4END[3]),
    .I2(Tile_X0Y0_EE4END[0]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q ),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4637_ (.I0(Tile_X0Y1_N2MID[7]),
    .I1(Tile_X0Y0_S2END[7]),
    .I2(Tile_X0Y0_E2END[7]),
    .I3(Tile_X0Y0_WW4END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q ),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4638_ (.I(_0524_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4639_ (.I0(_0459_),
    .I1(_0510_),
    .I2(_0524_),
    .I3(_0523_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q ),
    .Z(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4640_ (.A1(_0162_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4641_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[14] ),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4642_ (.A1(_0163_),
    .A2(_0526_),
    .A3(_0527_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4643_ (.A1(_0163_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[14] ),
    .B(_0528_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4644_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4645_ (.A1(_0091_),
    .A2(_0530_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4646_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4647_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ),
    .A2(_0532_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4648_ (.I0(Tile_X0Y0_E6END[1]),
    .I1(Tile_X0Y0_S2END[3]),
    .I2(Tile_X0Y0_W2END[3]),
    .I3(Tile_X0Y0_WW4END[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4649_ (.A1(_0091_),
    .A2(_0534_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4650_ (.I0(Tile_X0Y1_N2MID[3]),
    .I1(Tile_X0Y1_N4END[7]),
    .I2(Tile_X0Y0_E1END[1]),
    .I3(Tile_X0Y0_E2END[3]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4651_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ),
    .A2(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4652_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ),
    .A2(_0535_),
    .A3(_0537_),
    .B1(_0531_),
    .B2(_0533_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4653_ (.I0(Tile_X0Y1_NN4END[7]),
    .I1(Tile_X0Y0_S2END[6]),
    .I2(Tile_X0Y0_E2END[6]),
    .I3(Tile_X0Y0_W2END[6]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q ),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4654_ (.I0(Tile_X0Y0_E2END[3]),
    .I1(Tile_X0Y0_WW4END[2]),
    .I2(Tile_X0Y0_SS4END[3]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q ),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4655_ (.I0(_0538_),
    .I1(_0539_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4656_ (.A1(_0061_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q ),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4657_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ),
    .B(_0541_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4658_ (.A1(_0064_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4659_ (.A1(Tile_X0Y0_S2MID[7]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q ),
    .C(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4660_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ),
    .A2(_0542_),
    .A3(_0544_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4661_ (.I0(Tile_X0Y0_E2MID[6]),
    .I1(Tile_X0Y0_W2MID[6]),
    .I2(Tile_X0Y0_S2MID[6]),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q ),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4662_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ),
    .A2(_0546_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4663_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q ),
    .A2(_0547_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4664_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q ),
    .A2(_0540_),
    .B1(_0545_),
    .B2(_0548_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4665_ (.I(_0549_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4666_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[4] ),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4667_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .A2(_0549_),
    .B(_0550_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4668_ (.I(_0551_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4669_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4670_ (.A1(_0108_),
    .A2(_0553_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4671_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4672_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ),
    .A2(_0555_),
    .B(_0109_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4673_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .I1(Tile_X0Y0_E2END[4]),
    .I2(Tile_X0Y1_N2MID[4]),
    .I3(Tile_X0Y0_E6END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4674_ (.A1(_0108_),
    .A2(_0557_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4675_ (.I0(Tile_X0Y0_S2END[4]),
    .I1(Tile_X0Y0_W2END[4]),
    .I2(Tile_X0Y0_S4END[0]),
    .I3(Tile_X0Y0_W6END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4676_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ),
    .A2(_0559_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4677_ (.A1(_0554_),
    .A2(_0556_),
    .B1(_0558_),
    .B2(_0560_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4678_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4679_ (.A1(_0106_),
    .A2(_0562_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4680_ (.I0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .I1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .I2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .I3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4681_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .A2(_0564_),
    .B(_0107_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4682_ (.I0(Tile_X0Y1_N2END[1]),
    .I1(Tile_X0Y1_N4END[1]),
    .I2(Tile_X0Y1_E1END[3]),
    .I3(Tile_X0Y1_E2END[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4683_ (.A1(_0106_),
    .A2(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4684_ (.I0(Tile_X0Y1_E6END[1]),
    .I1(Tile_X0Y1_W2END[1]),
    .I2(Tile_X0Y0_SS4END[5]),
    .I3(Tile_X0Y1_W6END[1]),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4685_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .A2(_0568_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q ),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4686_ (.A1(_0563_),
    .A2(_0565_),
    .B1(_0567_),
    .B2(_0569_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4687_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .I1(Tile_X0Y0_E2MID[0]),
    .I2(Tile_X0Y0_S2MID[0]),
    .I3(_0561_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q ),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4688_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .I1(Tile_X0Y0_S2MID[1]),
    .I2(Tile_X0Y0_E2MID[1]),
    .I3(Tile_X0Y0_W2MID[1]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q ),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4689_ (.I(_0571_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4690_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ),
    .A2(_0572_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q ),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4691_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ),
    .A2(_0570_),
    .B(_0573_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4692_ (.I0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .I1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .I2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .I3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4693_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .A2(_0210_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4694_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .B(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4695_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .A2(_0214_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4696_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .B(_0578_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4697_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .A2(_0577_),
    .B(_0579_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4698_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ),
    .A2(_0575_),
    .B(_0580_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4699_ (.I0(_0255_),
    .I1(Tile_X0Y1_N2MID[2]),
    .I2(Tile_X0Y0_E2END[2]),
    .I3(Tile_X0Y0_E6END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4700_ (.I0(Tile_X0Y0_S2END[2]),
    .I1(Tile_X0Y0_W2END[2]),
    .I2(Tile_X0Y0_S4END[2]),
    .I3(Tile_X0Y0_W6END[0]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4701_ (.I(_0583_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4702_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ),
    .A2(_0584_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4703_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ),
    .A2(_0582_),
    .B(_0585_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4704_ (.A1(_0581_),
    .A2(_0586_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4705_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4706_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ),
    .A2(_0587_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4707_ (.A1(Tile_X0Y0_S4END[0]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q ),
    .C(_0588_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4708_ (.A1(_0028_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q ),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4709_ (.A1(Tile_X0Y1_N4END[4]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ),
    .B(_0590_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4710_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ),
    .A2(_0589_),
    .A3(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4711_ (.I0(Tile_X0Y1_N2MID[0]),
    .I1(Tile_X0Y0_E2END[0]),
    .I2(Tile_X0Y0_S2END[0]),
    .I3(Tile_X0Y0_WW4END[3]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q ),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4712_ (.I(_0593_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4713_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ),
    .A2(_0593_),
    .B(_0592_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q ),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4714_ (.A1(_0574_),
    .A2(_0595_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4715_ (.I(_0596_),
    .ZN(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4716_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[7] ),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4717_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(_0596_),
    .B(_0597_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4718_ (.I(_0598_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4719_ (.A1(_0551_),
    .A2(_0598_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4720_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ),
    .A2(_0253_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4721_ (.A1(Tile_X0Y0_W6END[1]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q ),
    .C(_0601_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4722_ (.A1(Tile_X0Y1_N4END[5]),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4723_ (.A1(_0058_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q ),
    .C(_0603_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4724_ (.A1(_0105_),
    .A2(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4725_ (.I0(Tile_X0Y1_N2MID[4]),
    .I1(Tile_X0Y0_S2END[4]),
    .I2(Tile_X0Y0_EE4END[0]),
    .I3(Tile_X0Y0_W2END[4]),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q ),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4726_ (.I(_0606_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4727_ (.A1(_0602_),
    .A2(_0605_),
    .B1(_0607_),
    .B2(_0105_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4728_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4729_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4730_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4731_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4732_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4733_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4734_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4735_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4736_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4737_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4738_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4739_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4740_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4741_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4742_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4743_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4744_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4745_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4746_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4747_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4748_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4749_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4750_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4751_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4752_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4753_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4754_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4755_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4756_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4757_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4758_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4759_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4760_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4761_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4762_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4763_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4764_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4765_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4766_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4767_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4768_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4769_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4770_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4771_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4772_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4773_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4774_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4775_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4776_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4777_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4778_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4779_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4780_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4781_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4782_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4783_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4784_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4785_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4786_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4787_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4788_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4789_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4790_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4791_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4792_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4793_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4794_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4795_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4796_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4797_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4798_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4799_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4800_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4801_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4802_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4803_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4804_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4805_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4806_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4807_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4808_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4809_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4810_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4811_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4812_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4813_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4814_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4815_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4816_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4817_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4818_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4819_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4820_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4821_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4822_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4823_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4824_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4825_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4826_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4827_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4828_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4829_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4830_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4831_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4832_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4833_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4834_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4835_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4836_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4837_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4838_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4839_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4840_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4841_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4842_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4843_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4844_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4845_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4846_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4847_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4848_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4849_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4850_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4851_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4852_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4853_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4854_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4855_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4856_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4857_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4858_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4859_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4860_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4861_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4862_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4863_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4864_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4865_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4866_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4867_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4868_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4869_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4870_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4871_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4872_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4873_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4874_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4875_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4876_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4877_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4878_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4879_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4880_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4881_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4882_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4883_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4884_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4885_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4886_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4887_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4888_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4889_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4890_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4891_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4892_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4893_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4894_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4895_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4896_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4897_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4898_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4899_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4900_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4901_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4902_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4903_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4904_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4905_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4906_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4907_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4908_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4909_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4910_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4911_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4912_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4913_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4914_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4915_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4916_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4917_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4918_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4919_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4920_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4921_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4922_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4923_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4924_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4925_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4926_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4927_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4928_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4929_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4930_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4931_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4932_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4933_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4934_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4935_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4936_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4937_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4938_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4939_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4940_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4941_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4942_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4943_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4944_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4945_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4946_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4947_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4948_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4949_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4950_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4951_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4952_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4953_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4954_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4955_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4956_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4957_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4958_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4959_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4960_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4961_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4962_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4963_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4964_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4965_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4966_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4967_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4968_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4969_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4970_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4971_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4972_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4973_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4974_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4975_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4976_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4977_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4978_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4979_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4980_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4981_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4982_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4983_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4984_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4985_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4986_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4987_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4988_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4989_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4990_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4991_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4992_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4993_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4994_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4995_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4996_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4997_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4998_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _4999_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5000_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5001_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5002_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5003_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5004_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5005_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5006_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5007_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5008_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5009_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5010_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5011_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5012_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5013_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5014_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5015_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5016_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5017_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5018_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5019_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5020_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5021_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5022_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5023_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5024_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5025_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5026_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5027_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5028_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5029_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5030_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5031_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5032_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5033_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5034_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5035_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5036_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5037_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5038_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5039_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5040_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5041_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5042_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5043_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5044_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5045_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5046_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5047_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5048_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5049_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5050_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5051_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5052_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5053_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5054_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5055_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5056_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5057_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5058_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5059_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5060_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5061_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5062_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5063_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5064_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5065_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5066_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5067_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5068_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5069_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5070_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5071_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5072_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5073_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5074_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5075_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5076_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5077_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5078_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5079_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5080_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5081_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5082_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5083_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5084_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5085_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5086_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5087_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5088_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5089_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5090_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5091_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5092_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5093_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5094_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5095_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5096_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5097_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5098_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5099_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5100_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5101_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5102_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5103_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5104_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5105_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5106_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5107_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5108_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5109_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5110_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5111_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5112_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5113_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5114_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5115_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5116_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5117_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5118_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5119_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5120_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5121_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5122_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5123_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5124_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5125_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5126_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5127_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5128_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5129_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5130_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5131_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5132_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5133_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5134_ (.D(_0000_),
    .CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5135_ (.D(_0001_),
    .CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5136_ (.D(_0002_),
    .CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5137_ (.D(_0003_),
    .CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5138_ (.D(_0004_),
    .CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5139_ (.D(_0005_),
    .CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5140_ (.D(_0006_),
    .CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5141_ (.D(_0007_),
    .CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5142_ (.D(_0008_),
    .CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5143_ (.D(_0009_),
    .CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5144_ (.D(_0010_),
    .CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5145_ (.D(_0011_),
    .CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5146_ (.D(_0012_),
    .CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5147_ (.D(_0013_),
    .CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5148_ (.D(_0014_),
    .CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5149_ (.D(_0015_),
    .CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5150_ (.D(_0016_),
    .CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5151_ (.D(_0017_),
    .CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5152_ (.D(_0018_),
    .CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5153_ (.D(_0019_),
    .CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5154_ (.D(\Tile_X0Y1_DSP_bot.A0 ),
    .CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5155_ (.D(\Tile_X0Y1_DSP_bot.A1 ),
    .CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5156_ (.D(\Tile_X0Y1_DSP_bot.A2 ),
    .CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5157_ (.D(\Tile_X0Y1_DSP_bot.A3 ),
    .CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5158_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X ),
    .CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5159_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X ),
    .CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5160_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ),
    .CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5161_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X ),
    .CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5162_ (.D(\Tile_X0Y1_DSP_bot.B0 ),
    .CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5163_ (.D(\Tile_X0Y1_DSP_bot.B1 ),
    .CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5164_ (.D(\Tile_X0Y1_DSP_bot.B2 ),
    .CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5165_ (.D(\Tile_X0Y1_DSP_bot.B3 ),
    .CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5166_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X ),
    .CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5167_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ),
    .CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5168_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X ),
    .CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5169_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X ),
    .CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5170_ (.D(\Tile_X0Y1_DSP_bot.C0 ),
    .CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5171_ (.D(\Tile_X0Y1_DSP_bot.C1 ),
    .CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5172_ (.D(\Tile_X0Y1_DSP_bot.C2 ),
    .CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5173_ (.D(\Tile_X0Y1_DSP_bot.C3 ),
    .CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5174_ (.D(\Tile_X0Y1_DSP_bot.C4 ),
    .CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5175_ (.D(\Tile_X0Y1_DSP_bot.C5 ),
    .CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5176_ (.D(\Tile_X0Y1_DSP_bot.C6 ),
    .CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5177_ (.D(\Tile_X0Y1_DSP_bot.C7 ),
    .CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5178_ (.D(\Tile_X0Y1_DSP_bot.C8 ),
    .CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5179_ (.D(\Tile_X0Y1_DSP_bot.C9 ),
    .CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5180_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ),
    .CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5181_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X ),
    .CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5182_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ),
    .CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5183_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ),
    .CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5184_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ),
    .CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5185_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ),
    .CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5186_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ),
    .CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5187_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ),
    .CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5188_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ),
    .CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _5189_ (.D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ),
    .CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[19] ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5190_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5191_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5192_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5193_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5194_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5195_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5196_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5197_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5198_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5199_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5200_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5201_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5202_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5203_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5204_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5205_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5206_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5207_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5208_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5209_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5210_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5211_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5212_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5213_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5214_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5215_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5216_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5217_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5218_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5219_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5220_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5221_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5222_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5223_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5224_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5225_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5226_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5227_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5228_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5229_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5230_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5231_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5232_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5233_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5234_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5235_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5236_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5237_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5238_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5239_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5240_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5241_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5242_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5243_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5244_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5245_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5246_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5247_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5248_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5249_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5250_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5251_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5252_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5253_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5254_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5255_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5256_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5257_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5258_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5259_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5260_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5261_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5262_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5263_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5264_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5265_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5266_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5267_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5268_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5269_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5270_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5271_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5272_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5273_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5274_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5275_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5276_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5277_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5278_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5279_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5280_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5281_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5282_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5283_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5284_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5285_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5286_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5287_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5288_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5289_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5290_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5291_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5292_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5293_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5294_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5295_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5296_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5297_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5298_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5299_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5300_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5301_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5302_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5303_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5304_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5305_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5306_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5307_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5308_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5309_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5310_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5311_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5312_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5313_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5314_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5315_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5316_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5317_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5318_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5319_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5320_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5321_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5322_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5323_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5324_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5325_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5326_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5327_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5328_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5329_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5330_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5331_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5332_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5333_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5334_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5335_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5336_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5337_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5338_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5339_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5340_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5341_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5342_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5343_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5344_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5345_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5346_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5347_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5348_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5349_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5350_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5351_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5352_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5353_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5354_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5355_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5356_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5357_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5358_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5359_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5360_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5361_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5362_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5363_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5364_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5365_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5366_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5367_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5368_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5369_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5370_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5371_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5372_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5373_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5374_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5375_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5376_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5377_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5378_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5379_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5380_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5381_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5382_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5383_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5384_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5385_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5386_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5387_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5388_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5389_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5390_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5391_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5392_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5393_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5394_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5395_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5396_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5397_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5398_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5399_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5400_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5401_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5402_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5403_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5404_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5405_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5406_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5407_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5408_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5409_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5410_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5411_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5412_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5413_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5414_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5415_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5416_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5417_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5418_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5419_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5420_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5421_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5422_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5423_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5424_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5425_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5426_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5427_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5428_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5429_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5430_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5431_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5432_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5433_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5434_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5435_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5436_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5437_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5438_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5439_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5440_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5441_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5442_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5443_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5444_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5445_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5446_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5447_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5448_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5449_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5450_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5451_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5452_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5453_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5454_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5455_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5456_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5457_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5458_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5459_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5460_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5461_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5462_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5463_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5464_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5465_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5466_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5467_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5468_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5469_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5470_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5471_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5472_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5473_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5474_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5475_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5476_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5477_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5478_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5479_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5480_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5481_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5482_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5483_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5484_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5485_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5486_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5487_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5488_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5489_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5490_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5491_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5492_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5493_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5494_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5495_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5496_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5497_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5498_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5499_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5500_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5501_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5502_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5503_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5504_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5505_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5506_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5507_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5508_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5509_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5510_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5511_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5512_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5513_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5514_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5515_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5516_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5517_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5518_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5519_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5520_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5521_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5522_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5523_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5524_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5525_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5526_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5527_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5528_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5529_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5530_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5531_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5532_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5533_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5534_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5535_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5536_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5537_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5538_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5539_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5540_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5541_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[10]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5542_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5543_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5544_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5545_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5546_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5547_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5548_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5549_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5550_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5551_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5552_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5553_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5554_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5555_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5556_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5557_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5558_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5559_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5560_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5561_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5562_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5563_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5564_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5565_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5566_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5567_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5568_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5569_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5570_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5571_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5572_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5573_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[11]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5574_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5575_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5576_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5577_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5578_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5579_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5580_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5581_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5582_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5583_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5584_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5585_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5586_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5587_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5588_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5589_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5590_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5591_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5592_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5593_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5594_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5595_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5596_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5597_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5598_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5599_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5600_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5601_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5602_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5603_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5604_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _5605_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[12]),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5606_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 ),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5607_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 ),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5608_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 ),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5609_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 ),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5610_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5611_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5612_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5613_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5614_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5615_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5616_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5617_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5618_ (.I(Tile_X0Y0_E2MID[0]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5619_ (.I(Tile_X0Y0_E2MID[1]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5620_ (.I(Tile_X0Y0_E2MID[2]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5621_ (.I(Tile_X0Y0_E2MID[3]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5622_ (.I(Tile_X0Y0_E2MID[4]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5623_ (.I(Tile_X0Y0_E2MID[5]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5624_ (.I(Tile_X0Y0_E2MID[6]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5625_ (.I(Tile_X0Y0_E2MID[7]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5626_ (.I(Tile_X0Y0_E6END[2]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5627_ (.I(Tile_X0Y0_E6END[3]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5628_ (.I(Tile_X0Y0_E6END[4]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5629_ (.I(Tile_X0Y0_E6END[5]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5630_ (.I(Tile_X0Y0_E6END[6]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5631_ (.I(Tile_X0Y0_E6END[7]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5632_ (.I(Tile_X0Y0_E6END[8]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5633_ (.I(Tile_X0Y0_E6END[9]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5634_ (.I(Tile_X0Y0_E6END[10]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5635_ (.I(Tile_X0Y0_E6END[11]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5636_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 ),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5637_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 ),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5638_ (.I(Tile_X0Y0_EE4END[4]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5639_ (.I(Tile_X0Y0_EE4END[5]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5640_ (.I(Tile_X0Y0_EE4END[6]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5641_ (.I(Tile_X0Y0_EE4END[7]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5642_ (.I(Tile_X0Y0_EE4END[8]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5643_ (.I(Tile_X0Y0_EE4END[9]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5644_ (.I(Tile_X0Y0_EE4END[10]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5645_ (.I(Tile_X0Y0_EE4END[11]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5646_ (.I(Tile_X0Y0_EE4END[12]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5647_ (.I(Tile_X0Y0_EE4END[13]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5648_ (.I(Tile_X0Y0_EE4END[14]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5649_ (.I(Tile_X0Y0_EE4END[15]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5650_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 ),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5651_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 ),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5652_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 ),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5653_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 ),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5654_ (.I(Tile_X0Y0_FrameData[0]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5655_ (.I(Tile_X0Y0_FrameData[1]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5656_ (.I(Tile_X0Y0_FrameData[2]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5657_ (.I(Tile_X0Y0_FrameData[3]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5658_ (.I(Tile_X0Y0_FrameData[4]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5659_ (.I(Tile_X0Y0_FrameData[5]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5660_ (.I(Tile_X0Y0_FrameData[6]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5661_ (.I(Tile_X0Y0_FrameData[7]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5662_ (.I(Tile_X0Y0_FrameData[8]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5663_ (.I(Tile_X0Y0_FrameData[9]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5664_ (.I(Tile_X0Y0_FrameData[10]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5665_ (.I(Tile_X0Y0_FrameData[11]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5666_ (.I(Tile_X0Y0_FrameData[12]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5667_ (.I(Tile_X0Y0_FrameData[13]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5668_ (.I(Tile_X0Y0_FrameData[14]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5669_ (.I(Tile_X0Y0_FrameData[15]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5670_ (.I(Tile_X0Y0_FrameData[16]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5671_ (.I(Tile_X0Y0_FrameData[17]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5672_ (.I(Tile_X0Y0_FrameData[18]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5673_ (.I(Tile_X0Y0_FrameData[19]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5674_ (.I(Tile_X0Y0_FrameData[20]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5675_ (.I(Tile_X0Y0_FrameData[21]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5676_ (.I(Tile_X0Y0_FrameData[22]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5677_ (.I(Tile_X0Y0_FrameData[23]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5678_ (.I(Tile_X0Y0_FrameData[24]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5679_ (.I(Tile_X0Y0_FrameData[25]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5680_ (.I(Tile_X0Y0_FrameData[26]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5681_ (.I(Tile_X0Y0_FrameData[27]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5682_ (.I(Tile_X0Y0_FrameData[28]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5683_ (.I(Tile_X0Y0_FrameData[29]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5684_ (.I(Tile_X0Y0_FrameData[30]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5685_ (.I(Tile_X0Y0_FrameData[31]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5686_ (.I(Tile_X0Y1_FrameStrobe[0]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5687_ (.I(Tile_X0Y1_FrameStrobe[1]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5688_ (.I(Tile_X0Y1_FrameStrobe[2]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5689_ (.I(Tile_X0Y1_FrameStrobe[3]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5690_ (.I(Tile_X0Y1_FrameStrobe[4]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5691_ (.I(Tile_X0Y1_FrameStrobe[5]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5692_ (.I(Tile_X0Y1_FrameStrobe[6]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5693_ (.I(Tile_X0Y1_FrameStrobe[7]),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5694_ (.I(Tile_X0Y1_FrameStrobe[8]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5695_ (.I(Tile_X0Y1_FrameStrobe[9]),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5696_ (.I(Tile_X0Y1_FrameStrobe[10]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5697_ (.I(Tile_X0Y1_FrameStrobe[11]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5698_ (.I(Tile_X0Y1_FrameStrobe[12]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5699_ (.I(Tile_X0Y1_FrameStrobe[13]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5700_ (.I(Tile_X0Y1_FrameStrobe[14]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5701_ (.I(Tile_X0Y1_FrameStrobe[15]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5702_ (.I(Tile_X0Y1_FrameStrobe[16]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5703_ (.I(Tile_X0Y1_FrameStrobe[17]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5704_ (.I(Tile_X0Y1_FrameStrobe[18]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5705_ (.I(Tile_X0Y1_FrameStrobe[19]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5706_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 ),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5707_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 ),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5708_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 ),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5709_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 ),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5710_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5711_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5712_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5713_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5714_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5715_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5716_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5717_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5718_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5719_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5720_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5721_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5722_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5723_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5724_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5725_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5726_ (.I(Tile_X0Y1_N4END[8]),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5727_ (.I(Tile_X0Y1_N4END[9]),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5728_ (.I(Tile_X0Y1_N4END[10]),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5729_ (.I(Tile_X0Y1_N4END[11]),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5730_ (.I(Tile_X0Y1_N4END[12]),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5731_ (.I(Tile_X0Y1_N4END[13]),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5732_ (.I(Tile_X0Y1_N4END[14]),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5733_ (.I(Tile_X0Y1_N4END[15]),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5734_ (.I(\Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A ),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5735_ (.I(\Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A ),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5736_ (.I(\Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A ),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5737_ (.I(\Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A ),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5738_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 ),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5739_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 ),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5740_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 ),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5741_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 ),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5742_ (.I(Tile_X0Y1_NN4END[8]),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5743_ (.I(Tile_X0Y1_NN4END[9]),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5744_ (.I(Tile_X0Y1_NN4END[10]),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5745_ (.I(Tile_X0Y1_NN4END[11]),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5746_ (.I(Tile_X0Y1_NN4END[12]),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5747_ (.I(Tile_X0Y1_NN4END[13]),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5748_ (.I(Tile_X0Y1_NN4END[14]),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5749_ (.I(Tile_X0Y1_NN4END[15]),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5750_ (.I(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A ),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5751_ (.I(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A ),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5752_ (.I(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A ),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5753_ (.I(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A ),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5754_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 ),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5755_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 ),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5756_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 ),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5757_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 ),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5758_ (.I(clknet_1_0__leaf_Tile_X0Y1_UserCLK),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5759_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 ),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5760_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 ),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5761_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 ),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5762_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 ),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5763_ (.I(Tile_X0Y0_W2END[0]),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5764_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5765_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5766_ (.I(Tile_X0Y0_W2END[3]),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5767_ (.I(Tile_X0Y0_W2END[4]),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5768_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5769_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5770_ (.I(Tile_X0Y0_W2END[7]),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5771_ (.I(Tile_X0Y0_W2MID[0]),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5772_ (.I(Tile_X0Y0_W2MID[1]),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5773_ (.I(Tile_X0Y0_W2MID[2]),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5774_ (.I(Tile_X0Y0_W2MID[3]),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5775_ (.I(Tile_X0Y0_W2MID[4]),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5776_ (.I(Tile_X0Y0_W2MID[5]),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5777_ (.I(Tile_X0Y0_W2MID[6]),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5778_ (.I(Tile_X0Y0_W2MID[7]),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5779_ (.I(Tile_X0Y0_W6END[2]),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5780_ (.I(Tile_X0Y0_W6END[3]),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5781_ (.I(Tile_X0Y0_W6END[4]),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5782_ (.I(Tile_X0Y0_W6END[5]),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5783_ (.I(Tile_X0Y0_W6END[6]),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5784_ (.I(Tile_X0Y0_W6END[7]),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5785_ (.I(Tile_X0Y0_W6END[8]),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5786_ (.I(Tile_X0Y0_W6END[9]),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5787_ (.I(Tile_X0Y0_W6END[10]),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5788_ (.I(Tile_X0Y0_W6END[11]),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5789_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 ),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5790_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 ),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5791_ (.I(Tile_X0Y0_WW4END[4]),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5792_ (.I(Tile_X0Y0_WW4END[5]),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5793_ (.I(Tile_X0Y0_WW4END[6]),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5794_ (.I(Tile_X0Y0_WW4END[7]),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5795_ (.I(Tile_X0Y0_WW4END[8]),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5796_ (.I(Tile_X0Y0_WW4END[9]),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5797_ (.I(Tile_X0Y0_WW4END[10]),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5798_ (.I(Tile_X0Y0_WW4END[11]),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5799_ (.I(Tile_X0Y0_WW4END[12]),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5800_ (.I(Tile_X0Y0_WW4END[13]),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5801_ (.I(Tile_X0Y0_WW4END[14]),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5802_ (.I(Tile_X0Y0_WW4END[15]),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5803_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 ),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5804_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 ),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5805_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 ),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5806_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 ),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5807_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 ),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5808_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 ),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5809_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 ),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5810_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 ),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5811_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5812_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5813_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5814_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5815_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5816_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5817_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5818_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 ),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5819_ (.I(Tile_X0Y1_E2MID[0]),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5820_ (.I(Tile_X0Y1_E2MID[1]),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5821_ (.I(Tile_X0Y1_E2MID[2]),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5822_ (.I(Tile_X0Y1_E2MID[3]),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5823_ (.I(Tile_X0Y1_E2MID[4]),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5824_ (.I(Tile_X0Y1_E2MID[5]),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5825_ (.I(Tile_X0Y1_E2MID[6]),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5826_ (.I(Tile_X0Y1_E2MID[7]),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5827_ (.I(Tile_X0Y1_E6END[2]),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5828_ (.I(Tile_X0Y1_E6END[3]),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5829_ (.I(Tile_X0Y1_E6END[4]),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5830_ (.I(Tile_X0Y1_E6END[5]),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5831_ (.I(Tile_X0Y1_E6END[6]),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5832_ (.I(Tile_X0Y1_E6END[7]),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5833_ (.I(Tile_X0Y1_E6END[8]),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5834_ (.I(Tile_X0Y1_E6END[9]),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5835_ (.I(Tile_X0Y1_E6END[10]),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5836_ (.I(Tile_X0Y1_E6END[11]),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5837_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 ),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5838_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 ),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5839_ (.I(Tile_X0Y1_EE4END[4]),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5840_ (.I(Tile_X0Y1_EE4END[5]),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5841_ (.I(Tile_X0Y1_EE4END[6]),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5842_ (.I(Tile_X0Y1_EE4END[7]),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5843_ (.I(Tile_X0Y1_EE4END[8]),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5844_ (.I(Tile_X0Y1_EE4END[9]),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5845_ (.I(Tile_X0Y1_EE4END[10]),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5846_ (.I(Tile_X0Y1_EE4END[11]),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5847_ (.I(Tile_X0Y1_EE4END[12]),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5848_ (.I(Tile_X0Y1_EE4END[13]),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5849_ (.I(Tile_X0Y1_EE4END[14]),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5850_ (.I(Tile_X0Y1_EE4END[15]),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5851_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 ),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5852_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 ),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5853_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 ),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5854_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 ),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5855_ (.I(Tile_X0Y1_FrameData[0]),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5856_ (.I(Tile_X0Y1_FrameData[1]),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5857_ (.I(Tile_X0Y1_FrameData[2]),
    .Z(net272));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5858_ (.I(Tile_X0Y1_FrameData[3]),
    .Z(net275));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5859_ (.I(Tile_X0Y1_FrameData[4]),
    .Z(net276));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5860_ (.I(Tile_X0Y1_FrameData[5]),
    .Z(net277));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5861_ (.I(Tile_X0Y1_FrameData[6]),
    .Z(net278));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5862_ (.I(Tile_X0Y1_FrameData[7]),
    .Z(net279));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5863_ (.I(Tile_X0Y1_FrameData[8]),
    .Z(net280));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5864_ (.I(Tile_X0Y1_FrameData[9]),
    .Z(net281));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5865_ (.I(Tile_X0Y1_FrameData[10]),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5866_ (.I(Tile_X0Y1_FrameData[11]),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5867_ (.I(Tile_X0Y1_FrameData[12]),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5868_ (.I(Tile_X0Y1_FrameData[13]),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5869_ (.I(Tile_X0Y1_FrameData[14]),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5870_ (.I(Tile_X0Y1_FrameData[15]),
    .Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5871_ (.I(Tile_X0Y1_FrameData[16]),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5872_ (.I(Tile_X0Y1_FrameData[17]),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5873_ (.I(Tile_X0Y1_FrameData[18]),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5874_ (.I(Tile_X0Y1_FrameData[19]),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5875_ (.I(Tile_X0Y1_FrameData[20]),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5876_ (.I(Tile_X0Y1_FrameData[21]),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5877_ (.I(Tile_X0Y1_FrameData[22]),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5878_ (.I(Tile_X0Y1_FrameData[23]),
    .Z(net265));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5879_ (.I(Tile_X0Y1_FrameData[24]),
    .Z(net266));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5880_ (.I(Tile_X0Y1_FrameData[25]),
    .Z(net267));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5881_ (.I(Tile_X0Y1_FrameData[26]),
    .Z(net268));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5882_ (.I(Tile_X0Y1_FrameData[27]),
    .Z(net269));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5883_ (.I(Tile_X0Y1_FrameData[28]),
    .Z(net270));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5884_ (.I(Tile_X0Y1_FrameData[29]),
    .Z(net271));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5885_ (.I(Tile_X0Y1_FrameData[30]),
    .Z(net273));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5886_ (.I(Tile_X0Y1_FrameData[31]),
    .Z(net274));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5887_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 ),
    .Z(net282));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5888_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 ),
    .Z(net283));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5889_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 ),
    .Z(net284));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5890_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 ),
    .Z(net285));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5891_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ),
    .Z(net286));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5892_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ),
    .Z(net287));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5893_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .Z(net288));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5894_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .Z(net289));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5895_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ),
    .Z(net290));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5896_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ),
    .Z(net291));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5897_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ),
    .Z(net292));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5898_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ),
    .Z(net293));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5899_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .Z(net294));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5900_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5901_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .Z(net296));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5902_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .Z(net297));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5903_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .Z(net298));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5904_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .Z(net299));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5905_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .Z(net300));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5906_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .Z(net301));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5907_ (.I(Tile_X0Y0_S4END[8]),
    .Z(net302));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5908_ (.I(Tile_X0Y0_S4END[9]),
    .Z(net309));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5909_ (.I(Tile_X0Y0_S4END[10]),
    .Z(net310));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5910_ (.I(Tile_X0Y0_S4END[11]),
    .Z(net311));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5911_ (.I(Tile_X0Y0_S4END[12]),
    .Z(net312));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5912_ (.I(Tile_X0Y0_S4END[13]),
    .Z(net313));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5913_ (.I(Tile_X0Y0_S4END[14]),
    .Z(net314));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5914_ (.I(Tile_X0Y0_S4END[15]),
    .Z(net315));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5915_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 ),
    .Z(net316));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5916_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 ),
    .Z(net317));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5917_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 ),
    .Z(net303));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5918_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 ),
    .Z(net304));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5919_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 ),
    .Z(net305));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5920_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 ),
    .Z(net306));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5921_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 ),
    .Z(net307));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5922_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 ),
    .Z(net308));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5923_ (.I(Tile_X0Y0_SS4END[8]),
    .Z(net318));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5924_ (.I(Tile_X0Y0_SS4END[9]),
    .Z(net325));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5925_ (.I(Tile_X0Y0_SS4END[10]),
    .Z(net326));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5926_ (.I(Tile_X0Y0_SS4END[11]),
    .Z(net327));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5927_ (.I(Tile_X0Y0_SS4END[12]),
    .Z(net328));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5928_ (.I(Tile_X0Y0_SS4END[13]),
    .Z(net329));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5929_ (.I(Tile_X0Y0_SS4END[14]),
    .Z(net330));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5930_ (.I(Tile_X0Y0_SS4END[15]),
    .Z(net331));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5931_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 ),
    .Z(net332));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5932_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 ),
    .Z(net333));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5933_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 ),
    .Z(net319));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5934_ (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 ),
    .Z(net320));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5935_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 ),
    .Z(net321));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5936_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 ),
    .Z(net322));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5937_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 ),
    .Z(net323));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5938_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 ),
    .Z(net324));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5939_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 ),
    .Z(net334));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5940_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 ),
    .Z(net335));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5941_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 ),
    .Z(net336));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5942_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 ),
    .Z(net337));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5943_ (.I(Tile_X0Y1_W2END[0]),
    .Z(net338));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5944_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ),
    .Z(net339));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5945_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ),
    .Z(net340));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5946_ (.I(Tile_X0Y1_W2END[3]),
    .Z(net341));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5947_ (.I(Tile_X0Y1_W2END[4]),
    .Z(net342));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5948_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .Z(net343));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5949_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 ),
    .Z(net344));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5950_ (.I(Tile_X0Y1_W2END[7]),
    .Z(net345));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5951_ (.I(Tile_X0Y1_W2MID[0]),
    .Z(net346));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5952_ (.I(Tile_X0Y1_W2MID[1]),
    .Z(net347));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5953_ (.I(Tile_X0Y1_W2MID[2]),
    .Z(net348));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5954_ (.I(Tile_X0Y1_W2MID[3]),
    .Z(net349));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5955_ (.I(Tile_X0Y1_W2MID[4]),
    .Z(net350));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5956_ (.I(Tile_X0Y1_W2MID[5]),
    .Z(net351));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5957_ (.I(Tile_X0Y1_W2MID[6]),
    .Z(net352));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5958_ (.I(Tile_X0Y1_W2MID[7]),
    .Z(net353));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5959_ (.I(Tile_X0Y1_W6END[2]),
    .Z(net354));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5960_ (.I(Tile_X0Y1_W6END[3]),
    .Z(net357));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5961_ (.I(Tile_X0Y1_W6END[4]),
    .Z(net358));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5962_ (.I(Tile_X0Y1_W6END[5]),
    .Z(net359));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5963_ (.I(Tile_X0Y1_W6END[6]),
    .Z(net360));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5964_ (.I(Tile_X0Y1_W6END[7]),
    .Z(net361));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5965_ (.I(Tile_X0Y1_W6END[8]),
    .Z(net362));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5966_ (.I(Tile_X0Y1_W6END[9]),
    .Z(net363));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5967_ (.I(Tile_X0Y1_W6END[10]),
    .Z(net364));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5968_ (.I(Tile_X0Y1_W6END[11]),
    .Z(net365));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5969_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 ),
    .Z(net355));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5970_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 ),
    .Z(net356));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5971_ (.I(Tile_X0Y1_WW4END[4]),
    .Z(net366));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5972_ (.I(Tile_X0Y1_WW4END[5]),
    .Z(net373));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5973_ (.I(Tile_X0Y1_WW4END[6]),
    .Z(net374));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5974_ (.I(Tile_X0Y1_WW4END[7]),
    .Z(net375));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5975_ (.I(Tile_X0Y1_WW4END[8]),
    .Z(net376));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5976_ (.I(Tile_X0Y1_WW4END[9]),
    .Z(net377));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5977_ (.I(Tile_X0Y1_WW4END[10]),
    .Z(net378));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5978_ (.I(Tile_X0Y1_WW4END[11]),
    .Z(net379));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5979_ (.I(Tile_X0Y1_WW4END[12]),
    .Z(net380));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5980_ (.I(Tile_X0Y1_WW4END[13]),
    .Z(net381));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5981_ (.I(Tile_X0Y1_WW4END[14]),
    .Z(net367));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5982_ (.I(Tile_X0Y1_WW4END[15]),
    .Z(net368));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5983_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 ),
    .Z(net369));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5984_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 ),
    .Z(net370));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5985_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 ),
    .Z(net371));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5986_ (.I(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 ),
    .Z(net372));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output1 (.I(net1),
    .Z(Tile_X0Y0_E1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output2 (.I(net2),
    .Z(Tile_X0Y0_E1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output3 (.I(net3),
    .Z(Tile_X0Y0_E1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output4 (.I(net4),
    .Z(Tile_X0Y0_E1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output5 (.I(net5),
    .Z(Tile_X0Y0_E2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output6 (.I(net6),
    .Z(Tile_X0Y0_E2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output7 (.I(net7),
    .Z(Tile_X0Y0_E2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output8 (.I(net8),
    .Z(Tile_X0Y0_E2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output9 (.I(net9),
    .Z(Tile_X0Y0_E2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output10 (.I(net10),
    .Z(Tile_X0Y0_E2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output11 (.I(net11),
    .Z(Tile_X0Y0_E2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output12 (.I(net12),
    .Z(Tile_X0Y0_E2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output13 (.I(net13),
    .Z(Tile_X0Y0_E2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output14 (.I(net14),
    .Z(Tile_X0Y0_E2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output15 (.I(net15),
    .Z(Tile_X0Y0_E2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output16 (.I(net16),
    .Z(Tile_X0Y0_E2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output17 (.I(net17),
    .Z(Tile_X0Y0_E2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output18 (.I(net18),
    .Z(Tile_X0Y0_E2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output19 (.I(net19),
    .Z(Tile_X0Y0_E2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output20 (.I(net20),
    .Z(Tile_X0Y0_E2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output21 (.I(net21),
    .Z(Tile_X0Y0_E6BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output22 (.I(net22),
    .Z(Tile_X0Y0_E6BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output23 (.I(net23),
    .Z(Tile_X0Y0_E6BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output24 (.I(net24),
    .Z(Tile_X0Y0_E6BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output25 (.I(net25),
    .Z(Tile_X0Y0_E6BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output26 (.I(net26),
    .Z(Tile_X0Y0_E6BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output27 (.I(net27),
    .Z(Tile_X0Y0_E6BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output28 (.I(net28),
    .Z(Tile_X0Y0_E6BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output29 (.I(net29),
    .Z(Tile_X0Y0_E6BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output30 (.I(net30),
    .Z(Tile_X0Y0_E6BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output31 (.I(net31),
    .Z(Tile_X0Y0_E6BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output32 (.I(net32),
    .Z(Tile_X0Y0_E6BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output33 (.I(net33),
    .Z(Tile_X0Y0_EE4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output34 (.I(net34),
    .Z(Tile_X0Y0_EE4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output35 (.I(net35),
    .Z(Tile_X0Y0_EE4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output36 (.I(net36),
    .Z(Tile_X0Y0_EE4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output37 (.I(net37),
    .Z(Tile_X0Y0_EE4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output38 (.I(net38),
    .Z(Tile_X0Y0_EE4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output39 (.I(net39),
    .Z(Tile_X0Y0_EE4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output40 (.I(net40),
    .Z(Tile_X0Y0_EE4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output41 (.I(net41),
    .Z(Tile_X0Y0_EE4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output42 (.I(net42),
    .Z(Tile_X0Y0_EE4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output43 (.I(net43),
    .Z(Tile_X0Y0_EE4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output44 (.I(net44),
    .Z(Tile_X0Y0_EE4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output45 (.I(net45),
    .Z(Tile_X0Y0_EE4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output46 (.I(net46),
    .Z(Tile_X0Y0_EE4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output47 (.I(net47),
    .Z(Tile_X0Y0_EE4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output48 (.I(net48),
    .Z(Tile_X0Y0_EE4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output49 (.I(net49),
    .Z(Tile_X0Y0_FrameData_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output50 (.I(net50),
    .Z(Tile_X0Y0_FrameData_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output51 (.I(net51),
    .Z(Tile_X0Y0_FrameData_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output52 (.I(net52),
    .Z(Tile_X0Y0_FrameData_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output53 (.I(net53),
    .Z(Tile_X0Y0_FrameData_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output54 (.I(net54),
    .Z(Tile_X0Y0_FrameData_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output55 (.I(net55),
    .Z(Tile_X0Y0_FrameData_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output56 (.I(net56),
    .Z(Tile_X0Y0_FrameData_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output57 (.I(net57),
    .Z(Tile_X0Y0_FrameData_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output58 (.I(net58),
    .Z(Tile_X0Y0_FrameData_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output59 (.I(net59),
    .Z(Tile_X0Y0_FrameData_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output60 (.I(net60),
    .Z(Tile_X0Y0_FrameData_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output61 (.I(net61),
    .Z(Tile_X0Y0_FrameData_O[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output62 (.I(net62),
    .Z(Tile_X0Y0_FrameData_O[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output63 (.I(net63),
    .Z(Tile_X0Y0_FrameData_O[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output64 (.I(net64),
    .Z(Tile_X0Y0_FrameData_O[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output65 (.I(net65),
    .Z(Tile_X0Y0_FrameData_O[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output66 (.I(net66),
    .Z(Tile_X0Y0_FrameData_O[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output67 (.I(net67),
    .Z(Tile_X0Y0_FrameData_O[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output68 (.I(net68),
    .Z(Tile_X0Y0_FrameData_O[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output69 (.I(net69),
    .Z(Tile_X0Y0_FrameData_O[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output70 (.I(net70),
    .Z(Tile_X0Y0_FrameData_O[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output71 (.I(net71),
    .Z(Tile_X0Y0_FrameData_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output72 (.I(net72),
    .Z(Tile_X0Y0_FrameData_O[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output73 (.I(net73),
    .Z(Tile_X0Y0_FrameData_O[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output74 (.I(net74),
    .Z(Tile_X0Y0_FrameData_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output75 (.I(net75),
    .Z(Tile_X0Y0_FrameData_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output76 (.I(net76),
    .Z(Tile_X0Y0_FrameData_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output77 (.I(net77),
    .Z(Tile_X0Y0_FrameData_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output78 (.I(net78),
    .Z(Tile_X0Y0_FrameData_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output79 (.I(net79),
    .Z(Tile_X0Y0_FrameData_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output80 (.I(net80),
    .Z(Tile_X0Y0_FrameData_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output81 (.I(net81),
    .Z(Tile_X0Y0_FrameStrobe_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output82 (.I(net82),
    .Z(Tile_X0Y0_FrameStrobe_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output83 (.I(net83),
    .Z(Tile_X0Y0_FrameStrobe_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output84 (.I(net84),
    .Z(Tile_X0Y0_FrameStrobe_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output85 (.I(net85),
    .Z(Tile_X0Y0_FrameStrobe_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output86 (.I(net86),
    .Z(Tile_X0Y0_FrameStrobe_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output87 (.I(net87),
    .Z(Tile_X0Y0_FrameStrobe_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output88 (.I(net88),
    .Z(Tile_X0Y0_FrameStrobe_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output89 (.I(net89),
    .Z(Tile_X0Y0_FrameStrobe_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output90 (.I(net90),
    .Z(Tile_X0Y0_FrameStrobe_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output91 (.I(net91),
    .Z(Tile_X0Y0_FrameStrobe_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output92 (.I(net92),
    .Z(Tile_X0Y0_FrameStrobe_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output93 (.I(net93),
    .Z(Tile_X0Y0_FrameStrobe_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output94 (.I(net94),
    .Z(Tile_X0Y0_FrameStrobe_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output95 (.I(net95),
    .Z(Tile_X0Y0_FrameStrobe_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output96 (.I(net96),
    .Z(Tile_X0Y0_FrameStrobe_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output97 (.I(net97),
    .Z(Tile_X0Y0_FrameStrobe_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output98 (.I(net98),
    .Z(Tile_X0Y0_FrameStrobe_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output99 (.I(net99),
    .Z(Tile_X0Y0_FrameStrobe_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output100 (.I(net100),
    .Z(Tile_X0Y0_FrameStrobe_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output101 (.I(net101),
    .Z(Tile_X0Y0_N1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output102 (.I(net102),
    .Z(Tile_X0Y0_N1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output103 (.I(net103),
    .Z(Tile_X0Y0_N1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output104 (.I(net104),
    .Z(Tile_X0Y0_N1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output105 (.I(net105),
    .Z(Tile_X0Y0_N2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output106 (.I(net106),
    .Z(Tile_X0Y0_N2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output107 (.I(net107),
    .Z(Tile_X0Y0_N2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output108 (.I(net108),
    .Z(Tile_X0Y0_N2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output109 (.I(net109),
    .Z(Tile_X0Y0_N2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output110 (.I(net110),
    .Z(Tile_X0Y0_N2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output111 (.I(net111),
    .Z(Tile_X0Y0_N2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output112 (.I(net112),
    .Z(Tile_X0Y0_N2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output113 (.I(net113),
    .Z(Tile_X0Y0_N2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output114 (.I(net114),
    .Z(Tile_X0Y0_N2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output115 (.I(net115),
    .Z(Tile_X0Y0_N2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output116 (.I(net116),
    .Z(Tile_X0Y0_N2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output117 (.I(net117),
    .Z(Tile_X0Y0_N2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output118 (.I(net118),
    .Z(Tile_X0Y0_N2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output119 (.I(net119),
    .Z(Tile_X0Y0_N2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output120 (.I(net120),
    .Z(Tile_X0Y0_N2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output121 (.I(net121),
    .Z(Tile_X0Y0_N4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output122 (.I(net122),
    .Z(Tile_X0Y0_N4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output123 (.I(net123),
    .Z(Tile_X0Y0_N4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output124 (.I(net124),
    .Z(Tile_X0Y0_N4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output125 (.I(net125),
    .Z(Tile_X0Y0_N4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output126 (.I(net126),
    .Z(Tile_X0Y0_N4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output127 (.I(net127),
    .Z(Tile_X0Y0_N4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output128 (.I(net128),
    .Z(Tile_X0Y0_N4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output129 (.I(net129),
    .Z(Tile_X0Y0_N4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output130 (.I(net130),
    .Z(Tile_X0Y0_N4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output131 (.I(net131),
    .Z(Tile_X0Y0_N4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output132 (.I(net132),
    .Z(Tile_X0Y0_N4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output133 (.I(net133),
    .Z(Tile_X0Y0_N4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output134 (.I(net134),
    .Z(Tile_X0Y0_N4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output135 (.I(net135),
    .Z(Tile_X0Y0_N4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output136 (.I(net136),
    .Z(Tile_X0Y0_N4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output137 (.I(net137),
    .Z(Tile_X0Y0_NN4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output138 (.I(net138),
    .Z(Tile_X0Y0_NN4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output139 (.I(net139),
    .Z(Tile_X0Y0_NN4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output140 (.I(net140),
    .Z(Tile_X0Y0_NN4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output141 (.I(net141),
    .Z(Tile_X0Y0_NN4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output142 (.I(net142),
    .Z(Tile_X0Y0_NN4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output143 (.I(net143),
    .Z(Tile_X0Y0_NN4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output144 (.I(net144),
    .Z(Tile_X0Y0_NN4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output145 (.I(net145),
    .Z(Tile_X0Y0_NN4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output146 (.I(net146),
    .Z(Tile_X0Y0_NN4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output147 (.I(net147),
    .Z(Tile_X0Y0_NN4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output148 (.I(net148),
    .Z(Tile_X0Y0_NN4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output149 (.I(net149),
    .Z(Tile_X0Y0_NN4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output150 (.I(net150),
    .Z(Tile_X0Y0_NN4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output151 (.I(net151),
    .Z(Tile_X0Y0_NN4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output152 (.I(net152),
    .Z(Tile_X0Y0_NN4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output153 (.I(net153),
    .Z(Tile_X0Y0_UserCLKo));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output154 (.I(net154),
    .Z(Tile_X0Y0_W1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output155 (.I(net155),
    .Z(Tile_X0Y0_W1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output156 (.I(net156),
    .Z(Tile_X0Y0_W1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output157 (.I(net157),
    .Z(Tile_X0Y0_W1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output158 (.I(net158),
    .Z(Tile_X0Y0_W2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output159 (.I(net159),
    .Z(Tile_X0Y0_W2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output160 (.I(net160),
    .Z(Tile_X0Y0_W2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output161 (.I(net161),
    .Z(Tile_X0Y0_W2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output162 (.I(net162),
    .Z(Tile_X0Y0_W2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output163 (.I(net163),
    .Z(Tile_X0Y0_W2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output164 (.I(net164),
    .Z(Tile_X0Y0_W2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output165 (.I(net165),
    .Z(Tile_X0Y0_W2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output166 (.I(net166),
    .Z(Tile_X0Y0_W2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output167 (.I(net167),
    .Z(Tile_X0Y0_W2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output168 (.I(net168),
    .Z(Tile_X0Y0_W2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output169 (.I(net169),
    .Z(Tile_X0Y0_W2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output170 (.I(net170),
    .Z(Tile_X0Y0_W2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output171 (.I(net171),
    .Z(Tile_X0Y0_W2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output172 (.I(net172),
    .Z(Tile_X0Y0_W2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output173 (.I(net173),
    .Z(Tile_X0Y0_W2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output174 (.I(net174),
    .Z(Tile_X0Y0_W6BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output175 (.I(net175),
    .Z(Tile_X0Y0_W6BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output176 (.I(net176),
    .Z(Tile_X0Y0_W6BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output177 (.I(net177),
    .Z(Tile_X0Y0_W6BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output178 (.I(net178),
    .Z(Tile_X0Y0_W6BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output179 (.I(net179),
    .Z(Tile_X0Y0_W6BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output180 (.I(net180),
    .Z(Tile_X0Y0_W6BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output181 (.I(net181),
    .Z(Tile_X0Y0_W6BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output182 (.I(net182),
    .Z(Tile_X0Y0_W6BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output183 (.I(net183),
    .Z(Tile_X0Y0_W6BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output184 (.I(net184),
    .Z(Tile_X0Y0_W6BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output185 (.I(net185),
    .Z(Tile_X0Y0_W6BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output186 (.I(net186),
    .Z(Tile_X0Y0_WW4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output187 (.I(net187),
    .Z(Tile_X0Y0_WW4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output188 (.I(net188),
    .Z(Tile_X0Y0_WW4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output189 (.I(net189),
    .Z(Tile_X0Y0_WW4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output190 (.I(net190),
    .Z(Tile_X0Y0_WW4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output191 (.I(net191),
    .Z(Tile_X0Y0_WW4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output192 (.I(net192),
    .Z(Tile_X0Y0_WW4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output193 (.I(net193),
    .Z(Tile_X0Y0_WW4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output194 (.I(net194),
    .Z(Tile_X0Y0_WW4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output195 (.I(net195),
    .Z(Tile_X0Y0_WW4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output196 (.I(net196),
    .Z(Tile_X0Y0_WW4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output197 (.I(net197),
    .Z(Tile_X0Y0_WW4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output198 (.I(net198),
    .Z(Tile_X0Y0_WW4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output199 (.I(net199),
    .Z(Tile_X0Y0_WW4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output200 (.I(net200),
    .Z(Tile_X0Y0_WW4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output201 (.I(net201),
    .Z(Tile_X0Y0_WW4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output202 (.I(net202),
    .Z(Tile_X0Y1_E1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output203 (.I(net203),
    .Z(Tile_X0Y1_E1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output204 (.I(net204),
    .Z(Tile_X0Y1_E1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output205 (.I(net205),
    .Z(Tile_X0Y1_E1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output206 (.I(net206),
    .Z(Tile_X0Y1_E2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output207 (.I(net207),
    .Z(Tile_X0Y1_E2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output208 (.I(net208),
    .Z(Tile_X0Y1_E2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output209 (.I(net209),
    .Z(Tile_X0Y1_E2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output210 (.I(net210),
    .Z(Tile_X0Y1_E2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output211 (.I(net211),
    .Z(Tile_X0Y1_E2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output212 (.I(net212),
    .Z(Tile_X0Y1_E2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output213 (.I(net213),
    .Z(Tile_X0Y1_E2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output214 (.I(net214),
    .Z(Tile_X0Y1_E2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output215 (.I(net215),
    .Z(Tile_X0Y1_E2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output216 (.I(net216),
    .Z(Tile_X0Y1_E2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output217 (.I(net217),
    .Z(Tile_X0Y1_E2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output218 (.I(net218),
    .Z(Tile_X0Y1_E2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output219 (.I(net219),
    .Z(Tile_X0Y1_E2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output220 (.I(net220),
    .Z(Tile_X0Y1_E2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output221 (.I(net221),
    .Z(Tile_X0Y1_E2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output222 (.I(net222),
    .Z(Tile_X0Y1_E6BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output223 (.I(net223),
    .Z(Tile_X0Y1_E6BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output224 (.I(net224),
    .Z(Tile_X0Y1_E6BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output225 (.I(net225),
    .Z(Tile_X0Y1_E6BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output226 (.I(net226),
    .Z(Tile_X0Y1_E6BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output227 (.I(net227),
    .Z(Tile_X0Y1_E6BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output228 (.I(net228),
    .Z(Tile_X0Y1_E6BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output229 (.I(net229),
    .Z(Tile_X0Y1_E6BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output230 (.I(net230),
    .Z(Tile_X0Y1_E6BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output231 (.I(net231),
    .Z(Tile_X0Y1_E6BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output232 (.I(net232),
    .Z(Tile_X0Y1_E6BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output233 (.I(net233),
    .Z(Tile_X0Y1_E6BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output234 (.I(net234),
    .Z(Tile_X0Y1_EE4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output235 (.I(net235),
    .Z(Tile_X0Y1_EE4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output236 (.I(net236),
    .Z(Tile_X0Y1_EE4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output237 (.I(net237),
    .Z(Tile_X0Y1_EE4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output238 (.I(net238),
    .Z(Tile_X0Y1_EE4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output239 (.I(net239),
    .Z(Tile_X0Y1_EE4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output240 (.I(net240),
    .Z(Tile_X0Y1_EE4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output241 (.I(net241),
    .Z(Tile_X0Y1_EE4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output242 (.I(net242),
    .Z(Tile_X0Y1_EE4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output243 (.I(net243),
    .Z(Tile_X0Y1_EE4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output244 (.I(net244),
    .Z(Tile_X0Y1_EE4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output245 (.I(net245),
    .Z(Tile_X0Y1_EE4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output246 (.I(net246),
    .Z(Tile_X0Y1_EE4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output247 (.I(net247),
    .Z(Tile_X0Y1_EE4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output248 (.I(net248),
    .Z(Tile_X0Y1_EE4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output249 (.I(net249),
    .Z(Tile_X0Y1_EE4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output250 (.I(net250),
    .Z(Tile_X0Y1_FrameData_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output251 (.I(net251),
    .Z(Tile_X0Y1_FrameData_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output252 (.I(net252),
    .Z(Tile_X0Y1_FrameData_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output253 (.I(net253),
    .Z(Tile_X0Y1_FrameData_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output254 (.I(net254),
    .Z(Tile_X0Y1_FrameData_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output255 (.I(net255),
    .Z(Tile_X0Y1_FrameData_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output256 (.I(net256),
    .Z(Tile_X0Y1_FrameData_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output257 (.I(net257),
    .Z(Tile_X0Y1_FrameData_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output258 (.I(net258),
    .Z(Tile_X0Y1_FrameData_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output259 (.I(net259),
    .Z(Tile_X0Y1_FrameData_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output260 (.I(net260),
    .Z(Tile_X0Y1_FrameData_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output261 (.I(net261),
    .Z(Tile_X0Y1_FrameData_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output262 (.I(net262),
    .Z(Tile_X0Y1_FrameData_O[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output263 (.I(net263),
    .Z(Tile_X0Y1_FrameData_O[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output264 (.I(net264),
    .Z(Tile_X0Y1_FrameData_O[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output265 (.I(net265),
    .Z(Tile_X0Y1_FrameData_O[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output266 (.I(net266),
    .Z(Tile_X0Y1_FrameData_O[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output267 (.I(net267),
    .Z(Tile_X0Y1_FrameData_O[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output268 (.I(net268),
    .Z(Tile_X0Y1_FrameData_O[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output269 (.I(net269),
    .Z(Tile_X0Y1_FrameData_O[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output270 (.I(net270),
    .Z(Tile_X0Y1_FrameData_O[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output271 (.I(net271),
    .Z(Tile_X0Y1_FrameData_O[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output272 (.I(net272),
    .Z(Tile_X0Y1_FrameData_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output273 (.I(net273),
    .Z(Tile_X0Y1_FrameData_O[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output274 (.I(net274),
    .Z(Tile_X0Y1_FrameData_O[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output275 (.I(net275),
    .Z(Tile_X0Y1_FrameData_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output276 (.I(net276),
    .Z(Tile_X0Y1_FrameData_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output277 (.I(net277),
    .Z(Tile_X0Y1_FrameData_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output278 (.I(net278),
    .Z(Tile_X0Y1_FrameData_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output279 (.I(net279),
    .Z(Tile_X0Y1_FrameData_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output280 (.I(net280),
    .Z(Tile_X0Y1_FrameData_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output281 (.I(net281),
    .Z(Tile_X0Y1_FrameData_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output282 (.I(net282),
    .Z(Tile_X0Y1_S1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output283 (.I(net283),
    .Z(Tile_X0Y1_S1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output284 (.I(net284),
    .Z(Tile_X0Y1_S1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output285 (.I(net285),
    .Z(Tile_X0Y1_S1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output286 (.I(net286),
    .Z(Tile_X0Y1_S2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output287 (.I(net287),
    .Z(Tile_X0Y1_S2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output288 (.I(net288),
    .Z(Tile_X0Y1_S2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output289 (.I(net289),
    .Z(Tile_X0Y1_S2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output290 (.I(net290),
    .Z(Tile_X0Y1_S2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output291 (.I(net291),
    .Z(Tile_X0Y1_S2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output292 (.I(net292),
    .Z(Tile_X0Y1_S2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output293 (.I(net293),
    .Z(Tile_X0Y1_S2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output294 (.I(net294),
    .Z(Tile_X0Y1_S2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output295 (.I(net295),
    .Z(Tile_X0Y1_S2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output296 (.I(net296),
    .Z(Tile_X0Y1_S2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output297 (.I(net297),
    .Z(Tile_X0Y1_S2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output298 (.I(net298),
    .Z(Tile_X0Y1_S2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output299 (.I(net299),
    .Z(Tile_X0Y1_S2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output300 (.I(net300),
    .Z(Tile_X0Y1_S2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output301 (.I(net301),
    .Z(Tile_X0Y1_S2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output302 (.I(net302),
    .Z(Tile_X0Y1_S4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output303 (.I(net303),
    .Z(Tile_X0Y1_S4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output304 (.I(net304),
    .Z(Tile_X0Y1_S4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output305 (.I(net305),
    .Z(Tile_X0Y1_S4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output306 (.I(net306),
    .Z(Tile_X0Y1_S4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output307 (.I(net307),
    .Z(Tile_X0Y1_S4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output308 (.I(net308),
    .Z(Tile_X0Y1_S4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output309 (.I(net309),
    .Z(Tile_X0Y1_S4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output310 (.I(net310),
    .Z(Tile_X0Y1_S4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output311 (.I(net311),
    .Z(Tile_X0Y1_S4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output312 (.I(net312),
    .Z(Tile_X0Y1_S4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output313 (.I(net313),
    .Z(Tile_X0Y1_S4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output314 (.I(net314),
    .Z(Tile_X0Y1_S4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output315 (.I(net315),
    .Z(Tile_X0Y1_S4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output316 (.I(net316),
    .Z(Tile_X0Y1_S4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output317 (.I(net317),
    .Z(Tile_X0Y1_S4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output318 (.I(net318),
    .Z(Tile_X0Y1_SS4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output319 (.I(net319),
    .Z(Tile_X0Y1_SS4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output320 (.I(net320),
    .Z(Tile_X0Y1_SS4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output321 (.I(net321),
    .Z(Tile_X0Y1_SS4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output322 (.I(net322),
    .Z(Tile_X0Y1_SS4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output323 (.I(net323),
    .Z(Tile_X0Y1_SS4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output324 (.I(net324),
    .Z(Tile_X0Y1_SS4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output325 (.I(net325),
    .Z(Tile_X0Y1_SS4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output326 (.I(net326),
    .Z(Tile_X0Y1_SS4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output327 (.I(net327),
    .Z(Tile_X0Y1_SS4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output328 (.I(net328),
    .Z(Tile_X0Y1_SS4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output329 (.I(net329),
    .Z(Tile_X0Y1_SS4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output330 (.I(net330),
    .Z(Tile_X0Y1_SS4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output331 (.I(net331),
    .Z(Tile_X0Y1_SS4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output332 (.I(net332),
    .Z(Tile_X0Y1_SS4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output333 (.I(net333),
    .Z(Tile_X0Y1_SS4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output334 (.I(net334),
    .Z(Tile_X0Y1_W1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output335 (.I(net335),
    .Z(Tile_X0Y1_W1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output336 (.I(net336),
    .Z(Tile_X0Y1_W1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output337 (.I(net337),
    .Z(Tile_X0Y1_W1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output338 (.I(net338),
    .Z(Tile_X0Y1_W2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output339 (.I(net339),
    .Z(Tile_X0Y1_W2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output340 (.I(net340),
    .Z(Tile_X0Y1_W2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output341 (.I(net341),
    .Z(Tile_X0Y1_W2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output342 (.I(net342),
    .Z(Tile_X0Y1_W2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output343 (.I(net343),
    .Z(Tile_X0Y1_W2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output344 (.I(net344),
    .Z(Tile_X0Y1_W2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output345 (.I(net345),
    .Z(Tile_X0Y1_W2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output346 (.I(net346),
    .Z(Tile_X0Y1_W2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output347 (.I(net347),
    .Z(Tile_X0Y1_W2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output348 (.I(net348),
    .Z(Tile_X0Y1_W2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output349 (.I(net349),
    .Z(Tile_X0Y1_W2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output350 (.I(net350),
    .Z(Tile_X0Y1_W2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output351 (.I(net351),
    .Z(Tile_X0Y1_W2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output352 (.I(net352),
    .Z(Tile_X0Y1_W2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output353 (.I(net353),
    .Z(Tile_X0Y1_W2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output354 (.I(net354),
    .Z(Tile_X0Y1_W6BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output355 (.I(net355),
    .Z(Tile_X0Y1_W6BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output356 (.I(net356),
    .Z(Tile_X0Y1_W6BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output357 (.I(net357),
    .Z(Tile_X0Y1_W6BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output358 (.I(net358),
    .Z(Tile_X0Y1_W6BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output359 (.I(net359),
    .Z(Tile_X0Y1_W6BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output360 (.I(net360),
    .Z(Tile_X0Y1_W6BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output361 (.I(net361),
    .Z(Tile_X0Y1_W6BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output362 (.I(net362),
    .Z(Tile_X0Y1_W6BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output363 (.I(net363),
    .Z(Tile_X0Y1_W6BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output364 (.I(net364),
    .Z(Tile_X0Y1_W6BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output365 (.I(net365),
    .Z(Tile_X0Y1_W6BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output366 (.I(net366),
    .Z(Tile_X0Y1_WW4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output367 (.I(net367),
    .Z(Tile_X0Y1_WW4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output368 (.I(net368),
    .Z(Tile_X0Y1_WW4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output369 (.I(net369),
    .Z(Tile_X0Y1_WW4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output370 (.I(net370),
    .Z(Tile_X0Y1_WW4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output371 (.I(net371),
    .Z(Tile_X0Y1_WW4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output372 (.I(net372),
    .Z(Tile_X0Y1_WW4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output373 (.I(net373),
    .Z(Tile_X0Y1_WW4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output374 (.I(net374),
    .Z(Tile_X0Y1_WW4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output375 (.I(net375),
    .Z(Tile_X0Y1_WW4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output376 (.I(net376),
    .Z(Tile_X0Y1_WW4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output377 (.I(net377),
    .Z(Tile_X0Y1_WW4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output378 (.I(net378),
    .Z(Tile_X0Y1_WW4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output379 (.I(net379),
    .Z(Tile_X0Y1_WW4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output380 (.I(net380),
    .Z(Tile_X0Y1_WW4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output381 (.I(net381),
    .Z(Tile_X0Y1_WW4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_regs_0_Tile_X0Y1_UserCLK (.I(Tile_X0Y1_UserCLK),
    .Z(Tile_X0Y1_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_Tile_X0Y1_UserCLK (.I(Tile_X0Y1_UserCLK),
    .Z(clknet_0_Tile_X0Y1_UserCLK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_Tile_X0Y1_UserCLK (.I(clknet_0_Tile_X0Y1_UserCLK),
    .Z(clknet_1_0__leaf_Tile_X0Y1_UserCLK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_Tile_X0Y1_UserCLK_regs (.I(Tile_X0Y1_UserCLK_regs),
    .Z(clknet_0_Tile_X0Y1_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_Tile_X0Y1_UserCLK_regs (.I(clknet_0_Tile_X0Y1_UserCLK_regs),
    .Z(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_Tile_X0Y1_UserCLK_regs (.I(clknet_0_Tile_X0Y1_UserCLK_regs),
    .Z(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_Tile_X0Y1_UserCLK_regs (.I(clknet_0_Tile_X0Y1_UserCLK_regs),
    .Z(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_Tile_X0Y1_UserCLK_regs (.I(clknet_0_Tile_X0Y1_UserCLK_regs),
    .Z(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload0 (.I(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(Tile_X0Y0_E6END[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(Tile_X0Y0_E6END[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_3 (.I(Tile_X0Y0_E6END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_4 (.I(Tile_X0Y0_EE4END[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_5 (.I(Tile_X0Y0_EE4END[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_6 (.I(Tile_X0Y0_EE4END[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_7 (.I(Tile_X0Y0_EE4END[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_8 (.I(Tile_X0Y0_EE4END[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_9 (.I(Tile_X0Y0_EE4END[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_10 (.I(Tile_X0Y0_EE4END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_11 (.I(Tile_X0Y0_EE4END[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_12 (.I(Tile_X0Y0_W1END[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_13 (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_14 (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_15 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_16 (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_17 (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_18 (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_19 (.I(Tile_X0Y1_E6END[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_20 (.I(Tile_X0Y1_E6END[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_21 (.I(Tile_X0Y1_E6END[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_22 (.I(Tile_X0Y1_E6END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_23 (.I(Tile_X0Y1_EE4END[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_24 (.I(Tile_X0Y1_EE4END[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_25 (.I(Tile_X0Y1_EE4END[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_26 (.I(Tile_X0Y1_EE4END[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_27 (.I(Tile_X0Y1_EE4END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_28 (.I(Tile_X0Y1_EE4END[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_29 (.I(Tile_X0Y1_FrameStrobe[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_30 (.I(Tile_X0Y1_FrameStrobe[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_31 (.I(Tile_X0Y1_FrameStrobe[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_32 (.I(Tile_X0Y1_FrameStrobe[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_33 (.I(Tile_X0Y1_FrameStrobe[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_34 (.I(Tile_X0Y1_FrameStrobe[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_35 (.I(Tile_X0Y1_FrameStrobe[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_36 (.I(Tile_X0Y1_FrameStrobe[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_37 (.I(Tile_X0Y1_FrameStrobe[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_38 (.I(Tile_X0Y1_FrameStrobe[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_39 (.I(Tile_X0Y1_FrameStrobe[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_40 (.I(Tile_X0Y1_FrameStrobe[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_41 (.I(Tile_X0Y1_FrameStrobe[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_42 (.I(Tile_X0Y1_FrameStrobe[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_43 (.I(Tile_X0Y1_N4END[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_44 (.I(Tile_X0Y1_N4END[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_45 (.I(Tile_X0Y1_N4END[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_46 (.I(Tile_X0Y1_N4END[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_47 (.I(Tile_X0Y1_N4END[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_48 (.I(Tile_X0Y1_N4END[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_49 (.I(Tile_X0Y1_N4END[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_50 (.I(Tile_X0Y1_N4END[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_51 (.I(Tile_X0Y1_N4END[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_52 (.I(Tile_X0Y1_N4END[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_53 (.I(Tile_X0Y1_N4END[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_54 (.I(Tile_X0Y1_N4END[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_55 (.I(Tile_X0Y1_N4END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_56 (.I(Tile_X0Y1_N4END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_57 (.I(Tile_X0Y1_N4END[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_58 (.I(Tile_X0Y1_N4END[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_59 (.I(Tile_X0Y1_NN4END[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_60 (.I(Tile_X0Y1_NN4END[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_61 (.I(Tile_X0Y1_NN4END[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_62 (.I(Tile_X0Y1_NN4END[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_63 (.I(Tile_X0Y1_NN4END[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_64 (.I(Tile_X0Y1_NN4END[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_65 (.I(Tile_X0Y1_NN4END[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_66 (.I(Tile_X0Y1_NN4END[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_67 (.I(Tile_X0Y1_NN4END[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_68 (.I(Tile_X0Y1_NN4END[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_69 (.I(Tile_X0Y1_NN4END[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_70 (.I(Tile_X0Y1_NN4END[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_71 (.I(Tile_X0Y1_NN4END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_72 (.I(Tile_X0Y1_NN4END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_73 (.I(Tile_X0Y1_NN4END[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_74 (.I(Tile_X0Y1_NN4END[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_75 (.I(Tile_X0Y1_W2MID[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_76 (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_77 (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_78 (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_79 (.I(Tile_X0Y0_E6END[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_80 (.I(Tile_X0Y0_E6END[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_81 (.I(Tile_X0Y0_E6END[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_82 (.I(Tile_X0Y0_EE4END[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_83 (.I(Tile_X0Y0_EE4END[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_84 (.I(Tile_X0Y0_EE4END[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_85 (.I(Tile_X0Y0_SS4END[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_86 (.I(Tile_X0Y0_SS4END[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_87 (.I(Tile_X0Y0_SS4END[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_88 (.I(Tile_X0Y0_W2END[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_89 (.I(net365));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_90 (.I(net366));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_91 (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_92 (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_93 (.I(Tile_X0Y0_EE4END[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_94 (.I(Tile_X0Y0_W2END[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_95 (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_96 (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_97 (.I(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_98 (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_99 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_100 (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_101 (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_102 (.I(Tile_X0Y1_E6END[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_103 (.I(Tile_X0Y1_E6END[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_104 (.I(Tile_X0Y1_N4END[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_105 (.I(Tile_X0Y1_N4END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_106 (.I(Tile_X0Y1_NN4END[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_107 (.I(net373));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_108 (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_109 (.I(net380));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_110 (.I(net381));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_450 ();
endmodule
