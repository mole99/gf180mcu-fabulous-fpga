VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO W_IO4
  CLASS BLOCK ;
  FOREIGN W_IO4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 142.800 BY 287.280 ;
  PIN A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.680 0.560 16.240 ;
    END
  END A_I_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 11.200 0.560 11.760 ;
    END
  END A_O_top
  PIN A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.160 0.560 20.720 ;
    END
  END A_T_top
  PIN A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 64.960 0.560 65.520 ;
    END
  END A_config_C_bit0
  PIN A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 69.440 0.560 70.000 ;
    END
  END A_config_C_bit1
  PIN A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 73.920 0.560 74.480 ;
    END
  END A_config_C_bit2
  PIN A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.400 0.560 78.960 ;
    END
  END A_config_C_bit3
  PIN B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 29.120 0.560 29.680 ;
    END
  END B_I_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 24.640 0.560 25.200 ;
    END
  END B_O_top
  PIN B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.600 0.560 34.160 ;
    END
  END B_T_top
  PIN B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 82.880 0.560 83.440 ;
    END
  END B_config_C_bit0
  PIN B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 0.560 87.920 ;
    END
  END B_config_C_bit1
  PIN B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 91.840 0.560 92.400 ;
    END
  END B_config_C_bit2
  PIN B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.320 0.560 96.880 ;
    END
  END B_config_C_bit3
  PIN C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.560 0.560 43.120 ;
    END
  END C_I_top
  PIN C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 38.080 0.560 38.640 ;
    END
  END C_O_top
  PIN C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.040 0.560 47.600 ;
    END
  END C_T_top
  PIN C_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 0.560 101.360 ;
    END
  END C_config_C_bit0
  PIN C_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 105.280 0.560 105.840 ;
    END
  END C_config_C_bit1
  PIN C_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 109.760 0.560 110.320 ;
    END
  END C_config_C_bit2
  PIN C_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 0.560 114.800 ;
    END
  END C_config_C_bit3
  PIN D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 56.000 0.560 56.560 ;
    END
  END D_I_top
  PIN D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 51.520 0.560 52.080 ;
    END
  END D_O_top
  PIN D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.480 0.560 61.040 ;
    END
  END D_T_top
  PIN D_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.720 0.560 119.280 ;
    END
  END D_config_C_bit0
  PIN D_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 123.200 0.560 123.760 ;
    END
  END D_config_C_bit1
  PIN D_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 0.560 128.240 ;
    END
  END D_config_C_bit2
  PIN D_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.160 0.560 132.720 ;
    END
  END D_config_C_bit3
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 108.640 142.800 109.200 ;
    END
  END E1BEG[0]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 110.880 142.800 111.440 ;
    END
  END E1BEG[1]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 113.120 142.800 113.680 ;
    END
  END E1BEG[2]
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 115.360 142.800 115.920 ;
    END
  END E1BEG[3]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 117.600 142.800 118.160 ;
    END
  END E2BEG[0]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 119.840 142.800 120.400 ;
    END
  END E2BEG[1]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 122.080 142.800 122.640 ;
    END
  END E2BEG[2]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 124.320 142.800 124.880 ;
    END
  END E2BEG[3]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 126.560 142.800 127.120 ;
    END
  END E2BEG[4]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 128.800 142.800 129.360 ;
    END
  END E2BEG[5]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 131.040 142.800 131.600 ;
    END
  END E2BEG[6]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 133.280 142.800 133.840 ;
    END
  END E2BEG[7]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 135.520 142.800 136.080 ;
    END
  END E2BEGb[0]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 137.760 142.800 138.320 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 140.000 142.800 140.560 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 142.240 142.800 142.800 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 144.480 142.800 145.040 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 146.720 142.800 147.280 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 148.960 142.800 149.520 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 151.200 142.800 151.760 ;
    END
  END E2BEGb[7]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 189.280 142.800 189.840 ;
    END
  END E6BEG[0]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 211.680 142.800 212.240 ;
    END
  END E6BEG[10]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 213.920 142.800 214.480 ;
    END
  END E6BEG[11]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 191.520 142.800 192.080 ;
    END
  END E6BEG[1]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 193.760 142.800 194.320 ;
    END
  END E6BEG[2]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 196.000 142.800 196.560 ;
    END
  END E6BEG[3]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 198.240 142.800 198.800 ;
    END
  END E6BEG[4]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 200.480 142.800 201.040 ;
    END
  END E6BEG[5]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 202.720 142.800 203.280 ;
    END
  END E6BEG[6]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 204.960 142.800 205.520 ;
    END
  END E6BEG[7]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 207.200 142.800 207.760 ;
    END
  END E6BEG[8]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 209.440 142.800 210.000 ;
    END
  END E6BEG[9]
  PIN EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 153.440 142.800 154.000 ;
    END
  END EE4BEG[0]
  PIN EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 175.840 142.800 176.400 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 178.080 142.800 178.640 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 180.320 142.800 180.880 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 182.560 142.800 183.120 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 184.800 142.800 185.360 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 187.040 142.800 187.600 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 155.680 142.800 156.240 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 157.920 142.800 158.480 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 160.160 142.800 160.720 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 162.400 142.800 162.960 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 164.640 142.800 165.200 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 166.880 142.800 167.440 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 169.120 142.800 169.680 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 171.360 142.800 171.920 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 173.600 142.800 174.160 ;
    END
  END EE4BEG[9]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 136.640 0.560 137.200 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 181.440 0.560 182.000 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 185.920 0.560 186.480 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 190.400 0.560 190.960 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.880 0.560 195.440 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 199.360 0.560 199.920 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 203.840 0.560 204.400 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 208.320 0.560 208.880 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 212.800 0.560 213.360 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 217.280 0.560 217.840 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.760 0.560 222.320 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 0.560 141.680 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 226.240 0.560 226.800 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.720 0.560 231.280 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 235.200 0.560 235.760 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 239.680 0.560 240.240 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 244.160 0.560 244.720 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 248.640 0.560 249.200 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 253.120 0.560 253.680 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 257.600 0.560 258.160 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.080 0.560 262.640 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 266.560 0.560 267.120 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 145.600 0.560 146.160 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 271.040 0.560 271.600 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 275.520 0.560 276.080 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.080 0.560 150.640 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 0.560 155.120 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 159.040 0.560 159.600 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 163.520 0.560 164.080 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 0.560 168.560 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 172.480 0.560 173.040 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 176.960 0.560 177.520 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 216.160 142.800 216.720 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 238.560 142.800 239.120 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 240.800 142.800 241.360 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 243.040 142.800 243.600 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 245.280 142.800 245.840 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 247.520 142.800 248.080 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 249.760 142.800 250.320 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 252.000 142.800 252.560 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 254.240 142.800 254.800 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 256.480 142.800 257.040 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 258.720 142.800 259.280 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 218.400 142.800 218.960 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 260.960 142.800 261.520 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 263.200 142.800 263.760 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 265.440 142.800 266.000 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 267.680 142.800 268.240 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 269.920 142.800 270.480 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 272.160 142.800 272.720 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 274.400 142.800 274.960 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 276.640 142.800 277.200 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 278.880 142.800 279.440 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 281.120 142.800 281.680 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 220.640 142.800 221.200 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 283.360 142.800 283.920 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 285.600 142.800 286.160 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 222.880 142.800 223.440 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 225.120 142.800 225.680 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 227.360 142.800 227.920 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 229.600 142.800 230.160 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 231.840 142.800 232.400 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 234.080 142.800 234.640 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 236.320 142.800 236.880 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 0.000 10.640 0.560 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 0.560 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 0.560 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 0.560 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 0.560 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 0.560 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 0.560 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 0.000 118.160 0.560 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 0.560 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 0.560 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 0.000 138.320 0.560 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 0.000 17.360 0.560 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 0.560 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.510000 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 0.560 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 0.560 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 0.560 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 0.560 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 0.000 57.680 0.560 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 0.560 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 0.560 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 286.720 10.640 287.280 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 286.720 77.840 287.280 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 286.720 84.560 287.280 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 286.720 91.280 287.280 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 286.720 98.000 287.280 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 286.720 104.720 287.280 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 286.720 111.440 287.280 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 286.720 118.160 287.280 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 286.720 124.880 287.280 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 286.720 131.600 287.280 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 286.720 138.320 287.280 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 286.720 17.360 287.280 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 286.720 24.080 287.280 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 286.720 30.800 287.280 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 286.720 37.520 287.280 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 286.720 44.240 287.280 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 286.720 50.960 287.280 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 286.720 57.680 287.280 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 286.720 64.400 287.280 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 286.720 71.120 287.280 ;
    END
  END FrameStrobe_O[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.476000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 0.560 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 286.720 3.920 287.280 ;
    END
  END UserCLKo
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.880 0.000 20.480 287.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 118.880 0.000 120.480 287.280 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.180 0.000 23.780 287.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.180 0.000 123.780 287.280 ;
    END
  END VSS
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 1.120 142.800 1.680 ;
    END
  END W1END[0]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 3.360 142.800 3.920 ;
    END
  END W1END[1]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 5.600 142.800 6.160 ;
    END
  END W1END[2]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 7.840 142.800 8.400 ;
    END
  END W1END[3]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 28.000 142.800 28.560 ;
    END
  END W2END[0]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 30.240 142.800 30.800 ;
    END
  END W2END[1]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 32.480 142.800 33.040 ;
    END
  END W2END[2]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 34.720 142.800 35.280 ;
    END
  END W2END[3]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 36.960 142.800 37.520 ;
    END
  END W2END[4]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 39.200 142.800 39.760 ;
    END
  END W2END[5]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 41.440 142.800 42.000 ;
    END
  END W2END[6]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 43.680 142.800 44.240 ;
    END
  END W2END[7]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 10.080 142.800 10.640 ;
    END
  END W2MID[0]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 12.320 142.800 12.880 ;
    END
  END W2MID[1]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 14.560 142.800 15.120 ;
    END
  END W2MID[2]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 16.800 142.800 17.360 ;
    END
  END W2MID[3]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 19.040 142.800 19.600 ;
    END
  END W2MID[4]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 21.280 142.800 21.840 ;
    END
  END W2MID[5]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 23.520 142.800 24.080 ;
    END
  END W2MID[6]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 25.760 142.800 26.320 ;
    END
  END W2MID[7]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 81.760 142.800 82.320 ;
    END
  END W6END[0]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 104.160 142.800 104.720 ;
    END
  END W6END[10]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 106.400 142.800 106.960 ;
    END
  END W6END[11]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 84.000 142.800 84.560 ;
    END
  END W6END[1]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 86.240 142.800 86.800 ;
    END
  END W6END[2]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 88.480 142.800 89.040 ;
    END
  END W6END[3]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 90.720 142.800 91.280 ;
    END
  END W6END[4]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 92.960 142.800 93.520 ;
    END
  END W6END[5]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 95.200 142.800 95.760 ;
    END
  END W6END[6]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 97.440 142.800 98.000 ;
    END
  END W6END[7]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 99.680 142.800 100.240 ;
    END
  END W6END[8]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 101.920 142.800 102.480 ;
    END
  END W6END[9]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 45.920 142.800 46.480 ;
    END
  END WW4END[0]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 68.320 142.800 68.880 ;
    END
  END WW4END[10]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 70.560 142.800 71.120 ;
    END
  END WW4END[11]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 72.800 142.800 73.360 ;
    END
  END WW4END[12]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 75.040 142.800 75.600 ;
    END
  END WW4END[13]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 77.280 142.800 77.840 ;
    END
  END WW4END[14]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 79.520 142.800 80.080 ;
    END
  END WW4END[15]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 48.160 142.800 48.720 ;
    END
  END WW4END[1]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 50.400 142.800 50.960 ;
    END
  END WW4END[2]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 52.640 142.800 53.200 ;
    END
  END WW4END[3]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 54.880 142.800 55.440 ;
    END
  END WW4END[4]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 57.120 142.800 57.680 ;
    END
  END WW4END[5]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 59.360 142.800 59.920 ;
    END
  END WW4END[6]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 61.600 142.800 62.160 ;
    END
  END WW4END[7]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 63.840 142.800 64.400 ;
    END
  END WW4END[8]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 142.240 66.080 142.800 66.640 ;
    END
  END WW4END[9]
  OBS
      LAYER Nwell ;
        RECT 2.930 3.490 139.870 282.670 ;
      LAYER Metal1 ;
        RECT 3.360 3.620 139.440 282.540 ;
      LAYER Metal2 ;
        RECT 0.140 286.420 3.060 287.140 ;
        RECT 4.220 286.420 9.780 287.140 ;
        RECT 10.940 286.420 16.500 287.140 ;
        RECT 17.660 286.420 23.220 287.140 ;
        RECT 24.380 286.420 29.940 287.140 ;
        RECT 31.100 286.420 36.660 287.140 ;
        RECT 37.820 286.420 43.380 287.140 ;
        RECT 44.540 286.420 50.100 287.140 ;
        RECT 51.260 286.420 56.820 287.140 ;
        RECT 57.980 286.420 63.540 287.140 ;
        RECT 64.700 286.420 70.260 287.140 ;
        RECT 71.420 286.420 76.980 287.140 ;
        RECT 78.140 286.420 83.700 287.140 ;
        RECT 84.860 286.420 90.420 287.140 ;
        RECT 91.580 286.420 97.140 287.140 ;
        RECT 98.300 286.420 103.860 287.140 ;
        RECT 105.020 286.420 110.580 287.140 ;
        RECT 111.740 286.420 117.300 287.140 ;
        RECT 118.460 286.420 124.020 287.140 ;
        RECT 125.180 286.420 130.740 287.140 ;
        RECT 131.900 286.420 137.460 287.140 ;
        RECT 138.620 286.420 141.540 287.140 ;
        RECT 0.140 0.860 141.540 286.420 ;
        RECT 0.140 0.560 3.060 0.860 ;
        RECT 4.220 0.560 9.780 0.860 ;
        RECT 10.940 0.560 16.500 0.860 ;
        RECT 17.660 0.560 23.220 0.860 ;
        RECT 24.380 0.560 29.940 0.860 ;
        RECT 31.100 0.560 36.660 0.860 ;
        RECT 37.820 0.560 43.380 0.860 ;
        RECT 44.540 0.560 50.100 0.860 ;
        RECT 51.260 0.560 56.820 0.860 ;
        RECT 57.980 0.560 63.540 0.860 ;
        RECT 64.700 0.560 70.260 0.860 ;
        RECT 71.420 0.560 76.980 0.860 ;
        RECT 78.140 0.560 83.700 0.860 ;
        RECT 84.860 0.560 90.420 0.860 ;
        RECT 91.580 0.560 97.140 0.860 ;
        RECT 98.300 0.560 103.860 0.860 ;
        RECT 105.020 0.560 110.580 0.860 ;
        RECT 111.740 0.560 117.300 0.860 ;
        RECT 118.460 0.560 124.020 0.860 ;
        RECT 125.180 0.560 130.740 0.860 ;
        RECT 131.900 0.560 137.460 0.860 ;
        RECT 138.620 0.560 141.540 0.860 ;
      LAYER Metal3 ;
        RECT 0.560 286.460 142.240 286.580 ;
        RECT 0.560 285.300 141.940 286.460 ;
        RECT 0.560 284.220 142.240 285.300 ;
        RECT 0.560 283.060 141.940 284.220 ;
        RECT 0.560 281.980 142.240 283.060 ;
        RECT 0.560 280.820 141.940 281.980 ;
        RECT 0.560 279.740 142.240 280.820 ;
        RECT 0.560 278.580 141.940 279.740 ;
        RECT 0.560 277.500 142.240 278.580 ;
        RECT 0.560 276.380 141.940 277.500 ;
        RECT 0.860 276.340 141.940 276.380 ;
        RECT 0.860 275.260 142.240 276.340 ;
        RECT 0.860 275.220 141.940 275.260 ;
        RECT 0.560 274.100 141.940 275.220 ;
        RECT 0.560 273.020 142.240 274.100 ;
        RECT 0.560 271.900 141.940 273.020 ;
        RECT 0.860 271.860 141.940 271.900 ;
        RECT 0.860 270.780 142.240 271.860 ;
        RECT 0.860 270.740 141.940 270.780 ;
        RECT 0.560 269.620 141.940 270.740 ;
        RECT 0.560 268.540 142.240 269.620 ;
        RECT 0.560 267.420 141.940 268.540 ;
        RECT 0.860 267.380 141.940 267.420 ;
        RECT 0.860 266.300 142.240 267.380 ;
        RECT 0.860 266.260 141.940 266.300 ;
        RECT 0.560 265.140 141.940 266.260 ;
        RECT 0.560 264.060 142.240 265.140 ;
        RECT 0.560 262.940 141.940 264.060 ;
        RECT 0.860 262.900 141.940 262.940 ;
        RECT 0.860 261.820 142.240 262.900 ;
        RECT 0.860 261.780 141.940 261.820 ;
        RECT 0.560 260.660 141.940 261.780 ;
        RECT 0.560 259.580 142.240 260.660 ;
        RECT 0.560 258.460 141.940 259.580 ;
        RECT 0.860 258.420 141.940 258.460 ;
        RECT 0.860 257.340 142.240 258.420 ;
        RECT 0.860 257.300 141.940 257.340 ;
        RECT 0.560 256.180 141.940 257.300 ;
        RECT 0.560 255.100 142.240 256.180 ;
        RECT 0.560 253.980 141.940 255.100 ;
        RECT 0.860 253.940 141.940 253.980 ;
        RECT 0.860 252.860 142.240 253.940 ;
        RECT 0.860 252.820 141.940 252.860 ;
        RECT 0.560 251.700 141.940 252.820 ;
        RECT 0.560 250.620 142.240 251.700 ;
        RECT 0.560 249.500 141.940 250.620 ;
        RECT 0.860 249.460 141.940 249.500 ;
        RECT 0.860 248.380 142.240 249.460 ;
        RECT 0.860 248.340 141.940 248.380 ;
        RECT 0.560 247.220 141.940 248.340 ;
        RECT 0.560 246.140 142.240 247.220 ;
        RECT 0.560 245.020 141.940 246.140 ;
        RECT 0.860 244.980 141.940 245.020 ;
        RECT 0.860 243.900 142.240 244.980 ;
        RECT 0.860 243.860 141.940 243.900 ;
        RECT 0.560 242.740 141.940 243.860 ;
        RECT 0.560 241.660 142.240 242.740 ;
        RECT 0.560 240.540 141.940 241.660 ;
        RECT 0.860 240.500 141.940 240.540 ;
        RECT 0.860 239.420 142.240 240.500 ;
        RECT 0.860 239.380 141.940 239.420 ;
        RECT 0.560 238.260 141.940 239.380 ;
        RECT 0.560 237.180 142.240 238.260 ;
        RECT 0.560 236.060 141.940 237.180 ;
        RECT 0.860 236.020 141.940 236.060 ;
        RECT 0.860 234.940 142.240 236.020 ;
        RECT 0.860 234.900 141.940 234.940 ;
        RECT 0.560 233.780 141.940 234.900 ;
        RECT 0.560 232.700 142.240 233.780 ;
        RECT 0.560 231.580 141.940 232.700 ;
        RECT 0.860 231.540 141.940 231.580 ;
        RECT 0.860 230.460 142.240 231.540 ;
        RECT 0.860 230.420 141.940 230.460 ;
        RECT 0.560 229.300 141.940 230.420 ;
        RECT 0.560 228.220 142.240 229.300 ;
        RECT 0.560 227.100 141.940 228.220 ;
        RECT 0.860 227.060 141.940 227.100 ;
        RECT 0.860 225.980 142.240 227.060 ;
        RECT 0.860 225.940 141.940 225.980 ;
        RECT 0.560 224.820 141.940 225.940 ;
        RECT 0.560 223.740 142.240 224.820 ;
        RECT 0.560 222.620 141.940 223.740 ;
        RECT 0.860 222.580 141.940 222.620 ;
        RECT 0.860 221.500 142.240 222.580 ;
        RECT 0.860 221.460 141.940 221.500 ;
        RECT 0.560 220.340 141.940 221.460 ;
        RECT 0.560 219.260 142.240 220.340 ;
        RECT 0.560 218.140 141.940 219.260 ;
        RECT 0.860 218.100 141.940 218.140 ;
        RECT 0.860 217.020 142.240 218.100 ;
        RECT 0.860 216.980 141.940 217.020 ;
        RECT 0.560 215.860 141.940 216.980 ;
        RECT 0.560 214.780 142.240 215.860 ;
        RECT 0.560 213.660 141.940 214.780 ;
        RECT 0.860 213.620 141.940 213.660 ;
        RECT 0.860 212.540 142.240 213.620 ;
        RECT 0.860 212.500 141.940 212.540 ;
        RECT 0.560 211.380 141.940 212.500 ;
        RECT 0.560 210.300 142.240 211.380 ;
        RECT 0.560 209.180 141.940 210.300 ;
        RECT 0.860 209.140 141.940 209.180 ;
        RECT 0.860 208.060 142.240 209.140 ;
        RECT 0.860 208.020 141.940 208.060 ;
        RECT 0.560 206.900 141.940 208.020 ;
        RECT 0.560 205.820 142.240 206.900 ;
        RECT 0.560 204.700 141.940 205.820 ;
        RECT 0.860 204.660 141.940 204.700 ;
        RECT 0.860 203.580 142.240 204.660 ;
        RECT 0.860 203.540 141.940 203.580 ;
        RECT 0.560 202.420 141.940 203.540 ;
        RECT 0.560 201.340 142.240 202.420 ;
        RECT 0.560 200.220 141.940 201.340 ;
        RECT 0.860 200.180 141.940 200.220 ;
        RECT 0.860 199.100 142.240 200.180 ;
        RECT 0.860 199.060 141.940 199.100 ;
        RECT 0.560 197.940 141.940 199.060 ;
        RECT 0.560 196.860 142.240 197.940 ;
        RECT 0.560 195.740 141.940 196.860 ;
        RECT 0.860 195.700 141.940 195.740 ;
        RECT 0.860 194.620 142.240 195.700 ;
        RECT 0.860 194.580 141.940 194.620 ;
        RECT 0.560 193.460 141.940 194.580 ;
        RECT 0.560 192.380 142.240 193.460 ;
        RECT 0.560 191.260 141.940 192.380 ;
        RECT 0.860 191.220 141.940 191.260 ;
        RECT 0.860 190.140 142.240 191.220 ;
        RECT 0.860 190.100 141.940 190.140 ;
        RECT 0.560 188.980 141.940 190.100 ;
        RECT 0.560 187.900 142.240 188.980 ;
        RECT 0.560 186.780 141.940 187.900 ;
        RECT 0.860 186.740 141.940 186.780 ;
        RECT 0.860 185.660 142.240 186.740 ;
        RECT 0.860 185.620 141.940 185.660 ;
        RECT 0.560 184.500 141.940 185.620 ;
        RECT 0.560 183.420 142.240 184.500 ;
        RECT 0.560 182.300 141.940 183.420 ;
        RECT 0.860 182.260 141.940 182.300 ;
        RECT 0.860 181.180 142.240 182.260 ;
        RECT 0.860 181.140 141.940 181.180 ;
        RECT 0.560 180.020 141.940 181.140 ;
        RECT 0.560 178.940 142.240 180.020 ;
        RECT 0.560 177.820 141.940 178.940 ;
        RECT 0.860 177.780 141.940 177.820 ;
        RECT 0.860 176.700 142.240 177.780 ;
        RECT 0.860 176.660 141.940 176.700 ;
        RECT 0.560 175.540 141.940 176.660 ;
        RECT 0.560 174.460 142.240 175.540 ;
        RECT 0.560 173.340 141.940 174.460 ;
        RECT 0.860 173.300 141.940 173.340 ;
        RECT 0.860 172.220 142.240 173.300 ;
        RECT 0.860 172.180 141.940 172.220 ;
        RECT 0.560 171.060 141.940 172.180 ;
        RECT 0.560 169.980 142.240 171.060 ;
        RECT 0.560 168.860 141.940 169.980 ;
        RECT 0.860 168.820 141.940 168.860 ;
        RECT 0.860 167.740 142.240 168.820 ;
        RECT 0.860 167.700 141.940 167.740 ;
        RECT 0.560 166.580 141.940 167.700 ;
        RECT 0.560 165.500 142.240 166.580 ;
        RECT 0.560 164.380 141.940 165.500 ;
        RECT 0.860 164.340 141.940 164.380 ;
        RECT 0.860 163.260 142.240 164.340 ;
        RECT 0.860 163.220 141.940 163.260 ;
        RECT 0.560 162.100 141.940 163.220 ;
        RECT 0.560 161.020 142.240 162.100 ;
        RECT 0.560 159.900 141.940 161.020 ;
        RECT 0.860 159.860 141.940 159.900 ;
        RECT 0.860 158.780 142.240 159.860 ;
        RECT 0.860 158.740 141.940 158.780 ;
        RECT 0.560 157.620 141.940 158.740 ;
        RECT 0.560 156.540 142.240 157.620 ;
        RECT 0.560 155.420 141.940 156.540 ;
        RECT 0.860 155.380 141.940 155.420 ;
        RECT 0.860 154.300 142.240 155.380 ;
        RECT 0.860 154.260 141.940 154.300 ;
        RECT 0.560 153.140 141.940 154.260 ;
        RECT 0.560 152.060 142.240 153.140 ;
        RECT 0.560 150.940 141.940 152.060 ;
        RECT 0.860 150.900 141.940 150.940 ;
        RECT 0.860 149.820 142.240 150.900 ;
        RECT 0.860 149.780 141.940 149.820 ;
        RECT 0.560 148.660 141.940 149.780 ;
        RECT 0.560 147.580 142.240 148.660 ;
        RECT 0.560 146.460 141.940 147.580 ;
        RECT 0.860 146.420 141.940 146.460 ;
        RECT 0.860 145.340 142.240 146.420 ;
        RECT 0.860 145.300 141.940 145.340 ;
        RECT 0.560 144.180 141.940 145.300 ;
        RECT 0.560 143.100 142.240 144.180 ;
        RECT 0.560 141.980 141.940 143.100 ;
        RECT 0.860 141.940 141.940 141.980 ;
        RECT 0.860 140.860 142.240 141.940 ;
        RECT 0.860 140.820 141.940 140.860 ;
        RECT 0.560 139.700 141.940 140.820 ;
        RECT 0.560 138.620 142.240 139.700 ;
        RECT 0.560 137.500 141.940 138.620 ;
        RECT 0.860 137.460 141.940 137.500 ;
        RECT 0.860 136.380 142.240 137.460 ;
        RECT 0.860 136.340 141.940 136.380 ;
        RECT 0.560 135.220 141.940 136.340 ;
        RECT 0.560 134.140 142.240 135.220 ;
        RECT 0.560 133.020 141.940 134.140 ;
        RECT 0.860 132.980 141.940 133.020 ;
        RECT 0.860 131.900 142.240 132.980 ;
        RECT 0.860 131.860 141.940 131.900 ;
        RECT 0.560 130.740 141.940 131.860 ;
        RECT 0.560 129.660 142.240 130.740 ;
        RECT 0.560 128.540 141.940 129.660 ;
        RECT 0.860 128.500 141.940 128.540 ;
        RECT 0.860 127.420 142.240 128.500 ;
        RECT 0.860 127.380 141.940 127.420 ;
        RECT 0.560 126.260 141.940 127.380 ;
        RECT 0.560 125.180 142.240 126.260 ;
        RECT 0.560 124.060 141.940 125.180 ;
        RECT 0.860 124.020 141.940 124.060 ;
        RECT 0.860 122.940 142.240 124.020 ;
        RECT 0.860 122.900 141.940 122.940 ;
        RECT 0.560 121.780 141.940 122.900 ;
        RECT 0.560 120.700 142.240 121.780 ;
        RECT 0.560 119.580 141.940 120.700 ;
        RECT 0.860 119.540 141.940 119.580 ;
        RECT 0.860 118.460 142.240 119.540 ;
        RECT 0.860 118.420 141.940 118.460 ;
        RECT 0.560 117.300 141.940 118.420 ;
        RECT 0.560 116.220 142.240 117.300 ;
        RECT 0.560 115.100 141.940 116.220 ;
        RECT 0.860 115.060 141.940 115.100 ;
        RECT 0.860 113.980 142.240 115.060 ;
        RECT 0.860 113.940 141.940 113.980 ;
        RECT 0.560 112.820 141.940 113.940 ;
        RECT 0.560 111.740 142.240 112.820 ;
        RECT 0.560 110.620 141.940 111.740 ;
        RECT 0.860 110.580 141.940 110.620 ;
        RECT 0.860 109.500 142.240 110.580 ;
        RECT 0.860 109.460 141.940 109.500 ;
        RECT 0.560 108.340 141.940 109.460 ;
        RECT 0.560 107.260 142.240 108.340 ;
        RECT 0.560 106.140 141.940 107.260 ;
        RECT 0.860 106.100 141.940 106.140 ;
        RECT 0.860 105.020 142.240 106.100 ;
        RECT 0.860 104.980 141.940 105.020 ;
        RECT 0.560 103.860 141.940 104.980 ;
        RECT 0.560 102.780 142.240 103.860 ;
        RECT 0.560 101.660 141.940 102.780 ;
        RECT 0.860 101.620 141.940 101.660 ;
        RECT 0.860 100.540 142.240 101.620 ;
        RECT 0.860 100.500 141.940 100.540 ;
        RECT 0.560 99.380 141.940 100.500 ;
        RECT 0.560 98.300 142.240 99.380 ;
        RECT 0.560 97.180 141.940 98.300 ;
        RECT 0.860 97.140 141.940 97.180 ;
        RECT 0.860 96.060 142.240 97.140 ;
        RECT 0.860 96.020 141.940 96.060 ;
        RECT 0.560 94.900 141.940 96.020 ;
        RECT 0.560 93.820 142.240 94.900 ;
        RECT 0.560 92.700 141.940 93.820 ;
        RECT 0.860 92.660 141.940 92.700 ;
        RECT 0.860 91.580 142.240 92.660 ;
        RECT 0.860 91.540 141.940 91.580 ;
        RECT 0.560 90.420 141.940 91.540 ;
        RECT 0.560 89.340 142.240 90.420 ;
        RECT 0.560 88.220 141.940 89.340 ;
        RECT 0.860 88.180 141.940 88.220 ;
        RECT 0.860 87.100 142.240 88.180 ;
        RECT 0.860 87.060 141.940 87.100 ;
        RECT 0.560 85.940 141.940 87.060 ;
        RECT 0.560 84.860 142.240 85.940 ;
        RECT 0.560 83.740 141.940 84.860 ;
        RECT 0.860 83.700 141.940 83.740 ;
        RECT 0.860 82.620 142.240 83.700 ;
        RECT 0.860 82.580 141.940 82.620 ;
        RECT 0.560 81.460 141.940 82.580 ;
        RECT 0.560 80.380 142.240 81.460 ;
        RECT 0.560 79.260 141.940 80.380 ;
        RECT 0.860 79.220 141.940 79.260 ;
        RECT 0.860 78.140 142.240 79.220 ;
        RECT 0.860 78.100 141.940 78.140 ;
        RECT 0.560 76.980 141.940 78.100 ;
        RECT 0.560 75.900 142.240 76.980 ;
        RECT 0.560 74.780 141.940 75.900 ;
        RECT 0.860 74.740 141.940 74.780 ;
        RECT 0.860 73.660 142.240 74.740 ;
        RECT 0.860 73.620 141.940 73.660 ;
        RECT 0.560 72.500 141.940 73.620 ;
        RECT 0.560 71.420 142.240 72.500 ;
        RECT 0.560 70.300 141.940 71.420 ;
        RECT 0.860 70.260 141.940 70.300 ;
        RECT 0.860 69.180 142.240 70.260 ;
        RECT 0.860 69.140 141.940 69.180 ;
        RECT 0.560 68.020 141.940 69.140 ;
        RECT 0.560 66.940 142.240 68.020 ;
        RECT 0.560 65.820 141.940 66.940 ;
        RECT 0.860 65.780 141.940 65.820 ;
        RECT 0.860 64.700 142.240 65.780 ;
        RECT 0.860 64.660 141.940 64.700 ;
        RECT 0.560 63.540 141.940 64.660 ;
        RECT 0.560 62.460 142.240 63.540 ;
        RECT 0.560 61.340 141.940 62.460 ;
        RECT 0.860 61.300 141.940 61.340 ;
        RECT 0.860 60.220 142.240 61.300 ;
        RECT 0.860 60.180 141.940 60.220 ;
        RECT 0.560 59.060 141.940 60.180 ;
        RECT 0.560 57.980 142.240 59.060 ;
        RECT 0.560 56.860 141.940 57.980 ;
        RECT 0.860 56.820 141.940 56.860 ;
        RECT 0.860 55.740 142.240 56.820 ;
        RECT 0.860 55.700 141.940 55.740 ;
        RECT 0.560 54.580 141.940 55.700 ;
        RECT 0.560 53.500 142.240 54.580 ;
        RECT 0.560 52.380 141.940 53.500 ;
        RECT 0.860 52.340 141.940 52.380 ;
        RECT 0.860 51.260 142.240 52.340 ;
        RECT 0.860 51.220 141.940 51.260 ;
        RECT 0.560 50.100 141.940 51.220 ;
        RECT 0.560 49.020 142.240 50.100 ;
        RECT 0.560 47.900 141.940 49.020 ;
        RECT 0.860 47.860 141.940 47.900 ;
        RECT 0.860 46.780 142.240 47.860 ;
        RECT 0.860 46.740 141.940 46.780 ;
        RECT 0.560 45.620 141.940 46.740 ;
        RECT 0.560 44.540 142.240 45.620 ;
        RECT 0.560 43.420 141.940 44.540 ;
        RECT 0.860 43.380 141.940 43.420 ;
        RECT 0.860 42.300 142.240 43.380 ;
        RECT 0.860 42.260 141.940 42.300 ;
        RECT 0.560 41.140 141.940 42.260 ;
        RECT 0.560 40.060 142.240 41.140 ;
        RECT 0.560 38.940 141.940 40.060 ;
        RECT 0.860 38.900 141.940 38.940 ;
        RECT 0.860 37.820 142.240 38.900 ;
        RECT 0.860 37.780 141.940 37.820 ;
        RECT 0.560 36.660 141.940 37.780 ;
        RECT 0.560 35.580 142.240 36.660 ;
        RECT 0.560 34.460 141.940 35.580 ;
        RECT 0.860 34.420 141.940 34.460 ;
        RECT 0.860 33.340 142.240 34.420 ;
        RECT 0.860 33.300 141.940 33.340 ;
        RECT 0.560 32.180 141.940 33.300 ;
        RECT 0.560 31.100 142.240 32.180 ;
        RECT 0.560 29.980 141.940 31.100 ;
        RECT 0.860 29.940 141.940 29.980 ;
        RECT 0.860 28.860 142.240 29.940 ;
        RECT 0.860 28.820 141.940 28.860 ;
        RECT 0.560 27.700 141.940 28.820 ;
        RECT 0.560 26.620 142.240 27.700 ;
        RECT 0.560 25.500 141.940 26.620 ;
        RECT 0.860 25.460 141.940 25.500 ;
        RECT 0.860 24.380 142.240 25.460 ;
        RECT 0.860 24.340 141.940 24.380 ;
        RECT 0.560 23.220 141.940 24.340 ;
        RECT 0.560 22.140 142.240 23.220 ;
        RECT 0.560 21.020 141.940 22.140 ;
        RECT 0.860 20.980 141.940 21.020 ;
        RECT 0.860 19.900 142.240 20.980 ;
        RECT 0.860 19.860 141.940 19.900 ;
        RECT 0.560 18.740 141.940 19.860 ;
        RECT 0.560 17.660 142.240 18.740 ;
        RECT 0.560 16.540 141.940 17.660 ;
        RECT 0.860 16.500 141.940 16.540 ;
        RECT 0.860 15.420 142.240 16.500 ;
        RECT 0.860 15.380 141.940 15.420 ;
        RECT 0.560 14.260 141.940 15.380 ;
        RECT 0.560 13.180 142.240 14.260 ;
        RECT 0.560 12.060 141.940 13.180 ;
        RECT 0.860 12.020 141.940 12.060 ;
        RECT 0.860 10.940 142.240 12.020 ;
        RECT 0.860 10.900 141.940 10.940 ;
        RECT 0.560 9.780 141.940 10.900 ;
        RECT 0.560 8.700 142.240 9.780 ;
        RECT 0.560 7.540 141.940 8.700 ;
        RECT 0.560 6.460 142.240 7.540 ;
        RECT 0.560 5.300 141.940 6.460 ;
        RECT 0.560 4.220 142.240 5.300 ;
        RECT 0.560 3.060 141.940 4.220 ;
        RECT 0.560 1.980 142.240 3.060 ;
        RECT 0.560 0.820 141.940 1.980 ;
        RECT 0.560 0.700 142.240 0.820 ;
      LAYER Metal4 ;
        RECT 6.300 1.770 18.580 279.910 ;
        RECT 20.780 1.770 21.880 279.910 ;
        RECT 24.080 1.770 118.580 279.910 ;
        RECT 120.780 1.770 121.880 279.910 ;
        RECT 124.080 1.770 137.620 279.910 ;
  END
END W_IO4
END LIBRARY

