* NGSPICE file created from S_term_SRAM.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

.subckt S_term_SRAM FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0]
+ N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10]
+ N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4]
+ N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3]
+ S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0]
+ S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10]
+ S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4]
+ S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] UserCLK UserCLKo VDD VSS
XFILLER_13_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_83_ S4END[4] net75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_66_ S2END[5] net67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_49_ FrameStrobe[17] net41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput42 net42 FrameStrobe_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput20 net20 FrameData_O[27] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput75 net75 N4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput64 net64 N2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput31 net31 FrameData_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput7 net7 FrameData_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput53 net53 N1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput86 net86 N4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_13_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_82_ S4END[5] net74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_12_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_65_ S2END[6] net66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_5_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Right_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_48_ FrameStrobe[16] net40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_15_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Right_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput76 net76 N4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput87 net87 N4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput32 net32 FrameData_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput8 net8 FrameData_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput10 net10 FrameData_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput54 net54 N1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput21 net21 FrameData_O[28] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput43 net43 FrameStrobe_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput65 net65 N2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_81_ S4END[6] net88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_8_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_64_ S2END[7] net65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_5_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_47_ FrameStrobe[15] net39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput33 net33 FrameStrobe_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput44 net44 FrameStrobe_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput77 net77 N4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput22 net22 FrameData_O[29] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput9 net9 FrameData_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput11 net11 FrameData_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput55 net55 N1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput66 net66 N2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput88 net88 N4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_11_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_80_ S4END[7] net87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_12_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_63_ S2MID[0] net64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_2_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_46_ FrameStrobe[14] net38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_12_Left_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_29_ FrameData[29] net22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput45 net45 FrameStrobe_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput78 net78 N4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput34 net34 FrameStrobe_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput23 net23 FrameData_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput12 net12 FrameData_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput56 net56 N1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput67 net67 N2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput89 net89 UserCLKo VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_15_Left_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_0_Left_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_62_ S2MID[1] net63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_45_ FrameStrobe[13] net37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_1_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_28_ FrameData[28] net21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput57 net57 N2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_15_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput24 net24 FrameData_O[30] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput46 net46 FrameStrobe_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput13 net13 FrameData_O[20] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput35 net35 FrameStrobe_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput79 net79 N4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput68 net68 N2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_13_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_61_ S2MID[2] net62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_2_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_44_ FrameStrobe[12] net36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_1_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_27_ FrameData[27] net20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_10_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput36 net36 FrameStrobe_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput47 net47 FrameStrobe_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput69 net69 N2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput58 net58 N2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput14 net14 FrameData_O[21] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput25 net25 FrameData_O[31] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_13_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_60_ S2MID[3] net61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_13_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_43_ FrameStrobe[11] net35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_26_ FrameData[26] net19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_10_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09_ FrameData[9] net32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput59 net59 N2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput15 net15 FrameData_O[22] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput37 net37 FrameStrobe_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_1_Right_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput26 net26 FrameData_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput48 net48 FrameStrobe_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_7_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_13_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_42_ FrameStrobe[10] net34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_25_ FrameData[25] net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_7_Left_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_10_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08_ FrameData[8] net31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput49 net49 FrameStrobe_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput16 net16 FrameData_O[23] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput27 net27 FrameData_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput38 net38 FrameStrobe_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_15_Right_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_13_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_41_ FrameStrobe[9] net52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_24_ FrameData[24] net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_10_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput39 net39 FrameStrobe_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07_ FrameData[7] net30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput28 net28 FrameData_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput17 net17 FrameData_O[24] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_15_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_40_ FrameStrobe[8] net51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_0_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_23_ FrameData[23] net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06_ FrameData[6] net29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput29 net29 FrameData_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput18 net18 FrameData_O[25] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_5_Right_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_22_ FrameData[22] net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05_ FrameData[5] net28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput19 net19 FrameData_O[26] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_15_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_11_Right_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_21_ FrameData[21] net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04_ FrameData[4] net27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_11_Left_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_14_Left_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_20_ FrameData[20] net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_03_ FrameData[3] net26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_6_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_3_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_9_Right_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_79_ S4END[8] net86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_6_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_02_ FrameData[2] net23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_8_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_3_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_78_ S4END[9] net85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_6_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_01_ FrameData[1] net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_2_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_0_Right_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_3_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Left_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_77_ S4END[10] net84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_6_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_00_ FrameData[0] net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_15_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_6_Left_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_76_ S4END[11] net83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_59_ S2MID[4] net60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_75_ S4END[12] net82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_14_Right_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_58_ S2MID[5] net59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_15_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Right_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_74_ S4END[13] net81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_1_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_57_ S2MID[6] net58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_15_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_73_ S4END[14] net80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_56_ S2MID[7] net57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_39_ FrameStrobe[7] net50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_7_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Left_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_72_ S4END[15] net73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_55_ S1END[0] net56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_10_Right_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_38_ FrameStrobe[6] net49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_8_Right_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_71_ S2END[0] net72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_54_ S1END[1] net55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_11_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_37_ FrameStrobe[5] net48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_70_ S2END[1] net71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_53_ S1END[2] net54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_11_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_36_ FrameStrobe[4] net47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_19_ FrameData[19] net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_5_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_2_Left_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_52_ S1END[3] net53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_11_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_35_ FrameStrobe[3] net46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_5_Left_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_18_ FrameData[18] net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_51_ FrameStrobe[19] net43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_34_ FrameStrobe[2] net45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_17_ FrameData[17] net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_13_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_50_ FrameStrobe[18] net42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_33_ FrameStrobe[1] net44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16_ FrameData[16] net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_3_Right_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_32_ FrameStrobe[0] net33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15_ FrameData[15] net7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_9_Left_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_13_Right_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_5_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_31_ FrameData[31] net25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14_ FrameData[14] net6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_4_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_30_ FrameData[30] net24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13_ FrameData[13] net5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_7_Right_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_5_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12_ FrameData[12] net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput1 net1 FrameData_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput80 net80 N4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_7_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_88_ UserCLK net89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11_ FrameData[11] net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_13_Left_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput81 net81 N4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput2 net2 FrameData_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_11_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput70 net70 N2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_14_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_1_Left_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_87_ S4END[0] net79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10_ FrameData[10] net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_5_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Left_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput71 net71 N2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_2_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput3 net3 FrameData_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput60 net60 N2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput82 net82 N4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_9_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_86_ S4END[1] net78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_69_ S2END[2] net70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_5_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput50 net50 FrameStrobe_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_2_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput4 net4 FrameData_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput61 net61 N2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput72 net72 N2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput83 net83 N4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_13_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_85_ S4END[2] net77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_68_ S2END[3] net69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_2_Right_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput40 net40 FrameStrobe_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput51 net51 FrameStrobe_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput84 net84 N4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_2_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput5 net5 FrameData_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput62 net62 N2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput73 net73 N4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_84_ S4END[3] net76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_67_ S2END[4] net68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_8_Left_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput41 net41 FrameStrobe_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput52 net52 FrameStrobe_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput30 net30 FrameData_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_1_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput6 net6 FrameData_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput63 net63 N2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput85 net85 N4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput74 net74 N4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

