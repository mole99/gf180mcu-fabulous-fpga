magic
tech gf180mcuD
magscale 1 5
timestamp 1764970794
<< metal1 >>
rect 336 6677 31864 6694
rect 336 6651 2233 6677
rect 2259 6651 2285 6677
rect 2311 6651 2337 6677
rect 2363 6651 12233 6677
rect 12259 6651 12285 6677
rect 12311 6651 12337 6677
rect 12363 6651 22233 6677
rect 22259 6651 22285 6677
rect 22311 6651 22337 6677
rect 22363 6651 31864 6677
rect 336 6634 31864 6651
rect 7519 6593 7545 6599
rect 1577 6567 1583 6593
rect 1609 6567 1615 6593
rect 7519 6561 7545 6567
rect 9143 6593 9169 6599
rect 9143 6561 9169 6567
rect 10599 6593 10625 6599
rect 10599 6561 10625 6567
rect 12223 6593 12249 6599
rect 12223 6561 12249 6567
rect 13231 6593 13257 6599
rect 13231 6561 13257 6567
rect 31263 6593 31289 6599
rect 31263 6561 31289 6567
rect 5105 6511 5111 6537
rect 5137 6511 5143 6537
rect 6449 6511 6455 6537
rect 6481 6511 6487 6537
rect 7233 6511 7239 6537
rect 7265 6511 7271 6537
rect 1751 6481 1777 6487
rect 3649 6455 3655 6481
rect 3681 6455 3687 6481
rect 6841 6455 6847 6481
rect 6873 6455 6879 6481
rect 8857 6455 8863 6481
rect 8889 6455 8895 6481
rect 10313 6455 10319 6481
rect 10345 6455 10351 6481
rect 11937 6455 11943 6481
rect 11969 6455 11975 6481
rect 12945 6455 12951 6481
rect 12977 6455 12983 6481
rect 15297 6455 15303 6481
rect 15329 6455 15335 6481
rect 16753 6455 16759 6481
rect 16785 6455 16791 6481
rect 18265 6455 18271 6481
rect 18297 6455 18303 6481
rect 21121 6455 21127 6481
rect 21153 6455 21159 6481
rect 22577 6455 22583 6481
rect 22609 6455 22615 6481
rect 24033 6455 24039 6481
rect 24065 6455 24071 6481
rect 26889 6455 26895 6481
rect 26921 6455 26927 6481
rect 28401 6455 28407 6481
rect 28433 6455 28439 6481
rect 29745 6455 29751 6481
rect 29777 6455 29783 6481
rect 30081 6455 30087 6481
rect 30113 6455 30119 6481
rect 30977 6455 30983 6481
rect 31009 6455 31015 6481
rect 1751 6449 1777 6455
rect 3151 6425 3177 6431
rect 3151 6393 3177 6399
rect 4607 6425 4633 6431
rect 4607 6393 4633 6399
rect 14799 6425 14825 6431
rect 14799 6393 14825 6399
rect 16255 6425 16281 6431
rect 16255 6393 16281 6399
rect 17767 6425 17793 6431
rect 17767 6393 17793 6399
rect 20623 6425 20649 6431
rect 20623 6393 20649 6399
rect 22079 6425 22105 6431
rect 22079 6393 22105 6399
rect 23535 6425 23561 6431
rect 23535 6393 23561 6399
rect 26391 6425 26417 6431
rect 26391 6393 26417 6399
rect 27903 6425 27929 6431
rect 27903 6393 27929 6399
rect 29359 6425 29385 6431
rect 29359 6393 29385 6399
rect 30591 6369 30617 6375
rect 30591 6337 30617 6343
rect 336 6285 31864 6302
rect 336 6259 1903 6285
rect 1929 6259 1955 6285
rect 1981 6259 2007 6285
rect 2033 6259 11903 6285
rect 11929 6259 11955 6285
rect 11981 6259 12007 6285
rect 12033 6259 21903 6285
rect 21929 6259 21955 6285
rect 21981 6259 22007 6285
rect 22033 6259 31864 6285
rect 336 6242 31864 6259
rect 19167 6201 19193 6207
rect 19167 6169 19193 6175
rect 24991 6201 25017 6207
rect 24991 6169 25017 6175
rect 29527 6201 29553 6207
rect 29527 6169 29553 6175
rect 30759 6145 30785 6151
rect 6897 6119 6903 6145
rect 6929 6119 6935 6145
rect 8521 6119 8527 6145
rect 8553 6119 8559 6145
rect 30759 6113 30785 6119
rect 31543 6145 31569 6151
rect 31543 6113 31569 6119
rect 7127 6089 7153 6095
rect 7127 6057 7153 6063
rect 8751 6089 8777 6095
rect 8751 6057 8777 6063
rect 17319 6089 17345 6095
rect 17319 6057 17345 6063
rect 18607 6089 18633 6095
rect 18607 6057 18633 6063
rect 20847 6089 20873 6095
rect 20847 6057 20873 6063
rect 21127 6089 21153 6095
rect 30249 6063 30255 6089
rect 30281 6063 30287 6089
rect 21127 6057 21153 6063
rect 16759 6033 16785 6039
rect 16759 6001 16785 6007
rect 17599 6033 17625 6039
rect 17599 6001 17625 6007
rect 18887 6033 18913 6039
rect 20679 6033 20705 6039
rect 27567 6033 27593 6039
rect 19665 6007 19671 6033
rect 19697 6007 19703 6033
rect 25489 6007 25495 6033
rect 25521 6007 25527 6033
rect 29017 6007 29023 6033
rect 29049 6007 29055 6033
rect 31033 6007 31039 6033
rect 31065 6007 31071 6033
rect 18887 6001 18913 6007
rect 20679 6001 20705 6007
rect 27567 6001 27593 6007
rect 16479 5977 16505 5983
rect 16479 5945 16505 5951
rect 20399 5977 20425 5983
rect 20399 5945 20425 5951
rect 27847 5977 27873 5983
rect 27847 5945 27873 5951
rect 336 5893 31864 5910
rect 336 5867 2233 5893
rect 2259 5867 2285 5893
rect 2311 5867 2337 5893
rect 2363 5867 12233 5893
rect 12259 5867 12285 5893
rect 12311 5867 12337 5893
rect 12363 5867 22233 5893
rect 22259 5867 22285 5893
rect 22311 5867 22337 5893
rect 22363 5867 31864 5893
rect 336 5850 31864 5867
rect 9927 5753 9953 5759
rect 9927 5721 9953 5727
rect 11047 5753 11073 5759
rect 11047 5721 11073 5727
rect 12279 5753 12305 5759
rect 12279 5721 12305 5727
rect 14967 5753 14993 5759
rect 14967 5721 14993 5727
rect 16199 5753 16225 5759
rect 16199 5721 16225 5727
rect 10207 5697 10233 5703
rect 10207 5665 10233 5671
rect 11327 5697 11353 5703
rect 11327 5665 11353 5671
rect 12559 5697 12585 5703
rect 12559 5665 12585 5671
rect 12783 5697 12809 5703
rect 12783 5665 12809 5671
rect 14687 5697 14713 5703
rect 14687 5665 14713 5671
rect 16479 5697 16505 5703
rect 16479 5665 16505 5671
rect 19447 5697 19473 5703
rect 19447 5665 19473 5671
rect 21743 5697 21769 5703
rect 29353 5671 29359 5697
rect 29385 5671 29391 5697
rect 30137 5671 30143 5697
rect 30169 5671 30175 5697
rect 30921 5671 30927 5697
rect 30953 5671 30959 5697
rect 21743 5665 21769 5671
rect 13063 5641 13089 5647
rect 13063 5609 13089 5615
rect 19727 5641 19753 5647
rect 19727 5609 19753 5615
rect 22023 5641 22049 5647
rect 22023 5609 22049 5615
rect 29863 5641 29889 5647
rect 29863 5609 29889 5615
rect 30647 5641 30673 5647
rect 31369 5615 31375 5641
rect 31401 5615 31407 5641
rect 30647 5609 30673 5615
rect 336 5501 31864 5518
rect 336 5475 1903 5501
rect 1929 5475 1955 5501
rect 1981 5475 2007 5501
rect 2033 5475 11903 5501
rect 11929 5475 11955 5501
rect 11981 5475 12007 5501
rect 12033 5475 21903 5501
rect 21929 5475 21955 5501
rect 21981 5475 22007 5501
rect 22033 5475 31864 5501
rect 336 5458 31864 5475
rect 18719 5361 18745 5367
rect 18719 5329 18745 5335
rect 18489 5279 18495 5305
rect 18521 5279 18527 5305
rect 31089 5279 31095 5305
rect 31121 5279 31127 5305
rect 15919 5249 15945 5255
rect 30249 5223 30255 5249
rect 30281 5223 30287 5249
rect 30641 5223 30647 5249
rect 30673 5223 30679 5249
rect 31425 5223 31431 5249
rect 31457 5223 31463 5249
rect 15919 5217 15945 5223
rect 15639 5193 15665 5199
rect 15639 5161 15665 5167
rect 336 5109 31864 5126
rect 336 5083 2233 5109
rect 2259 5083 2285 5109
rect 2311 5083 2337 5109
rect 2363 5083 12233 5109
rect 12259 5083 12285 5109
rect 12311 5083 12337 5109
rect 12363 5083 22233 5109
rect 22259 5083 22285 5109
rect 22311 5083 22337 5109
rect 22363 5083 31864 5109
rect 336 5066 31864 5083
rect 16535 5025 16561 5031
rect 16535 4993 16561 4999
rect 12783 4969 12809 4975
rect 12783 4937 12809 4943
rect 18719 4969 18745 4975
rect 30529 4943 30535 4969
rect 30561 4943 30567 4969
rect 18719 4937 18745 4943
rect 4159 4913 4185 4919
rect 4159 4881 4185 4887
rect 12503 4913 12529 4919
rect 18489 4887 18495 4913
rect 18521 4887 18527 4913
rect 30137 4887 30143 4913
rect 30169 4887 30175 4913
rect 30921 4887 30927 4913
rect 30953 4887 30959 4913
rect 12503 4881 12529 4887
rect 3929 4831 3935 4857
rect 3961 4831 3967 4857
rect 16753 4831 16759 4857
rect 16785 4831 16791 4857
rect 31369 4831 31375 4857
rect 31401 4831 31407 4857
rect 336 4717 31864 4734
rect 336 4691 1903 4717
rect 1929 4691 1955 4717
rect 1981 4691 2007 4717
rect 2033 4691 11903 4717
rect 11929 4691 11955 4717
rect 11981 4691 12007 4717
rect 12033 4691 21903 4717
rect 21929 4691 21955 4717
rect 21981 4691 22007 4717
rect 22033 4691 31864 4717
rect 336 4674 31864 4691
rect 30759 4633 30785 4639
rect 30759 4601 30785 4607
rect 14519 4577 14545 4583
rect 14519 4545 14545 4551
rect 20287 4577 20313 4583
rect 20287 4545 20313 4551
rect 11663 4521 11689 4527
rect 17263 4521 17289 4527
rect 14289 4495 14295 4521
rect 14321 4495 14327 4521
rect 30249 4495 30255 4521
rect 30281 4495 30287 4521
rect 31089 4495 31095 4521
rect 31121 4495 31127 4521
rect 11663 4489 11689 4495
rect 17263 4489 17289 4495
rect 967 4465 993 4471
rect 967 4433 993 4439
rect 11943 4465 11969 4471
rect 31425 4439 31431 4465
rect 31457 4439 31463 4465
rect 11943 4433 11969 4439
rect 1247 4409 1273 4415
rect 1247 4377 1273 4383
rect 16983 4409 17009 4415
rect 16983 4377 17009 4383
rect 20007 4409 20033 4415
rect 20007 4377 20033 4383
rect 336 4325 31864 4342
rect 336 4299 2233 4325
rect 2259 4299 2285 4325
rect 2311 4299 2337 4325
rect 2363 4299 12233 4325
rect 12259 4299 12285 4325
rect 12311 4299 12337 4325
rect 12363 4299 22233 4325
rect 22259 4299 22285 4325
rect 22311 4299 22337 4325
rect 22363 4299 31864 4325
rect 336 4282 31864 4299
rect 18887 4241 18913 4247
rect 18887 4209 18913 4215
rect 19167 4185 19193 4191
rect 19167 4153 19193 4159
rect 30479 4129 30505 4135
rect 30921 4103 30927 4129
rect 30953 4103 30959 4129
rect 30479 4097 30505 4103
rect 30697 4047 30703 4073
rect 30729 4047 30735 4073
rect 31431 4017 31457 4023
rect 31431 3985 31457 3991
rect 336 3933 31864 3950
rect 336 3907 1903 3933
rect 1929 3907 1955 3933
rect 1981 3907 2007 3933
rect 2033 3907 11903 3933
rect 11929 3907 11955 3933
rect 11981 3907 12007 3933
rect 12033 3907 21903 3933
rect 21929 3907 21955 3933
rect 21981 3907 22007 3933
rect 22033 3907 31864 3933
rect 336 3890 31864 3907
rect 31543 3849 31569 3855
rect 31543 3817 31569 3823
rect 6119 3793 6145 3799
rect 6119 3761 6145 3767
rect 13063 3793 13089 3799
rect 13063 3761 13089 3767
rect 17487 3793 17513 3799
rect 17487 3761 17513 3767
rect 30759 3793 30785 3799
rect 30759 3761 30785 3767
rect 4439 3737 4465 3743
rect 12783 3737 12809 3743
rect 5889 3711 5895 3737
rect 5921 3711 5927 3737
rect 4439 3705 4465 3711
rect 12783 3705 12809 3711
rect 13679 3737 13705 3743
rect 13679 3705 13705 3711
rect 14743 3737 14769 3743
rect 14743 3705 14769 3711
rect 15023 3737 15049 3743
rect 15023 3705 15049 3711
rect 17767 3737 17793 3743
rect 17767 3705 17793 3711
rect 20567 3737 20593 3743
rect 29409 3711 29415 3737
rect 29441 3711 29447 3737
rect 31089 3711 31095 3737
rect 31121 3711 31127 3737
rect 20567 3705 20593 3711
rect 10039 3681 10065 3687
rect 10039 3649 10065 3655
rect 10431 3681 10457 3687
rect 10431 3649 10457 3655
rect 13959 3681 13985 3687
rect 13959 3649 13985 3655
rect 18495 3681 18521 3687
rect 18495 3649 18521 3655
rect 20847 3681 20873 3687
rect 20847 3649 20873 3655
rect 29639 3681 29665 3687
rect 30249 3655 30255 3681
rect 30281 3655 30287 3681
rect 29639 3649 29665 3655
rect 4719 3625 4745 3631
rect 4719 3593 4745 3599
rect 9759 3625 9785 3631
rect 9759 3593 9785 3599
rect 10711 3625 10737 3631
rect 10711 3593 10737 3599
rect 18215 3625 18241 3631
rect 18215 3593 18241 3599
rect 336 3541 31864 3558
rect 336 3515 2233 3541
rect 2259 3515 2285 3541
rect 2311 3515 2337 3541
rect 2363 3515 12233 3541
rect 12259 3515 12285 3541
rect 12311 3515 12337 3541
rect 12363 3515 22233 3541
rect 22259 3515 22285 3541
rect 22311 3515 22337 3541
rect 22363 3515 31864 3541
rect 336 3498 31864 3515
rect 15639 3401 15665 3407
rect 15639 3369 15665 3375
rect 2647 3345 2673 3351
rect 2647 3313 2673 3319
rect 6455 3345 6481 3351
rect 15359 3345 15385 3351
rect 6673 3319 6679 3345
rect 6705 3319 6711 3345
rect 6455 3313 6481 3319
rect 15359 3313 15385 3319
rect 24487 3345 24513 3351
rect 30137 3319 30143 3345
rect 30169 3319 30175 3345
rect 30921 3319 30927 3345
rect 30953 3319 30959 3345
rect 24487 3313 24513 3319
rect 31431 3289 31457 3295
rect 2417 3263 2423 3289
rect 2449 3263 2455 3289
rect 24705 3263 24711 3289
rect 24737 3263 24743 3289
rect 31431 3257 31457 3263
rect 30647 3233 30673 3239
rect 30647 3201 30673 3207
rect 336 3149 31864 3166
rect 336 3123 1903 3149
rect 1929 3123 1955 3149
rect 1981 3123 2007 3149
rect 2033 3123 11903 3149
rect 11929 3123 11955 3149
rect 11981 3123 12007 3149
rect 12033 3123 21903 3149
rect 21929 3123 21955 3149
rect 21981 3123 22007 3149
rect 22033 3123 31864 3149
rect 336 3106 31864 3123
rect 31543 3065 31569 3071
rect 31543 3033 31569 3039
rect 20679 3009 20705 3015
rect 30809 2983 30815 3009
rect 30841 2983 30847 3009
rect 20679 2977 20705 2983
rect 17543 2953 17569 2959
rect 17543 2921 17569 2927
rect 20399 2953 20425 2959
rect 20399 2921 20425 2927
rect 22527 2953 22553 2959
rect 22527 2921 22553 2927
rect 23423 2953 23449 2959
rect 23423 2921 23449 2927
rect 25439 2953 25465 2959
rect 31089 2927 31095 2953
rect 31121 2927 31127 2953
rect 25439 2921 25465 2927
rect 17823 2897 17849 2903
rect 17823 2865 17849 2871
rect 22807 2897 22833 2903
rect 22807 2865 22833 2871
rect 23703 2897 23729 2903
rect 23703 2865 23729 2871
rect 25719 2897 25745 2903
rect 25719 2865 25745 2871
rect 27063 2897 27089 2903
rect 27063 2865 27089 2871
rect 26783 2841 26809 2847
rect 26783 2809 26809 2815
rect 30591 2841 30617 2847
rect 30591 2809 30617 2815
rect 336 2757 31864 2774
rect 336 2731 2233 2757
rect 2259 2731 2285 2757
rect 2311 2731 2337 2757
rect 2363 2731 12233 2757
rect 12259 2731 12285 2757
rect 12311 2731 12337 2757
rect 12363 2731 22233 2757
rect 22259 2731 22285 2757
rect 22311 2731 22337 2757
rect 22363 2731 31864 2757
rect 336 2714 31864 2731
rect 11327 2673 11353 2679
rect 11327 2641 11353 2647
rect 13119 2673 13145 2679
rect 13119 2641 13145 2647
rect 16983 2673 17009 2679
rect 16983 2641 17009 2647
rect 22191 2673 22217 2679
rect 22191 2641 22217 2647
rect 27399 2673 27425 2679
rect 27399 2641 27425 2647
rect 911 2617 937 2623
rect 911 2585 937 2591
rect 4439 2617 4465 2623
rect 4439 2585 4465 2591
rect 10319 2617 10345 2623
rect 10319 2585 10345 2591
rect 10599 2617 10625 2623
rect 10599 2585 10625 2591
rect 13399 2617 13425 2623
rect 13399 2585 13425 2591
rect 19167 2617 19193 2623
rect 19167 2585 19193 2591
rect 19447 2617 19473 2623
rect 21625 2591 21631 2617
rect 21657 2591 21663 2617
rect 30137 2591 30143 2617
rect 30169 2591 30175 2617
rect 30921 2591 30927 2617
rect 30953 2591 30959 2617
rect 31313 2591 31319 2617
rect 31345 2591 31351 2617
rect 19447 2585 19473 2591
rect 1191 2561 1217 2567
rect 1191 2529 1217 2535
rect 4719 2561 4745 2567
rect 4719 2529 4745 2535
rect 11047 2561 11073 2567
rect 11047 2529 11073 2535
rect 21799 2561 21825 2567
rect 21799 2529 21825 2535
rect 22471 2561 22497 2567
rect 22471 2529 22497 2535
rect 27679 2561 27705 2567
rect 30529 2535 30535 2561
rect 30561 2535 30567 2561
rect 27679 2529 27705 2535
rect 10767 2505 10793 2511
rect 10767 2473 10793 2479
rect 11607 2505 11633 2511
rect 17201 2479 17207 2505
rect 17233 2479 17239 2505
rect 11607 2473 11633 2479
rect 336 2365 31864 2382
rect 336 2339 1903 2365
rect 1929 2339 1955 2365
rect 1981 2339 2007 2365
rect 2033 2339 11903 2365
rect 11929 2339 11955 2365
rect 11981 2339 12007 2365
rect 12033 2339 21903 2365
rect 21929 2339 21955 2365
rect 21981 2339 22007 2365
rect 22033 2339 31864 2365
rect 336 2322 31864 2339
rect 31543 2281 31569 2287
rect 31543 2249 31569 2255
rect 24095 2225 24121 2231
rect 7681 2199 7687 2225
rect 7713 2199 7719 2225
rect 9193 2199 9199 2225
rect 9225 2199 9231 2225
rect 11713 2199 11719 2225
rect 11745 2199 11751 2225
rect 13897 2199 13903 2225
rect 13929 2199 13935 2225
rect 21737 2199 21743 2225
rect 21769 2199 21775 2225
rect 23585 2199 23591 2225
rect 23617 2199 23623 2225
rect 29577 2199 29583 2225
rect 29609 2199 29615 2225
rect 24095 2193 24121 2199
rect 16479 2169 16505 2175
rect 16479 2137 16505 2143
rect 18831 2169 18857 2175
rect 18831 2137 18857 2143
rect 21519 2169 21545 2175
rect 24313 2143 24319 2169
rect 24345 2143 24351 2169
rect 25097 2143 25103 2169
rect 25129 2143 25135 2169
rect 29409 2143 29415 2169
rect 29441 2143 29447 2169
rect 30249 2143 30255 2169
rect 30281 2143 30287 2169
rect 31089 2143 31095 2169
rect 31121 2143 31127 2169
rect 21519 2137 21545 2143
rect 11495 2113 11521 2119
rect 11495 2081 11521 2087
rect 12895 2113 12921 2119
rect 12895 2081 12921 2087
rect 15975 2113 16001 2119
rect 15975 2081 16001 2087
rect 16255 2113 16281 2119
rect 16255 2081 16281 2087
rect 16759 2113 16785 2119
rect 16759 2081 16785 2087
rect 19111 2113 19137 2119
rect 19111 2081 19137 2087
rect 20455 2113 20481 2119
rect 20455 2081 20481 2087
rect 21071 2113 21097 2119
rect 23921 2087 23927 2113
rect 23953 2087 23959 2113
rect 30641 2087 30647 2113
rect 30673 2087 30679 2113
rect 21071 2081 21097 2087
rect 7911 2057 7937 2063
rect 7911 2025 7937 2031
rect 8975 2057 9001 2063
rect 8975 2025 9001 2031
rect 12615 2057 12641 2063
rect 12615 2025 12641 2031
rect 13679 2057 13705 2063
rect 13679 2025 13705 2031
rect 20175 2057 20201 2063
rect 20175 2025 20201 2031
rect 20791 2057 20817 2063
rect 20791 2025 20817 2031
rect 25383 2057 25409 2063
rect 25383 2025 25409 2031
rect 336 1973 31864 1990
rect 336 1947 2233 1973
rect 2259 1947 2285 1973
rect 2311 1947 2337 1973
rect 2363 1947 12233 1973
rect 12259 1947 12285 1973
rect 12311 1947 12337 1973
rect 12363 1947 22233 1973
rect 22259 1947 22285 1973
rect 22311 1947 22337 1973
rect 22363 1947 31864 1973
rect 336 1930 31864 1947
rect 15639 1889 15665 1895
rect 15639 1857 15665 1863
rect 16199 1889 16225 1895
rect 16199 1857 16225 1863
rect 17935 1889 17961 1895
rect 17935 1857 17961 1863
rect 6007 1833 6033 1839
rect 6007 1801 6033 1807
rect 13959 1833 13985 1839
rect 15919 1833 15945 1839
rect 14121 1807 14127 1833
rect 14153 1807 14159 1833
rect 13959 1801 13985 1807
rect 15919 1801 15945 1807
rect 16479 1833 16505 1839
rect 25607 1833 25633 1839
rect 18377 1807 18383 1833
rect 18409 1807 18415 1833
rect 20729 1807 20735 1833
rect 20761 1807 20767 1833
rect 23081 1807 23087 1833
rect 23113 1807 23119 1833
rect 24033 1807 24039 1833
rect 24065 1807 24071 1833
rect 24817 1807 24823 1833
rect 24849 1807 24855 1833
rect 16479 1801 16505 1807
rect 25607 1801 25633 1807
rect 27959 1833 27985 1839
rect 27959 1801 27985 1807
rect 28463 1833 28489 1839
rect 30137 1807 30143 1833
rect 30169 1807 30175 1833
rect 30921 1807 30927 1833
rect 30953 1807 30959 1833
rect 28463 1801 28489 1807
rect 6287 1777 6313 1783
rect 6287 1745 6313 1751
rect 7015 1777 7041 1783
rect 15191 1777 15217 1783
rect 13729 1751 13735 1777
rect 13761 1751 13767 1777
rect 7015 1745 7041 1751
rect 15191 1745 15217 1751
rect 19167 1777 19193 1783
rect 25887 1777 25913 1783
rect 21457 1751 21463 1777
rect 21489 1751 21495 1777
rect 22297 1751 22303 1777
rect 22329 1751 22335 1777
rect 19167 1745 19193 1751
rect 25887 1745 25913 1751
rect 28239 1777 28265 1783
rect 28239 1745 28265 1751
rect 28743 1777 28769 1783
rect 28743 1745 28769 1751
rect 7295 1721 7321 1727
rect 7295 1689 7321 1695
rect 15471 1721 15497 1727
rect 15471 1689 15497 1695
rect 18215 1721 18241 1727
rect 18215 1689 18241 1695
rect 19447 1721 19473 1727
rect 19447 1689 19473 1695
rect 20231 1721 20257 1727
rect 20231 1689 20257 1695
rect 21015 1721 21041 1727
rect 21015 1689 21041 1695
rect 21799 1721 21825 1727
rect 30647 1721 30673 1727
rect 22745 1695 22751 1721
rect 22777 1695 22783 1721
rect 24369 1695 24375 1721
rect 24401 1695 24407 1721
rect 25265 1695 25271 1721
rect 25297 1695 25303 1721
rect 21799 1689 21825 1695
rect 30647 1689 30673 1695
rect 31431 1721 31457 1727
rect 31431 1689 31457 1695
rect 14407 1665 14433 1671
rect 14407 1633 14433 1639
rect 18663 1665 18689 1671
rect 18663 1633 18689 1639
rect 336 1581 31864 1598
rect 336 1555 1903 1581
rect 1929 1555 1955 1581
rect 1981 1555 2007 1581
rect 2033 1555 11903 1581
rect 11929 1555 11955 1581
rect 11981 1555 12007 1581
rect 12033 1555 21903 1581
rect 21929 1555 21955 1581
rect 21981 1555 22007 1581
rect 22033 1555 31864 1581
rect 336 1538 31864 1555
rect 31543 1497 31569 1503
rect 31543 1465 31569 1471
rect 22975 1441 23001 1447
rect 22975 1409 23001 1415
rect 26111 1441 26137 1447
rect 26111 1409 26137 1415
rect 26727 1441 26753 1447
rect 26727 1409 26753 1415
rect 25215 1385 25241 1391
rect 14345 1359 14351 1385
rect 14377 1359 14383 1385
rect 15969 1359 15975 1385
rect 16001 1359 16007 1385
rect 16809 1359 16815 1385
rect 16841 1359 16847 1385
rect 17257 1359 17263 1385
rect 17289 1359 17295 1385
rect 18153 1359 18159 1385
rect 18185 1359 18191 1385
rect 18937 1359 18943 1385
rect 18969 1359 18975 1385
rect 19721 1359 19727 1385
rect 19753 1359 19759 1385
rect 20505 1359 20511 1385
rect 20537 1359 20543 1385
rect 22577 1359 22583 1385
rect 22609 1359 22615 1385
rect 23473 1359 23479 1385
rect 23505 1359 23511 1385
rect 24481 1359 24487 1385
rect 24513 1359 24519 1385
rect 30249 1359 30255 1385
rect 30281 1359 30287 1385
rect 31089 1359 31095 1385
rect 31121 1359 31127 1385
rect 25215 1353 25241 1359
rect 911 1329 937 1335
rect 911 1297 937 1303
rect 13959 1329 13985 1335
rect 17039 1329 17065 1335
rect 21295 1329 21321 1335
rect 15129 1303 15135 1329
rect 15161 1303 15167 1329
rect 17649 1303 17655 1329
rect 17681 1303 17687 1329
rect 18545 1303 18551 1329
rect 18577 1303 18583 1329
rect 13959 1297 13985 1303
rect 17039 1297 17065 1303
rect 21295 1297 21321 1303
rect 21575 1329 21601 1335
rect 29359 1329 29385 1335
rect 22297 1303 22303 1329
rect 22329 1303 22335 1329
rect 23641 1303 23647 1329
rect 23673 1303 23679 1329
rect 30641 1303 30647 1329
rect 30673 1303 30679 1329
rect 21575 1297 21601 1303
rect 29359 1297 29385 1303
rect 1191 1273 1217 1279
rect 1191 1241 1217 1247
rect 13679 1273 13705 1279
rect 13679 1241 13705 1247
rect 14631 1273 14657 1279
rect 14631 1241 14657 1247
rect 15415 1273 15441 1279
rect 15415 1241 15441 1247
rect 16199 1273 16225 1279
rect 16199 1241 16225 1247
rect 19223 1273 19249 1279
rect 19223 1241 19249 1247
rect 20007 1273 20033 1279
rect 20007 1241 20033 1247
rect 20791 1273 20817 1279
rect 20791 1241 20817 1247
rect 23927 1273 23953 1279
rect 23927 1241 23953 1247
rect 24711 1273 24737 1279
rect 24711 1241 24737 1247
rect 25495 1273 25521 1279
rect 25495 1241 25521 1247
rect 26391 1273 26417 1279
rect 26391 1241 26417 1247
rect 27007 1273 27033 1279
rect 27007 1241 27033 1247
rect 29639 1273 29665 1279
rect 29639 1241 29665 1247
rect 336 1189 31864 1206
rect 336 1163 2233 1189
rect 2259 1163 2285 1189
rect 2311 1163 2337 1189
rect 2363 1163 12233 1189
rect 12259 1163 12285 1189
rect 12311 1163 12337 1189
rect 12363 1163 22233 1189
rect 22259 1163 22285 1189
rect 22311 1163 22337 1189
rect 22363 1163 31864 1189
rect 336 1146 31864 1163
rect 10543 1105 10569 1111
rect 10543 1073 10569 1079
rect 12839 1105 12865 1111
rect 12839 1073 12865 1079
rect 13287 1105 13313 1111
rect 13287 1073 13313 1079
rect 21183 1105 21209 1111
rect 21183 1073 21209 1079
rect 29639 1105 29665 1111
rect 29639 1073 29665 1079
rect 2367 1049 2393 1055
rect 2367 1017 2393 1023
rect 10823 1049 10849 1055
rect 23255 1049 23281 1055
rect 14513 1023 14519 1049
rect 14545 1023 14551 1049
rect 16361 1023 16367 1049
rect 16393 1023 16399 1049
rect 17145 1023 17151 1049
rect 17177 1023 17183 1049
rect 17929 1023 17935 1049
rect 17961 1023 17967 1049
rect 18713 1023 18719 1049
rect 18745 1023 18751 1049
rect 20897 1023 20903 1049
rect 20929 1023 20935 1049
rect 23081 1023 23087 1049
rect 23113 1023 23119 1049
rect 10823 1017 10849 1023
rect 23255 1017 23281 1023
rect 29191 1049 29217 1055
rect 29191 1017 29217 1023
rect 29919 1049 29945 1055
rect 30921 1023 30927 1049
rect 30953 1023 30959 1049
rect 29919 1017 29945 1023
rect 1191 993 1217 999
rect 1191 961 1217 967
rect 2647 993 2673 999
rect 2647 961 2673 967
rect 10375 993 10401 999
rect 10375 961 10401 967
rect 12615 993 12641 999
rect 19503 993 19529 999
rect 13729 967 13735 993
rect 13761 967 13767 993
rect 15409 967 15415 993
rect 15441 967 15447 993
rect 12615 961 12641 967
rect 19503 961 19529 967
rect 19783 993 19809 999
rect 29471 993 29497 999
rect 20113 967 20119 993
rect 20145 967 20151 993
rect 21737 967 21743 993
rect 21769 967 21775 993
rect 23473 967 23479 993
rect 23505 967 23511 993
rect 24033 967 24039 993
rect 24065 967 24071 993
rect 24873 967 24879 993
rect 24905 967 24911 993
rect 25713 967 25719 993
rect 25745 967 25751 993
rect 26441 967 26447 993
rect 26473 967 26479 993
rect 30137 967 30143 993
rect 30169 967 30175 993
rect 19783 961 19809 967
rect 29471 961 29497 967
rect 13119 937 13145 943
rect 961 911 967 937
rect 993 911 999 937
rect 10145 911 10151 937
rect 10177 911 10183 937
rect 12385 911 12391 937
rect 12417 911 12423 937
rect 13119 905 13145 911
rect 13567 937 13593 943
rect 18215 937 18241 943
rect 25887 937 25913 943
rect 14905 911 14911 937
rect 14937 911 14943 937
rect 22689 911 22695 937
rect 22721 911 22727 937
rect 24425 911 24431 937
rect 24457 911 24463 937
rect 25209 911 25215 937
rect 25241 911 25247 937
rect 13567 905 13593 911
rect 18215 905 18241 911
rect 25887 905 25913 911
rect 31431 937 31457 943
rect 31431 905 31457 911
rect 14239 881 14265 887
rect 14239 849 14265 855
rect 15583 881 15609 887
rect 15583 849 15609 855
rect 16647 881 16673 887
rect 16647 849 16673 855
rect 17431 881 17457 887
rect 17431 849 17457 855
rect 18999 881 19025 887
rect 18999 849 19025 855
rect 20399 881 20425 887
rect 20399 849 20425 855
rect 21967 881 21993 887
rect 21967 849 21993 855
rect 26671 881 26697 887
rect 26671 849 26697 855
rect 30647 881 30673 887
rect 30647 849 30673 855
rect 336 797 31864 814
rect 336 771 1903 797
rect 1929 771 1955 797
rect 1981 771 2007 797
rect 2033 771 11903 797
rect 11929 771 11955 797
rect 11981 771 12007 797
rect 12033 771 21903 797
rect 21929 771 21955 797
rect 21981 771 22007 797
rect 22033 771 31864 797
rect 336 754 31864 771
rect 31543 713 31569 719
rect 31543 681 31569 687
rect 14575 657 14601 663
rect 14575 625 14601 631
rect 15359 657 15385 663
rect 15359 625 15385 631
rect 16703 657 16729 663
rect 16703 625 16729 631
rect 22359 657 22385 663
rect 22359 625 22385 631
rect 29807 657 29833 663
rect 29807 625 29833 631
rect 30591 657 30617 663
rect 30591 625 30617 631
rect 12945 575 12951 601
rect 12977 575 12983 601
rect 14065 575 14071 601
rect 14097 575 14103 601
rect 14849 575 14855 601
rect 14881 575 14887 601
rect 15801 575 15807 601
rect 15833 575 15839 601
rect 17089 575 17095 601
rect 17121 575 17127 601
rect 18433 575 18439 601
rect 18465 575 18471 601
rect 19553 575 19559 601
rect 19585 575 19591 601
rect 20337 575 20343 601
rect 20369 575 20375 601
rect 21569 575 21575 601
rect 21601 575 21607 601
rect 22801 575 22807 601
rect 22833 575 22839 601
rect 23977 575 23983 601
rect 24009 575 24015 601
rect 24761 575 24767 601
rect 24793 575 24799 601
rect 25377 575 25383 601
rect 25409 575 25415 601
rect 26161 575 26167 601
rect 26193 575 26199 601
rect 29297 575 29303 601
rect 29329 575 29335 601
rect 31089 575 31095 601
rect 31121 575 31127 601
rect 13337 519 13343 545
rect 13369 519 13375 545
rect 17649 519 17655 545
rect 17681 519 17687 545
rect 21849 519 21855 545
rect 21881 519 21887 545
rect 23585 519 23591 545
rect 23617 519 23623 545
rect 24369 519 24375 545
rect 24401 519 24407 545
rect 26441 519 26447 545
rect 26473 519 26479 545
rect 30081 519 30087 545
rect 30113 519 30119 545
rect 16087 489 16113 495
rect 16087 457 16113 463
rect 17935 489 17961 495
rect 17935 457 17961 463
rect 18719 489 18745 495
rect 18719 457 18745 463
rect 19839 489 19865 495
rect 19839 457 19865 463
rect 20623 489 20649 495
rect 20623 457 20649 463
rect 25551 489 25577 495
rect 25551 457 25577 463
rect 336 405 31864 422
rect 336 379 2233 405
rect 2259 379 2285 405
rect 2311 379 2337 405
rect 2363 379 12233 405
rect 12259 379 12285 405
rect 12311 379 12337 405
rect 12363 379 22233 405
rect 22259 379 22285 405
rect 22311 379 22337 405
rect 22363 379 31864 405
rect 336 362 31864 379
<< via1 >>
rect 2233 6651 2259 6677
rect 2285 6651 2311 6677
rect 2337 6651 2363 6677
rect 12233 6651 12259 6677
rect 12285 6651 12311 6677
rect 12337 6651 12363 6677
rect 22233 6651 22259 6677
rect 22285 6651 22311 6677
rect 22337 6651 22363 6677
rect 1583 6567 1609 6593
rect 7519 6567 7545 6593
rect 9143 6567 9169 6593
rect 10599 6567 10625 6593
rect 12223 6567 12249 6593
rect 13231 6567 13257 6593
rect 31263 6567 31289 6593
rect 5111 6511 5137 6537
rect 6455 6511 6481 6537
rect 7239 6511 7265 6537
rect 1751 6455 1777 6481
rect 3655 6455 3681 6481
rect 6847 6455 6873 6481
rect 8863 6455 8889 6481
rect 10319 6455 10345 6481
rect 11943 6455 11969 6481
rect 12951 6455 12977 6481
rect 15303 6455 15329 6481
rect 16759 6455 16785 6481
rect 18271 6455 18297 6481
rect 21127 6455 21153 6481
rect 22583 6455 22609 6481
rect 24039 6455 24065 6481
rect 26895 6455 26921 6481
rect 28407 6455 28433 6481
rect 29751 6455 29777 6481
rect 30087 6455 30113 6481
rect 30983 6455 31009 6481
rect 3151 6399 3177 6425
rect 4607 6399 4633 6425
rect 14799 6399 14825 6425
rect 16255 6399 16281 6425
rect 17767 6399 17793 6425
rect 20623 6399 20649 6425
rect 22079 6399 22105 6425
rect 23535 6399 23561 6425
rect 26391 6399 26417 6425
rect 27903 6399 27929 6425
rect 29359 6399 29385 6425
rect 30591 6343 30617 6369
rect 1903 6259 1929 6285
rect 1955 6259 1981 6285
rect 2007 6259 2033 6285
rect 11903 6259 11929 6285
rect 11955 6259 11981 6285
rect 12007 6259 12033 6285
rect 21903 6259 21929 6285
rect 21955 6259 21981 6285
rect 22007 6259 22033 6285
rect 19167 6175 19193 6201
rect 24991 6175 25017 6201
rect 29527 6175 29553 6201
rect 6903 6119 6929 6145
rect 8527 6119 8553 6145
rect 30759 6119 30785 6145
rect 31543 6119 31569 6145
rect 7127 6063 7153 6089
rect 8751 6063 8777 6089
rect 17319 6063 17345 6089
rect 18607 6063 18633 6089
rect 20847 6063 20873 6089
rect 21127 6063 21153 6089
rect 30255 6063 30281 6089
rect 16759 6007 16785 6033
rect 17599 6007 17625 6033
rect 18887 6007 18913 6033
rect 19671 6007 19697 6033
rect 20679 6007 20705 6033
rect 25495 6007 25521 6033
rect 27567 6007 27593 6033
rect 29023 6007 29049 6033
rect 31039 6007 31065 6033
rect 16479 5951 16505 5977
rect 20399 5951 20425 5977
rect 27847 5951 27873 5977
rect 2233 5867 2259 5893
rect 2285 5867 2311 5893
rect 2337 5867 2363 5893
rect 12233 5867 12259 5893
rect 12285 5867 12311 5893
rect 12337 5867 12363 5893
rect 22233 5867 22259 5893
rect 22285 5867 22311 5893
rect 22337 5867 22363 5893
rect 9927 5727 9953 5753
rect 11047 5727 11073 5753
rect 12279 5727 12305 5753
rect 14967 5727 14993 5753
rect 16199 5727 16225 5753
rect 10207 5671 10233 5697
rect 11327 5671 11353 5697
rect 12559 5671 12585 5697
rect 12783 5671 12809 5697
rect 14687 5671 14713 5697
rect 16479 5671 16505 5697
rect 19447 5671 19473 5697
rect 21743 5671 21769 5697
rect 29359 5671 29385 5697
rect 30143 5671 30169 5697
rect 30927 5671 30953 5697
rect 13063 5615 13089 5641
rect 19727 5615 19753 5641
rect 22023 5615 22049 5641
rect 29863 5615 29889 5641
rect 30647 5615 30673 5641
rect 31375 5615 31401 5641
rect 1903 5475 1929 5501
rect 1955 5475 1981 5501
rect 2007 5475 2033 5501
rect 11903 5475 11929 5501
rect 11955 5475 11981 5501
rect 12007 5475 12033 5501
rect 21903 5475 21929 5501
rect 21955 5475 21981 5501
rect 22007 5475 22033 5501
rect 18719 5335 18745 5361
rect 18495 5279 18521 5305
rect 31095 5279 31121 5305
rect 15919 5223 15945 5249
rect 30255 5223 30281 5249
rect 30647 5223 30673 5249
rect 31431 5223 31457 5249
rect 15639 5167 15665 5193
rect 2233 5083 2259 5109
rect 2285 5083 2311 5109
rect 2337 5083 2363 5109
rect 12233 5083 12259 5109
rect 12285 5083 12311 5109
rect 12337 5083 12363 5109
rect 22233 5083 22259 5109
rect 22285 5083 22311 5109
rect 22337 5083 22363 5109
rect 16535 4999 16561 5025
rect 12783 4943 12809 4969
rect 18719 4943 18745 4969
rect 30535 4943 30561 4969
rect 4159 4887 4185 4913
rect 12503 4887 12529 4913
rect 18495 4887 18521 4913
rect 30143 4887 30169 4913
rect 30927 4887 30953 4913
rect 3935 4831 3961 4857
rect 16759 4831 16785 4857
rect 31375 4831 31401 4857
rect 1903 4691 1929 4717
rect 1955 4691 1981 4717
rect 2007 4691 2033 4717
rect 11903 4691 11929 4717
rect 11955 4691 11981 4717
rect 12007 4691 12033 4717
rect 21903 4691 21929 4717
rect 21955 4691 21981 4717
rect 22007 4691 22033 4717
rect 30759 4607 30785 4633
rect 14519 4551 14545 4577
rect 20287 4551 20313 4577
rect 11663 4495 11689 4521
rect 14295 4495 14321 4521
rect 17263 4495 17289 4521
rect 30255 4495 30281 4521
rect 31095 4495 31121 4521
rect 967 4439 993 4465
rect 11943 4439 11969 4465
rect 31431 4439 31457 4465
rect 1247 4383 1273 4409
rect 16983 4383 17009 4409
rect 20007 4383 20033 4409
rect 2233 4299 2259 4325
rect 2285 4299 2311 4325
rect 2337 4299 2363 4325
rect 12233 4299 12259 4325
rect 12285 4299 12311 4325
rect 12337 4299 12363 4325
rect 22233 4299 22259 4325
rect 22285 4299 22311 4325
rect 22337 4299 22363 4325
rect 18887 4215 18913 4241
rect 19167 4159 19193 4185
rect 30479 4103 30505 4129
rect 30927 4103 30953 4129
rect 30703 4047 30729 4073
rect 31431 3991 31457 4017
rect 1903 3907 1929 3933
rect 1955 3907 1981 3933
rect 2007 3907 2033 3933
rect 11903 3907 11929 3933
rect 11955 3907 11981 3933
rect 12007 3907 12033 3933
rect 21903 3907 21929 3933
rect 21955 3907 21981 3933
rect 22007 3907 22033 3933
rect 31543 3823 31569 3849
rect 6119 3767 6145 3793
rect 13063 3767 13089 3793
rect 17487 3767 17513 3793
rect 30759 3767 30785 3793
rect 4439 3711 4465 3737
rect 5895 3711 5921 3737
rect 12783 3711 12809 3737
rect 13679 3711 13705 3737
rect 14743 3711 14769 3737
rect 15023 3711 15049 3737
rect 17767 3711 17793 3737
rect 20567 3711 20593 3737
rect 29415 3711 29441 3737
rect 31095 3711 31121 3737
rect 10039 3655 10065 3681
rect 10431 3655 10457 3681
rect 13959 3655 13985 3681
rect 18495 3655 18521 3681
rect 20847 3655 20873 3681
rect 29639 3655 29665 3681
rect 30255 3655 30281 3681
rect 4719 3599 4745 3625
rect 9759 3599 9785 3625
rect 10711 3599 10737 3625
rect 18215 3599 18241 3625
rect 2233 3515 2259 3541
rect 2285 3515 2311 3541
rect 2337 3515 2363 3541
rect 12233 3515 12259 3541
rect 12285 3515 12311 3541
rect 12337 3515 12363 3541
rect 22233 3515 22259 3541
rect 22285 3515 22311 3541
rect 22337 3515 22363 3541
rect 15639 3375 15665 3401
rect 2647 3319 2673 3345
rect 6455 3319 6481 3345
rect 6679 3319 6705 3345
rect 15359 3319 15385 3345
rect 24487 3319 24513 3345
rect 30143 3319 30169 3345
rect 30927 3319 30953 3345
rect 2423 3263 2449 3289
rect 24711 3263 24737 3289
rect 31431 3263 31457 3289
rect 30647 3207 30673 3233
rect 1903 3123 1929 3149
rect 1955 3123 1981 3149
rect 2007 3123 2033 3149
rect 11903 3123 11929 3149
rect 11955 3123 11981 3149
rect 12007 3123 12033 3149
rect 21903 3123 21929 3149
rect 21955 3123 21981 3149
rect 22007 3123 22033 3149
rect 31543 3039 31569 3065
rect 20679 2983 20705 3009
rect 30815 2983 30841 3009
rect 17543 2927 17569 2953
rect 20399 2927 20425 2953
rect 22527 2927 22553 2953
rect 23423 2927 23449 2953
rect 25439 2927 25465 2953
rect 31095 2927 31121 2953
rect 17823 2871 17849 2897
rect 22807 2871 22833 2897
rect 23703 2871 23729 2897
rect 25719 2871 25745 2897
rect 27063 2871 27089 2897
rect 26783 2815 26809 2841
rect 30591 2815 30617 2841
rect 2233 2731 2259 2757
rect 2285 2731 2311 2757
rect 2337 2731 2363 2757
rect 12233 2731 12259 2757
rect 12285 2731 12311 2757
rect 12337 2731 12363 2757
rect 22233 2731 22259 2757
rect 22285 2731 22311 2757
rect 22337 2731 22363 2757
rect 11327 2647 11353 2673
rect 13119 2647 13145 2673
rect 16983 2647 17009 2673
rect 22191 2647 22217 2673
rect 27399 2647 27425 2673
rect 911 2591 937 2617
rect 4439 2591 4465 2617
rect 10319 2591 10345 2617
rect 10599 2591 10625 2617
rect 13399 2591 13425 2617
rect 19167 2591 19193 2617
rect 19447 2591 19473 2617
rect 21631 2591 21657 2617
rect 30143 2591 30169 2617
rect 30927 2591 30953 2617
rect 31319 2591 31345 2617
rect 1191 2535 1217 2561
rect 4719 2535 4745 2561
rect 11047 2535 11073 2561
rect 21799 2535 21825 2561
rect 22471 2535 22497 2561
rect 27679 2535 27705 2561
rect 30535 2535 30561 2561
rect 10767 2479 10793 2505
rect 11607 2479 11633 2505
rect 17207 2479 17233 2505
rect 1903 2339 1929 2365
rect 1955 2339 1981 2365
rect 2007 2339 2033 2365
rect 11903 2339 11929 2365
rect 11955 2339 11981 2365
rect 12007 2339 12033 2365
rect 21903 2339 21929 2365
rect 21955 2339 21981 2365
rect 22007 2339 22033 2365
rect 31543 2255 31569 2281
rect 7687 2199 7713 2225
rect 9199 2199 9225 2225
rect 11719 2199 11745 2225
rect 13903 2199 13929 2225
rect 21743 2199 21769 2225
rect 23591 2199 23617 2225
rect 24095 2199 24121 2225
rect 29583 2199 29609 2225
rect 16479 2143 16505 2169
rect 18831 2143 18857 2169
rect 21519 2143 21545 2169
rect 24319 2143 24345 2169
rect 25103 2143 25129 2169
rect 29415 2143 29441 2169
rect 30255 2143 30281 2169
rect 31095 2143 31121 2169
rect 11495 2087 11521 2113
rect 12895 2087 12921 2113
rect 15975 2087 16001 2113
rect 16255 2087 16281 2113
rect 16759 2087 16785 2113
rect 19111 2087 19137 2113
rect 20455 2087 20481 2113
rect 21071 2087 21097 2113
rect 23927 2087 23953 2113
rect 30647 2087 30673 2113
rect 7911 2031 7937 2057
rect 8975 2031 9001 2057
rect 12615 2031 12641 2057
rect 13679 2031 13705 2057
rect 20175 2031 20201 2057
rect 20791 2031 20817 2057
rect 25383 2031 25409 2057
rect 2233 1947 2259 1973
rect 2285 1947 2311 1973
rect 2337 1947 2363 1973
rect 12233 1947 12259 1973
rect 12285 1947 12311 1973
rect 12337 1947 12363 1973
rect 22233 1947 22259 1973
rect 22285 1947 22311 1973
rect 22337 1947 22363 1973
rect 15639 1863 15665 1889
rect 16199 1863 16225 1889
rect 17935 1863 17961 1889
rect 6007 1807 6033 1833
rect 13959 1807 13985 1833
rect 14127 1807 14153 1833
rect 15919 1807 15945 1833
rect 16479 1807 16505 1833
rect 18383 1807 18409 1833
rect 20735 1807 20761 1833
rect 23087 1807 23113 1833
rect 24039 1807 24065 1833
rect 24823 1807 24849 1833
rect 25607 1807 25633 1833
rect 27959 1807 27985 1833
rect 28463 1807 28489 1833
rect 30143 1807 30169 1833
rect 30927 1807 30953 1833
rect 6287 1751 6313 1777
rect 7015 1751 7041 1777
rect 13735 1751 13761 1777
rect 15191 1751 15217 1777
rect 19167 1751 19193 1777
rect 21463 1751 21489 1777
rect 22303 1751 22329 1777
rect 25887 1751 25913 1777
rect 28239 1751 28265 1777
rect 28743 1751 28769 1777
rect 7295 1695 7321 1721
rect 15471 1695 15497 1721
rect 18215 1695 18241 1721
rect 19447 1695 19473 1721
rect 20231 1695 20257 1721
rect 21015 1695 21041 1721
rect 21799 1695 21825 1721
rect 22751 1695 22777 1721
rect 24375 1695 24401 1721
rect 25271 1695 25297 1721
rect 30647 1695 30673 1721
rect 31431 1695 31457 1721
rect 14407 1639 14433 1665
rect 18663 1639 18689 1665
rect 1903 1555 1929 1581
rect 1955 1555 1981 1581
rect 2007 1555 2033 1581
rect 11903 1555 11929 1581
rect 11955 1555 11981 1581
rect 12007 1555 12033 1581
rect 21903 1555 21929 1581
rect 21955 1555 21981 1581
rect 22007 1555 22033 1581
rect 31543 1471 31569 1497
rect 22975 1415 23001 1441
rect 26111 1415 26137 1441
rect 26727 1415 26753 1441
rect 14351 1359 14377 1385
rect 15975 1359 16001 1385
rect 16815 1359 16841 1385
rect 17263 1359 17289 1385
rect 18159 1359 18185 1385
rect 18943 1359 18969 1385
rect 19727 1359 19753 1385
rect 20511 1359 20537 1385
rect 22583 1359 22609 1385
rect 23479 1359 23505 1385
rect 24487 1359 24513 1385
rect 25215 1359 25241 1385
rect 30255 1359 30281 1385
rect 31095 1359 31121 1385
rect 911 1303 937 1329
rect 13959 1303 13985 1329
rect 15135 1303 15161 1329
rect 17039 1303 17065 1329
rect 17655 1303 17681 1329
rect 18551 1303 18577 1329
rect 21295 1303 21321 1329
rect 21575 1303 21601 1329
rect 22303 1303 22329 1329
rect 23647 1303 23673 1329
rect 29359 1303 29385 1329
rect 30647 1303 30673 1329
rect 1191 1247 1217 1273
rect 13679 1247 13705 1273
rect 14631 1247 14657 1273
rect 15415 1247 15441 1273
rect 16199 1247 16225 1273
rect 19223 1247 19249 1273
rect 20007 1247 20033 1273
rect 20791 1247 20817 1273
rect 23927 1247 23953 1273
rect 24711 1247 24737 1273
rect 25495 1247 25521 1273
rect 26391 1247 26417 1273
rect 27007 1247 27033 1273
rect 29639 1247 29665 1273
rect 2233 1163 2259 1189
rect 2285 1163 2311 1189
rect 2337 1163 2363 1189
rect 12233 1163 12259 1189
rect 12285 1163 12311 1189
rect 12337 1163 12363 1189
rect 22233 1163 22259 1189
rect 22285 1163 22311 1189
rect 22337 1163 22363 1189
rect 10543 1079 10569 1105
rect 12839 1079 12865 1105
rect 13287 1079 13313 1105
rect 21183 1079 21209 1105
rect 29639 1079 29665 1105
rect 2367 1023 2393 1049
rect 10823 1023 10849 1049
rect 14519 1023 14545 1049
rect 16367 1023 16393 1049
rect 17151 1023 17177 1049
rect 17935 1023 17961 1049
rect 18719 1023 18745 1049
rect 20903 1023 20929 1049
rect 23087 1023 23113 1049
rect 23255 1023 23281 1049
rect 29191 1023 29217 1049
rect 29919 1023 29945 1049
rect 30927 1023 30953 1049
rect 1191 967 1217 993
rect 2647 967 2673 993
rect 10375 967 10401 993
rect 12615 967 12641 993
rect 13735 967 13761 993
rect 15415 967 15441 993
rect 19503 967 19529 993
rect 19783 967 19809 993
rect 20119 967 20145 993
rect 21743 967 21769 993
rect 23479 967 23505 993
rect 24039 967 24065 993
rect 24879 967 24905 993
rect 25719 967 25745 993
rect 26447 967 26473 993
rect 29471 967 29497 993
rect 30143 967 30169 993
rect 967 911 993 937
rect 10151 911 10177 937
rect 12391 911 12417 937
rect 13119 911 13145 937
rect 13567 911 13593 937
rect 14911 911 14937 937
rect 18215 911 18241 937
rect 22695 911 22721 937
rect 24431 911 24457 937
rect 25215 911 25241 937
rect 25887 911 25913 937
rect 31431 911 31457 937
rect 14239 855 14265 881
rect 15583 855 15609 881
rect 16647 855 16673 881
rect 17431 855 17457 881
rect 18999 855 19025 881
rect 20399 855 20425 881
rect 21967 855 21993 881
rect 26671 855 26697 881
rect 30647 855 30673 881
rect 1903 771 1929 797
rect 1955 771 1981 797
rect 2007 771 2033 797
rect 11903 771 11929 797
rect 11955 771 11981 797
rect 12007 771 12033 797
rect 21903 771 21929 797
rect 21955 771 21981 797
rect 22007 771 22033 797
rect 31543 687 31569 713
rect 14575 631 14601 657
rect 15359 631 15385 657
rect 16703 631 16729 657
rect 22359 631 22385 657
rect 29807 631 29833 657
rect 30591 631 30617 657
rect 12951 575 12977 601
rect 14071 575 14097 601
rect 14855 575 14881 601
rect 15807 575 15833 601
rect 17095 575 17121 601
rect 18439 575 18465 601
rect 19559 575 19585 601
rect 20343 575 20369 601
rect 21575 575 21601 601
rect 22807 575 22833 601
rect 23983 575 24009 601
rect 24767 575 24793 601
rect 25383 575 25409 601
rect 26167 575 26193 601
rect 29303 575 29329 601
rect 31095 575 31121 601
rect 13343 519 13369 545
rect 17655 519 17681 545
rect 21855 519 21881 545
rect 23591 519 23617 545
rect 24375 519 24401 545
rect 26447 519 26473 545
rect 30087 519 30113 545
rect 16087 463 16113 489
rect 17935 463 17961 489
rect 18719 463 18745 489
rect 19839 463 19865 489
rect 20623 463 20649 489
rect 25551 463 25577 489
rect 2233 379 2259 405
rect 2285 379 2311 405
rect 2337 379 2363 405
rect 12233 379 12259 405
rect 12285 379 12311 405
rect 12337 379 12363 405
rect 22233 379 22259 405
rect 22285 379 22311 405
rect 22337 379 22363 405
<< metal2 >>
rect 1456 7056 1512 7112
rect 2912 7056 2968 7112
rect 4368 7056 4424 7112
rect 5824 7056 5880 7112
rect 7280 7056 7336 7112
rect 8736 7056 8792 7112
rect 10192 7056 10248 7112
rect 11648 7056 11704 7112
rect 13104 7056 13160 7112
rect 14560 7056 14616 7112
rect 16016 7056 16072 7112
rect 17472 7056 17528 7112
rect 18928 7056 18984 7112
rect 20384 7056 20440 7112
rect 21840 7056 21896 7112
rect 23296 7056 23352 7112
rect 24752 7056 24808 7112
rect 26208 7056 26264 7112
rect 27664 7056 27720 7112
rect 29120 7056 29176 7112
rect 30576 7056 30632 7112
rect 910 6986 938 6991
rect 798 6762 826 6767
rect 798 5698 826 6734
rect 910 5810 938 6958
rect 1470 6818 1498 7056
rect 2926 7042 2954 7056
rect 2926 7009 2954 7014
rect 3150 7042 3178 7047
rect 1470 6790 1610 6818
rect 1582 6593 1610 6790
rect 2232 6678 2364 6683
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2232 6645 2364 6650
rect 1582 6567 1583 6593
rect 1609 6567 1610 6593
rect 1582 6561 1610 6567
rect 1750 6482 1778 6487
rect 1750 6435 1778 6454
rect 3150 6425 3178 7014
rect 4382 7042 4410 7056
rect 4382 7009 4410 7014
rect 4606 7042 4634 7047
rect 3822 6762 3850 6767
rect 3150 6399 3151 6425
rect 3177 6399 3178 6425
rect 3150 6393 3178 6399
rect 3654 6481 3682 6487
rect 3654 6455 3655 6481
rect 3681 6455 3682 6481
rect 3654 6370 3682 6455
rect 3654 6337 3682 6342
rect 1902 6286 2034 6291
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 1902 6253 2034 6258
rect 2232 5894 2364 5899
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2232 5861 2364 5866
rect 910 5777 938 5782
rect 798 5665 826 5670
rect 1902 5502 2034 5507
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 1902 5469 2034 5474
rect 2814 5306 2842 5311
rect 2232 5110 2364 5115
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2232 5077 2364 5082
rect 1902 4718 2034 4723
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 1902 4685 2034 4690
rect 966 4466 994 4471
rect 966 4419 994 4438
rect 1246 4410 1274 4415
rect 1246 4363 1274 4382
rect 2232 4326 2364 4331
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2232 4293 2364 4298
rect 1526 4018 1554 4023
rect 350 3066 378 3071
rect 350 1386 378 3038
rect 1526 2730 1554 3990
rect 1902 3934 2034 3939
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 1902 3901 2034 3906
rect 1526 2697 1554 2702
rect 1638 3794 1666 3799
rect 910 2618 938 2623
rect 910 2571 938 2590
rect 1190 2562 1218 2567
rect 1190 2515 1218 2534
rect 1022 2170 1050 2175
rect 350 1353 378 1358
rect 854 1778 882 1783
rect 854 938 882 1750
rect 910 1330 938 1335
rect 910 1283 938 1302
rect 854 905 882 910
rect 966 938 994 943
rect 966 891 994 910
rect 1022 882 1050 2142
rect 1190 1274 1218 1279
rect 1190 1227 1218 1246
rect 1638 1162 1666 3766
rect 2232 3542 2364 3547
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2232 3509 2364 3514
rect 2646 3345 2674 3351
rect 2646 3319 2647 3345
rect 2673 3319 2674 3345
rect 2422 3289 2450 3295
rect 2422 3263 2423 3289
rect 2449 3263 2450 3289
rect 1902 3150 2034 3155
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 1902 3117 2034 3122
rect 2422 2842 2450 3263
rect 2646 2898 2674 3319
rect 2646 2865 2674 2870
rect 2422 2809 2450 2814
rect 2232 2758 2364 2763
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2232 2725 2364 2730
rect 2534 2450 2562 2455
rect 1902 2366 2034 2371
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 1902 2333 2034 2338
rect 2086 2114 2114 2119
rect 1902 1582 2034 1587
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 1902 1549 2034 1554
rect 1638 1129 1666 1134
rect 1022 849 1050 854
rect 1190 993 1218 999
rect 1190 967 1191 993
rect 1217 967 1218 993
rect 1190 154 1218 967
rect 1902 798 2034 803
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 1902 765 2034 770
rect 2086 490 2114 2086
rect 2232 1974 2364 1979
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2232 1941 2364 1946
rect 2534 1498 2562 2422
rect 2814 2058 2842 5278
rect 2814 2025 2842 2030
rect 2926 3570 2954 3575
rect 2534 1465 2562 1470
rect 2534 1386 2562 1391
rect 2232 1190 2364 1195
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2232 1157 2364 1162
rect 2366 1106 2394 1111
rect 2366 1049 2394 1078
rect 2366 1023 2367 1049
rect 2393 1023 2394 1049
rect 2366 1017 2394 1023
rect 2086 457 2114 462
rect 2232 406 2364 411
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2232 373 2364 378
rect 2366 322 2394 327
rect 1190 121 1218 126
rect 2142 210 2170 215
rect 2142 56 2170 182
rect 2366 56 2394 294
rect 2534 266 2562 1358
rect 2646 993 2674 999
rect 2646 967 2647 993
rect 2673 967 2674 993
rect 2534 233 2562 238
rect 2590 826 2618 831
rect 2590 56 2618 798
rect 2646 602 2674 967
rect 2646 569 2674 574
rect 2926 322 2954 3542
rect 3822 2450 3850 6734
rect 4606 6425 4634 7014
rect 5110 6874 5138 6879
rect 5110 6537 5138 6846
rect 5110 6511 5111 6537
rect 5137 6511 5138 6537
rect 5110 6505 5138 6511
rect 5838 6538 5866 7056
rect 7294 7042 7322 7056
rect 7294 7009 7322 7014
rect 7518 7042 7546 7047
rect 6734 6650 6762 6655
rect 5838 6505 5866 6510
rect 6454 6538 6482 6543
rect 6454 6491 6482 6510
rect 4606 6399 4607 6425
rect 4633 6399 4634 6425
rect 4606 6393 4634 6399
rect 5838 6202 5866 6207
rect 5446 5922 5474 5927
rect 4214 5138 4242 5143
rect 4158 4914 4186 4919
rect 4158 4867 4186 4886
rect 3934 4858 3962 4863
rect 3934 4811 3962 4830
rect 4214 4018 4242 5110
rect 4214 3985 4242 3990
rect 4270 4746 4298 4751
rect 3822 2417 3850 2422
rect 3934 3346 3962 3351
rect 3486 1890 3514 1895
rect 3262 1554 3290 1559
rect 2926 289 2954 294
rect 3038 322 3066 327
rect 2814 266 2842 271
rect 2814 56 2842 238
rect 3038 56 3066 294
rect 3262 56 3290 1526
rect 3486 56 3514 1862
rect 3710 1834 3738 1839
rect 3710 56 3738 1806
rect 3934 56 3962 3318
rect 4270 3066 4298 4718
rect 4438 3738 4466 3743
rect 4438 3691 4466 3710
rect 4718 3625 4746 3631
rect 4718 3599 4719 3625
rect 4745 3599 4746 3625
rect 4718 3514 4746 3599
rect 4718 3481 4746 3486
rect 4830 3402 4858 3407
rect 4270 3033 4298 3038
rect 4606 3122 4634 3127
rect 4438 2618 4466 2623
rect 4438 2571 4466 2590
rect 4158 2058 4186 2063
rect 4158 56 4186 2030
rect 4382 1162 4410 1167
rect 4382 56 4410 1134
rect 4606 56 4634 3094
rect 4718 2561 4746 2567
rect 4718 2535 4719 2561
rect 4745 2535 4746 2561
rect 4718 210 4746 2535
rect 4718 177 4746 182
rect 4830 56 4858 3374
rect 5278 2674 5306 2679
rect 4998 2562 5026 2567
rect 4998 1218 5026 2534
rect 4998 1185 5026 1190
rect 5054 770 5082 775
rect 5054 56 5082 742
rect 5278 56 5306 2646
rect 5446 2282 5474 5894
rect 5838 5810 5866 6174
rect 5838 5777 5866 5782
rect 6510 6146 6538 6151
rect 6118 3906 6146 3911
rect 6118 3793 6146 3878
rect 6118 3767 6119 3793
rect 6145 3767 6146 3793
rect 6118 3761 6146 3767
rect 5446 2249 5474 2254
rect 5894 3737 5922 3743
rect 5894 3711 5895 3737
rect 5921 3711 5922 3737
rect 5726 2002 5754 2007
rect 5502 434 5530 439
rect 5502 56 5530 406
rect 5726 56 5754 1974
rect 5894 1722 5922 3711
rect 6454 3346 6482 3351
rect 6454 3299 6482 3318
rect 6454 2954 6482 2959
rect 6006 2506 6034 2511
rect 5838 1694 5922 1722
rect 5950 2226 5978 2231
rect 5838 826 5866 1694
rect 5838 793 5866 798
rect 5950 56 5978 2198
rect 6006 1833 6034 2478
rect 6454 2282 6482 2926
rect 6454 2249 6482 2254
rect 6006 1807 6007 1833
rect 6033 1807 6034 1833
rect 6006 1801 6034 1807
rect 6286 1777 6314 1783
rect 6286 1751 6287 1777
rect 6313 1751 6314 1777
rect 6286 770 6314 1751
rect 6510 1666 6538 6118
rect 6678 5026 6706 5031
rect 6510 1633 6538 1638
rect 6622 3962 6650 3967
rect 6286 737 6314 742
rect 6398 938 6426 943
rect 6174 714 6202 719
rect 6174 56 6202 686
rect 6398 56 6426 910
rect 6622 56 6650 3934
rect 6678 3458 6706 4998
rect 6734 4802 6762 6622
rect 7014 6594 7042 6599
rect 6902 6538 6930 6543
rect 6846 6481 6874 6487
rect 6846 6455 6847 6481
rect 6873 6455 6874 6481
rect 6846 6426 6874 6455
rect 6846 6393 6874 6398
rect 6790 6314 6818 6319
rect 6790 5866 6818 6286
rect 6902 6145 6930 6510
rect 6902 6119 6903 6145
rect 6929 6119 6930 6145
rect 6902 6113 6930 6119
rect 6790 5833 6818 5838
rect 6734 4769 6762 4774
rect 7014 4298 7042 6566
rect 7294 6594 7322 6599
rect 7238 6538 7266 6543
rect 7238 6491 7266 6510
rect 7294 6258 7322 6566
rect 7518 6593 7546 7014
rect 8750 7042 8778 7056
rect 8750 7009 8778 7014
rect 9142 7042 9170 7047
rect 7518 6567 7519 6593
rect 7545 6567 7546 6593
rect 7518 6561 7546 6567
rect 7742 6706 7770 6711
rect 7126 6230 7322 6258
rect 7350 6538 7378 6543
rect 7126 6089 7154 6230
rect 7126 6063 7127 6089
rect 7153 6063 7154 6089
rect 7126 6057 7154 6063
rect 7238 5586 7266 5591
rect 7238 4970 7266 5558
rect 7238 4937 7266 4942
rect 7350 4634 7378 6510
rect 7462 6482 7490 6487
rect 7462 5026 7490 6454
rect 7462 4993 7490 4998
rect 7686 5138 7714 5143
rect 7686 4970 7714 5110
rect 7686 4937 7714 4942
rect 7238 4606 7378 4634
rect 7406 4802 7434 4807
rect 7014 4265 7042 4270
rect 7126 4466 7154 4471
rect 6846 3794 6874 3799
rect 6678 3425 6706 3430
rect 6734 3682 6762 3687
rect 6678 3345 6706 3351
rect 6678 3319 6679 3345
rect 6705 3319 6706 3345
rect 6678 3290 6706 3319
rect 6678 3257 6706 3262
rect 6734 3066 6762 3654
rect 6734 3033 6762 3038
rect 6734 2898 6762 2903
rect 6734 2170 6762 2870
rect 6734 2137 6762 2142
rect 6790 1274 6818 1279
rect 6678 1050 6706 1055
rect 6678 546 6706 1022
rect 6790 658 6818 1246
rect 6846 826 6874 3766
rect 7070 2786 7098 2791
rect 7014 1777 7042 1783
rect 7014 1751 7015 1777
rect 7041 1751 7042 1777
rect 6846 793 6874 798
rect 6958 1442 6986 1447
rect 6790 625 6818 630
rect 6678 513 6706 518
rect 6846 490 6874 495
rect 6846 56 6874 462
rect 6958 378 6986 1414
rect 6958 345 6986 350
rect 7014 266 7042 1751
rect 7070 1330 7098 2758
rect 7126 2730 7154 4438
rect 7238 3850 7266 4606
rect 7238 3817 7266 3822
rect 7350 4354 7378 4359
rect 7126 2697 7154 2702
rect 7238 3234 7266 3239
rect 7126 1722 7154 1727
rect 7126 1386 7154 1694
rect 7126 1353 7154 1358
rect 7182 1610 7210 1615
rect 7070 1297 7098 1302
rect 7014 233 7042 238
rect 7070 826 7098 831
rect 7070 56 7098 798
rect 7182 322 7210 1582
rect 7238 1386 7266 3206
rect 7350 2730 7378 4326
rect 7350 2697 7378 2702
rect 7406 2674 7434 4774
rect 7462 4634 7490 4639
rect 7490 4606 7546 4634
rect 7462 4601 7490 4606
rect 7462 4466 7490 4471
rect 7462 4354 7490 4438
rect 7462 4321 7490 4326
rect 7462 4242 7490 4247
rect 7462 3626 7490 4214
rect 7518 4130 7546 4606
rect 7518 4097 7546 4102
rect 7574 4466 7602 4471
rect 7518 3850 7546 3855
rect 7518 3738 7546 3822
rect 7518 3705 7546 3710
rect 7462 3593 7490 3598
rect 7574 3402 7602 4438
rect 7406 2641 7434 2646
rect 7518 3374 7602 3402
rect 7686 3402 7714 3407
rect 7518 2618 7546 3374
rect 7518 2585 7546 2590
rect 7406 2394 7434 2399
rect 7238 1353 7266 1358
rect 7294 1721 7322 1727
rect 7294 1695 7295 1721
rect 7321 1695 7322 1721
rect 7294 546 7322 1695
rect 7350 1274 7378 1279
rect 7350 714 7378 1246
rect 7350 681 7378 686
rect 7294 513 7322 518
rect 7406 434 7434 2366
rect 7686 2225 7714 3374
rect 7686 2199 7687 2225
rect 7713 2199 7714 2225
rect 7686 2193 7714 2199
rect 7406 401 7434 406
rect 7462 1218 7490 1223
rect 7182 289 7210 294
rect 7294 378 7322 383
rect 7294 56 7322 350
rect 7462 322 7490 1190
rect 7462 289 7490 294
rect 7518 882 7546 887
rect 7518 56 7546 854
rect 7742 56 7770 6678
rect 9142 6593 9170 7014
rect 10206 7042 10234 7056
rect 10206 7009 10234 7014
rect 10598 7042 10626 7047
rect 9142 6567 9143 6593
rect 9169 6567 9170 6593
rect 9142 6561 9170 6567
rect 10262 6650 10290 6655
rect 8862 6482 8890 6487
rect 8526 6481 8890 6482
rect 8526 6455 8863 6481
rect 8889 6455 8890 6481
rect 8526 6454 8890 6455
rect 8526 6145 8554 6454
rect 8862 6449 8890 6454
rect 9926 6482 9954 6487
rect 8526 6119 8527 6145
rect 8553 6119 8554 6145
rect 8526 6113 8554 6119
rect 8750 6202 8778 6207
rect 8358 6090 8386 6095
rect 8246 5754 8274 5759
rect 8022 4522 8050 4527
rect 7910 2057 7938 2063
rect 7910 2031 7911 2057
rect 7937 2031 7938 2057
rect 7910 1778 7938 2031
rect 7910 1745 7938 1750
rect 8022 826 8050 4494
rect 8246 3346 8274 5726
rect 8246 3313 8274 3318
rect 8302 4858 8330 4863
rect 8078 3066 8106 3071
rect 8078 994 8106 3038
rect 8302 1106 8330 4830
rect 8358 4746 8386 6062
rect 8750 6089 8778 6174
rect 8750 6063 8751 6089
rect 8777 6063 8778 6089
rect 8750 6057 8778 6063
rect 9926 5753 9954 6454
rect 9926 5727 9927 5753
rect 9953 5727 9954 5753
rect 9926 5721 9954 5727
rect 10206 5697 10234 5703
rect 10206 5671 10207 5697
rect 10233 5671 10234 5697
rect 9086 5362 9114 5367
rect 9086 4914 9114 5334
rect 10038 5194 10066 5199
rect 9086 4881 9114 4886
rect 9982 5082 10010 5087
rect 8358 4713 8386 4718
rect 8862 4746 8890 4751
rect 8358 4634 8386 4639
rect 8358 3682 8386 4606
rect 8862 4242 8890 4718
rect 8862 4209 8890 4214
rect 9982 3962 10010 5054
rect 10038 4242 10066 5166
rect 10206 5082 10234 5671
rect 10206 5049 10234 5054
rect 10038 4209 10066 4214
rect 9982 3929 10010 3934
rect 8358 3649 8386 3654
rect 10038 3681 10066 3687
rect 10038 3655 10039 3681
rect 10065 3655 10066 3681
rect 9758 3625 9786 3631
rect 9758 3599 9759 3625
rect 9785 3599 9786 3625
rect 9758 3570 9786 3599
rect 9758 3537 9786 3542
rect 9198 3514 9226 3519
rect 9226 3486 9282 3514
rect 9198 3481 9226 3486
rect 8862 3234 8890 3239
rect 8470 2226 8498 2231
rect 8302 1073 8330 1078
rect 8414 1946 8442 1951
rect 8078 961 8106 966
rect 8190 994 8218 999
rect 8022 793 8050 798
rect 7966 714 7994 719
rect 7966 56 7994 686
rect 8190 56 8218 966
rect 8414 826 8442 1918
rect 8414 793 8442 798
rect 8470 154 8498 2198
rect 8414 126 8498 154
rect 8638 154 8666 159
rect 8414 56 8442 126
rect 8638 56 8666 126
rect 8862 56 8890 3206
rect 9086 2618 9114 2623
rect 8974 2058 9002 2063
rect 8974 2011 9002 2030
rect 9086 1442 9114 2590
rect 9198 2225 9226 2231
rect 9198 2199 9199 2225
rect 9225 2199 9226 2225
rect 9086 1409 9114 1414
rect 9142 1946 9170 1951
rect 9142 994 9170 1918
rect 9198 1330 9226 2199
rect 9254 1694 9282 3486
rect 9870 3458 9898 3463
rect 9870 2842 9898 3430
rect 9870 2809 9898 2814
rect 9926 2954 9954 2959
rect 9758 2730 9786 2735
rect 9254 1666 9450 1694
rect 9198 1297 9226 1302
rect 9142 961 9170 966
rect 9310 658 9338 663
rect 9086 434 9114 439
rect 9086 56 9114 406
rect 9310 56 9338 630
rect 9422 658 9450 1666
rect 9422 625 9450 630
rect 9534 322 9562 327
rect 9534 56 9562 294
rect 9758 56 9786 2702
rect 9926 1106 9954 2926
rect 9982 2282 10010 2287
rect 9982 1218 10010 2254
rect 9982 1185 10010 1190
rect 9926 1078 10010 1106
rect 9982 56 10010 1078
rect 10038 994 10066 3655
rect 10262 3346 10290 6622
rect 10598 6593 10626 7014
rect 10598 6567 10599 6593
rect 10625 6567 10626 6593
rect 10598 6561 10626 6567
rect 10990 6930 11018 6935
rect 10318 6482 10346 6487
rect 10318 6435 10346 6454
rect 10598 6370 10626 6375
rect 10598 5586 10626 6342
rect 10598 5553 10626 5558
rect 10934 5698 10962 5703
rect 10934 5474 10962 5670
rect 10934 5441 10962 5446
rect 10318 4578 10346 4583
rect 10318 3906 10346 4550
rect 10430 4578 10458 4583
rect 10430 4466 10458 4550
rect 10654 4522 10682 4527
rect 10430 4433 10458 4438
rect 10542 4466 10570 4471
rect 10542 4018 10570 4438
rect 10654 4354 10682 4494
rect 10654 4321 10682 4326
rect 10934 4522 10962 4527
rect 10598 4298 10626 4303
rect 10598 4074 10626 4270
rect 10822 4186 10850 4191
rect 10934 4186 10962 4494
rect 10850 4158 10962 4186
rect 10822 4153 10850 4158
rect 10598 4041 10626 4046
rect 10542 3985 10570 3990
rect 10598 3906 10626 3911
rect 10318 3878 10570 3906
rect 10430 3681 10458 3687
rect 10430 3655 10431 3681
rect 10457 3655 10458 3681
rect 10430 3626 10458 3655
rect 10430 3593 10458 3598
rect 10262 3313 10290 3318
rect 10374 2954 10402 2959
rect 10318 2618 10346 2623
rect 10318 2571 10346 2590
rect 10374 2226 10402 2926
rect 10486 2786 10514 2791
rect 10374 2193 10402 2198
rect 10430 2282 10458 2287
rect 10038 961 10066 966
rect 10374 993 10402 999
rect 10374 967 10375 993
rect 10401 967 10402 993
rect 10150 937 10178 943
rect 10150 911 10151 937
rect 10177 911 10178 937
rect 10094 714 10122 719
rect 10150 714 10178 911
rect 10206 714 10234 719
rect 10150 686 10206 714
rect 10094 322 10122 686
rect 10206 681 10234 686
rect 10094 289 10122 294
rect 10206 602 10234 607
rect 10206 56 10234 574
rect 10374 490 10402 967
rect 10374 457 10402 462
rect 10430 434 10458 2254
rect 10486 2226 10514 2758
rect 10486 2193 10514 2198
rect 10542 1386 10570 3878
rect 10598 3738 10626 3878
rect 10598 3705 10626 3710
rect 10654 3850 10682 3855
rect 10598 2842 10626 2847
rect 10598 2617 10626 2814
rect 10598 2591 10599 2617
rect 10625 2591 10626 2617
rect 10598 2585 10626 2591
rect 10654 2338 10682 3822
rect 10710 3625 10738 3631
rect 10710 3599 10711 3625
rect 10737 3599 10738 3625
rect 10710 3402 10738 3599
rect 10990 3570 11018 6902
rect 11662 6538 11690 7056
rect 12614 6818 12642 6823
rect 11662 6505 11690 6510
rect 12054 6706 12082 6711
rect 11046 6482 11074 6487
rect 11046 5753 11074 6454
rect 11942 6482 11970 6487
rect 11942 6435 11970 6454
rect 12054 6482 12082 6678
rect 12232 6678 12364 6683
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12232 6645 12364 6650
rect 12222 6593 12250 6599
rect 12222 6567 12223 6593
rect 12249 6567 12250 6593
rect 12222 6538 12250 6567
rect 12222 6505 12250 6510
rect 12054 6449 12082 6454
rect 11046 5727 11047 5753
rect 11073 5727 11074 5753
rect 11046 5721 11074 5727
rect 11718 6314 11746 6319
rect 12110 6314 12138 6319
rect 11326 5697 11354 5703
rect 11326 5671 11327 5697
rect 11353 5671 11354 5697
rect 11158 5362 11186 5367
rect 11102 5138 11130 5143
rect 11102 4746 11130 5110
rect 11158 5026 11186 5334
rect 11326 5362 11354 5671
rect 11718 5586 11746 6286
rect 11902 6286 12034 6291
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 11902 6253 12034 6258
rect 11774 6034 11802 6039
rect 11774 5866 11802 6006
rect 11774 5833 11802 5838
rect 11718 5553 11746 5558
rect 11902 5502 12034 5507
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 11902 5469 12034 5474
rect 11326 5329 11354 5334
rect 11158 4993 11186 4998
rect 12110 4802 12138 6286
rect 12232 5894 12364 5899
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12232 5861 12364 5866
rect 12166 5754 12194 5759
rect 12166 5474 12194 5726
rect 12278 5754 12306 5759
rect 12278 5707 12306 5726
rect 12166 5441 12194 5446
rect 12446 5698 12474 5703
rect 12222 5250 12250 5255
rect 12166 5222 12222 5250
rect 12166 5138 12194 5222
rect 12222 5217 12250 5222
rect 12446 5138 12474 5670
rect 12558 5698 12586 5703
rect 12558 5651 12586 5670
rect 12614 5418 12642 6790
rect 13118 6594 13146 7056
rect 14574 7042 14602 7056
rect 14574 7009 14602 7014
rect 14798 7042 14826 7047
rect 13566 6986 13594 6991
rect 13230 6594 13258 6599
rect 13118 6593 13258 6594
rect 13118 6567 13231 6593
rect 13257 6567 13258 6593
rect 13118 6566 13258 6567
rect 13230 6561 13258 6566
rect 12950 6481 12978 6487
rect 12950 6455 12951 6481
rect 12977 6455 12978 6481
rect 12726 6258 12754 6263
rect 12726 5922 12754 6230
rect 12726 5889 12754 5894
rect 12950 5754 12978 6455
rect 13454 5978 13482 5983
rect 12950 5721 12978 5726
rect 13342 5866 13370 5871
rect 12782 5697 12810 5703
rect 12782 5671 12783 5697
rect 12809 5671 12810 5697
rect 12782 5642 12810 5671
rect 12782 5609 12810 5614
rect 13062 5641 13090 5647
rect 13062 5615 13063 5641
rect 13089 5615 13090 5641
rect 12614 5385 12642 5390
rect 12166 5105 12194 5110
rect 12232 5110 12364 5115
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12446 5105 12474 5110
rect 12232 5077 12364 5082
rect 12558 5026 12586 5031
rect 12586 4998 12698 5026
rect 12558 4993 12586 4998
rect 12334 4970 12362 4975
rect 12278 4802 12306 4807
rect 12110 4769 12138 4774
rect 12166 4774 12278 4802
rect 11102 4713 11130 4718
rect 11902 4718 12034 4723
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 11902 4685 12034 4690
rect 11662 4634 11690 4639
rect 11662 4521 11690 4606
rect 11662 4495 11663 4521
rect 11689 4495 11690 4521
rect 11662 4489 11690 4495
rect 11942 4465 11970 4471
rect 11942 4439 11943 4465
rect 11969 4439 11970 4465
rect 11942 4018 11970 4439
rect 12166 4354 12194 4774
rect 12278 4769 12306 4774
rect 12334 4634 12362 4942
rect 12334 4601 12362 4606
rect 12502 4913 12530 4919
rect 12502 4887 12503 4913
rect 12529 4887 12530 4913
rect 12278 4578 12306 4583
rect 12278 4466 12306 4550
rect 12278 4433 12306 4438
rect 12446 4466 12474 4471
rect 12166 4321 12194 4326
rect 12232 4326 12364 4331
rect 11942 3985 11970 3990
rect 12110 4298 12138 4303
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12232 4293 12364 4298
rect 11902 3934 12034 3939
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 11902 3901 12034 3906
rect 10990 3537 11018 3542
rect 11830 3514 11858 3519
rect 10710 3369 10738 3374
rect 11774 3402 11802 3407
rect 11550 3290 11578 3295
rect 11326 3178 11354 3183
rect 10934 2898 10962 2903
rect 10934 2674 10962 2870
rect 10934 2641 10962 2646
rect 11326 2673 11354 3150
rect 11326 2647 11327 2673
rect 11353 2647 11354 2673
rect 11326 2641 11354 2647
rect 11158 2618 11186 2623
rect 11046 2561 11074 2567
rect 11046 2535 11047 2561
rect 11073 2535 11074 2561
rect 10766 2506 10794 2511
rect 10654 2305 10682 2310
rect 10710 2505 10794 2506
rect 10710 2479 10767 2505
rect 10793 2479 10794 2505
rect 10710 2478 10794 2479
rect 10542 1358 10682 1386
rect 10542 1162 10570 1167
rect 10542 1105 10570 1134
rect 10542 1079 10543 1105
rect 10569 1079 10570 1105
rect 10542 1073 10570 1079
rect 10430 401 10458 406
rect 10430 154 10458 159
rect 10430 56 10458 126
rect 10654 56 10682 1358
rect 10710 154 10738 2478
rect 10766 2473 10794 2478
rect 10934 2170 10962 2175
rect 10766 1666 10794 1671
rect 10766 1442 10794 1638
rect 10766 1409 10794 1414
rect 10822 1050 10850 1055
rect 10822 1003 10850 1022
rect 10934 882 10962 2142
rect 10822 854 10962 882
rect 10822 378 10850 854
rect 10822 345 10850 350
rect 10878 770 10906 775
rect 10710 121 10738 126
rect 10878 56 10906 742
rect 11046 658 11074 2535
rect 11046 625 11074 630
rect 11102 1778 11130 1783
rect 11102 56 11130 1750
rect 11158 1106 11186 2590
rect 11494 2114 11522 2119
rect 11494 2067 11522 2086
rect 11158 1073 11186 1078
rect 11214 1778 11242 1783
rect 11214 938 11242 1750
rect 11214 905 11242 910
rect 11326 602 11354 607
rect 11326 56 11354 574
rect 11550 56 11578 3262
rect 11606 2505 11634 2511
rect 11606 2479 11607 2505
rect 11633 2479 11634 2505
rect 11606 1106 11634 2479
rect 11718 2225 11746 2231
rect 11718 2199 11719 2225
rect 11745 2199 11746 2225
rect 11718 1694 11746 2199
rect 11606 1073 11634 1078
rect 11662 1666 11746 1694
rect 11662 602 11690 1666
rect 11662 569 11690 574
rect 11774 56 11802 3374
rect 11830 2674 11858 3486
rect 12110 3290 12138 4270
rect 12446 3794 12474 4438
rect 12502 4186 12530 4887
rect 12502 4153 12530 4158
rect 12614 4242 12642 4247
rect 12446 3761 12474 3766
rect 12232 3542 12364 3547
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12232 3509 12364 3514
rect 12110 3257 12138 3262
rect 12614 3178 12642 4214
rect 12670 3458 12698 4998
rect 12782 4970 12810 4975
rect 12782 4923 12810 4942
rect 13062 4914 13090 5615
rect 13062 4881 13090 4886
rect 12838 4690 12866 4695
rect 12726 4298 12754 4303
rect 12726 3850 12754 4270
rect 12726 3817 12754 3822
rect 12782 4130 12810 4135
rect 12782 3737 12810 4102
rect 12782 3711 12783 3737
rect 12809 3711 12810 3737
rect 12782 3705 12810 3711
rect 12670 3425 12698 3430
rect 12726 3570 12754 3575
rect 11902 3150 12034 3155
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12614 3145 12642 3150
rect 12670 3234 12698 3239
rect 11902 3117 12034 3122
rect 12614 3066 12642 3071
rect 12232 2758 12364 2763
rect 12166 2730 12194 2735
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12232 2725 12364 2730
rect 12446 2730 12474 2735
rect 12166 2674 12194 2702
rect 12446 2674 12474 2702
rect 12166 2646 12474 2674
rect 11830 2641 11858 2646
rect 12614 2394 12642 3038
rect 11902 2366 12034 2371
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12614 2361 12642 2366
rect 11902 2333 12034 2338
rect 12614 2057 12642 2063
rect 12614 2031 12615 2057
rect 12641 2031 12642 2057
rect 12232 1974 12364 1979
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12232 1941 12364 1946
rect 12614 1834 12642 2031
rect 12614 1801 12642 1806
rect 11902 1582 12034 1587
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 11902 1549 12034 1554
rect 12166 1554 12194 1559
rect 12166 1218 12194 1526
rect 12558 1554 12586 1559
rect 12670 1554 12698 3206
rect 12726 2282 12754 3542
rect 12838 3402 12866 4662
rect 13342 4354 13370 5838
rect 13454 5810 13482 5950
rect 13454 5777 13482 5782
rect 13454 5530 13482 5535
rect 13342 4321 13370 4326
rect 13398 5194 13426 5199
rect 13006 4242 13034 4247
rect 12838 3369 12866 3374
rect 12894 4018 12922 4023
rect 12894 2954 12922 3990
rect 12894 2921 12922 2926
rect 12726 2249 12754 2254
rect 12782 2786 12810 2791
rect 12586 1526 12698 1554
rect 12558 1521 12586 1526
rect 12166 1185 12194 1190
rect 12232 1190 12364 1195
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12232 1157 12364 1162
rect 12614 994 12642 999
rect 12614 993 12698 994
rect 12614 967 12615 993
rect 12641 967 12698 993
rect 12614 966 12698 967
rect 12614 961 12642 966
rect 12390 938 12418 943
rect 12390 891 12418 910
rect 11902 798 12034 803
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 11902 765 12034 770
rect 11998 658 12026 663
rect 11998 56 12026 630
rect 12446 490 12474 495
rect 12232 406 12364 411
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12232 373 12364 378
rect 12222 266 12250 271
rect 12222 56 12250 238
rect 12446 56 12474 462
rect 12670 56 12698 966
rect 12782 882 12810 2758
rect 12894 2113 12922 2119
rect 12894 2087 12895 2113
rect 12921 2087 12922 2113
rect 12894 1778 12922 2087
rect 12894 1745 12922 1750
rect 13006 1442 13034 4214
rect 13398 4186 13426 5166
rect 13454 5026 13482 5502
rect 13566 5530 13594 6958
rect 14798 6425 14826 7014
rect 16030 7042 16058 7056
rect 16030 7009 16058 7014
rect 16254 7042 16282 7047
rect 15750 6818 15778 6823
rect 14798 6399 14799 6425
rect 14825 6399 14826 6425
rect 14798 6393 14826 6399
rect 15302 6481 15330 6487
rect 15302 6455 15303 6481
rect 15329 6455 15330 6481
rect 14294 6370 14322 6375
rect 13566 5497 13594 5502
rect 13790 6258 13818 6263
rect 13454 4993 13482 4998
rect 13398 4153 13426 4158
rect 13678 4130 13706 4135
rect 13398 3962 13426 3967
rect 13062 3794 13090 3799
rect 13062 3747 13090 3766
rect 13342 3458 13370 3463
rect 13342 3346 13370 3430
rect 13342 3313 13370 3318
rect 13118 3290 13146 3295
rect 13118 2673 13146 3262
rect 13118 2647 13119 2673
rect 13145 2647 13146 2673
rect 13118 2641 13146 2647
rect 13398 2617 13426 3934
rect 13678 3737 13706 4102
rect 13678 3711 13679 3737
rect 13705 3711 13706 3737
rect 13678 3705 13706 3711
rect 13790 3682 13818 6230
rect 14238 6034 14266 6039
rect 14238 5642 14266 6006
rect 14238 5609 14266 5614
rect 14126 5474 14154 5479
rect 14014 4802 14042 4807
rect 13790 3649 13818 3654
rect 13846 4018 13874 4023
rect 13398 2591 13399 2617
rect 13425 2591 13426 2617
rect 13398 2585 13426 2591
rect 13734 2618 13762 2623
rect 13454 2562 13482 2567
rect 13454 2058 13482 2534
rect 13454 2025 13482 2030
rect 13510 2226 13538 2231
rect 13006 1409 13034 1414
rect 13174 1610 13202 1615
rect 12838 1386 12866 1391
rect 12838 1105 12866 1358
rect 12838 1079 12839 1105
rect 12865 1079 12866 1105
rect 12838 1073 12866 1079
rect 12782 849 12810 854
rect 13118 937 13146 943
rect 13118 911 13119 937
rect 13145 911 13146 937
rect 12950 602 12978 607
rect 12894 601 12978 602
rect 12894 575 12951 601
rect 12977 575 12978 601
rect 12894 574 12978 575
rect 12894 546 12922 574
rect 12950 569 12978 574
rect 13118 602 13146 911
rect 13118 569 13146 574
rect 12894 513 12922 518
rect 13174 490 13202 1582
rect 13286 1498 13314 1503
rect 13286 1105 13314 1470
rect 13510 1498 13538 2198
rect 13678 2057 13706 2063
rect 13678 2031 13679 2057
rect 13705 2031 13706 2057
rect 13678 1890 13706 2031
rect 13678 1857 13706 1862
rect 13734 1777 13762 2590
rect 13734 1751 13735 1777
rect 13761 1751 13762 1777
rect 13734 1745 13762 1751
rect 13846 1610 13874 3990
rect 13958 3682 13986 3687
rect 13958 3635 13986 3654
rect 14014 3122 14042 4774
rect 14014 3089 14042 3094
rect 14070 4522 14098 4527
rect 14070 2618 14098 4494
rect 14126 3906 14154 5446
rect 14238 5250 14266 5255
rect 14182 4634 14210 4639
rect 14182 4130 14210 4606
rect 14238 4214 14266 5222
rect 14294 4521 14322 6342
rect 14798 5922 14826 5927
rect 14686 5697 14714 5703
rect 14686 5671 14687 5697
rect 14713 5671 14714 5697
rect 14686 5306 14714 5671
rect 14686 5273 14714 5278
rect 14518 4578 14546 4583
rect 14518 4531 14546 4550
rect 14294 4495 14295 4521
rect 14321 4495 14322 4521
rect 14294 4489 14322 4495
rect 14238 4186 14770 4214
rect 14182 4097 14210 4102
rect 14126 3873 14154 3878
rect 14070 2585 14098 2590
rect 14126 3738 14154 3743
rect 14014 2282 14042 2287
rect 13846 1577 13874 1582
rect 13902 2225 13930 2231
rect 13902 2199 13903 2225
rect 13929 2199 13930 2225
rect 13510 1465 13538 1470
rect 13902 1386 13930 2199
rect 13958 1834 13986 1839
rect 14014 1834 14042 2254
rect 13958 1833 14042 1834
rect 13958 1807 13959 1833
rect 13985 1807 14042 1833
rect 13958 1806 14042 1807
rect 14126 1833 14154 3710
rect 14742 3737 14770 4186
rect 14742 3711 14743 3737
rect 14769 3711 14770 3737
rect 14742 3705 14770 3711
rect 14294 3514 14322 3519
rect 14126 1807 14127 1833
rect 14153 1807 14154 1833
rect 13958 1801 13986 1806
rect 14126 1801 14154 1807
rect 14182 3066 14210 3071
rect 14182 1610 14210 3038
rect 14294 1946 14322 3486
rect 14798 3066 14826 5894
rect 14966 5810 14994 5815
rect 14966 5753 14994 5782
rect 14966 5727 14967 5753
rect 14993 5727 14994 5753
rect 14966 5721 14994 5727
rect 15302 5754 15330 6455
rect 15302 5721 15330 5726
rect 15694 5418 15722 5423
rect 14966 5250 14994 5255
rect 14854 5194 14882 5199
rect 14854 3234 14882 5166
rect 14910 4242 14938 4247
rect 14910 3402 14938 4214
rect 14966 3794 14994 5222
rect 15638 5194 15666 5199
rect 15638 5147 15666 5166
rect 15190 5138 15218 5143
rect 15134 4522 15162 4527
rect 15134 4074 15162 4494
rect 15134 4041 15162 4046
rect 14966 3761 14994 3766
rect 15078 3850 15106 3855
rect 15022 3738 15050 3743
rect 15022 3691 15050 3710
rect 14910 3369 14938 3374
rect 14854 3201 14882 3206
rect 14798 3033 14826 3038
rect 15078 3010 15106 3822
rect 15190 3234 15218 5110
rect 15694 4214 15722 5390
rect 15638 4186 15722 4214
rect 15582 3402 15610 3407
rect 15358 3346 15386 3351
rect 15358 3299 15386 3318
rect 15190 3201 15218 3206
rect 15022 2982 15106 3010
rect 14294 1913 14322 1918
rect 14350 2842 14378 2847
rect 14182 1577 14210 1582
rect 14294 1834 14322 1839
rect 14294 1442 14322 1806
rect 14294 1409 14322 1414
rect 13902 1353 13930 1358
rect 14350 1385 14378 2814
rect 14742 2394 14770 2399
rect 14686 1890 14714 1895
rect 14350 1359 14351 1385
rect 14377 1359 14378 1385
rect 14350 1353 14378 1359
rect 14406 1665 14434 1671
rect 14406 1639 14407 1665
rect 14433 1639 14434 1665
rect 13958 1329 13986 1335
rect 13958 1303 13959 1329
rect 13985 1303 13986 1329
rect 13678 1274 13706 1279
rect 13678 1227 13706 1246
rect 13846 1274 13874 1279
rect 13286 1079 13287 1105
rect 13313 1079 13314 1105
rect 13286 1073 13314 1079
rect 13454 1162 13482 1167
rect 13342 546 13370 551
rect 13342 499 13370 518
rect 13118 462 13202 490
rect 12894 434 12922 439
rect 12894 56 12922 406
rect 13118 56 13146 462
rect 13454 210 13482 1134
rect 13734 994 13762 999
rect 13734 947 13762 966
rect 13566 937 13594 943
rect 13566 911 13567 937
rect 13593 911 13594 937
rect 13566 658 13594 911
rect 13566 625 13594 630
rect 13790 546 13818 551
rect 13454 177 13482 182
rect 13566 378 13594 383
rect 13342 154 13370 159
rect 13342 56 13370 126
rect 13566 56 13594 350
rect 13790 56 13818 518
rect 13846 322 13874 1246
rect 13958 1218 13986 1303
rect 13958 1185 13986 1190
rect 14070 1106 14098 1111
rect 14070 601 14098 1078
rect 14070 575 14071 601
rect 14097 575 14098 601
rect 14070 569 14098 575
rect 14238 881 14266 887
rect 14238 855 14239 881
rect 14265 855 14266 881
rect 13846 289 13874 294
rect 14014 490 14042 495
rect 14014 56 14042 462
rect 14238 56 14266 855
rect 14406 490 14434 1639
rect 14630 1274 14658 1279
rect 14406 457 14434 462
rect 14462 1273 14658 1274
rect 14462 1247 14631 1273
rect 14657 1247 14658 1273
rect 14462 1246 14658 1247
rect 14462 56 14490 1246
rect 14630 1241 14658 1246
rect 14686 1162 14714 1862
rect 14686 1129 14714 1134
rect 14518 1050 14546 1055
rect 14518 1003 14546 1022
rect 14742 714 14770 2366
rect 14742 681 14770 686
rect 14910 937 14938 943
rect 14910 911 14911 937
rect 14937 911 14938 937
rect 14574 658 14602 663
rect 14574 657 14714 658
rect 14574 631 14575 657
rect 14601 631 14714 657
rect 14574 630 14714 631
rect 14574 625 14602 630
rect 14686 56 14714 630
rect 14854 602 14882 607
rect 14854 555 14882 574
rect 14910 56 14938 911
rect 15022 434 15050 2982
rect 15078 2898 15106 2903
rect 15078 1554 15106 2870
rect 15582 1890 15610 3374
rect 15638 3401 15666 4186
rect 15638 3375 15639 3401
rect 15665 3375 15666 3401
rect 15638 3369 15666 3375
rect 15638 1890 15666 1895
rect 15582 1889 15666 1890
rect 15582 1863 15639 1889
rect 15665 1863 15666 1889
rect 15582 1862 15666 1863
rect 15638 1857 15666 1862
rect 15190 1777 15218 1783
rect 15190 1751 15191 1777
rect 15217 1751 15218 1777
rect 15190 1722 15218 1751
rect 15526 1778 15554 1783
rect 15190 1689 15218 1694
rect 15470 1721 15498 1727
rect 15470 1695 15471 1721
rect 15497 1695 15498 1721
rect 15078 1521 15106 1526
rect 15134 1330 15162 1335
rect 15134 1283 15162 1302
rect 15414 1274 15442 1279
rect 15190 1273 15442 1274
rect 15190 1247 15415 1273
rect 15441 1247 15442 1273
rect 15190 1246 15442 1247
rect 15190 658 15218 1246
rect 15414 1241 15442 1246
rect 15470 1050 15498 1695
rect 15470 1017 15498 1022
rect 15414 993 15442 999
rect 15414 967 15415 993
rect 15441 967 15442 993
rect 15414 938 15442 967
rect 15526 938 15554 1750
rect 15414 910 15554 938
rect 15638 1610 15666 1615
rect 15582 881 15610 887
rect 15582 855 15583 881
rect 15609 855 15610 881
rect 15022 401 15050 406
rect 15134 630 15218 658
rect 15358 657 15386 663
rect 15358 631 15359 657
rect 15385 631 15386 657
rect 15134 56 15162 630
rect 15358 56 15386 631
rect 15582 56 15610 855
rect 15638 490 15666 1582
rect 15750 1610 15778 6790
rect 16254 6425 16282 7014
rect 17486 7042 17514 7056
rect 17486 7009 17514 7014
rect 17766 7042 17794 7047
rect 16254 6399 16255 6425
rect 16281 6399 16282 6425
rect 16254 6393 16282 6399
rect 16702 6818 16730 6823
rect 16534 6314 16562 6319
rect 16478 5978 16506 5983
rect 16422 5977 16506 5978
rect 16422 5951 16479 5977
rect 16505 5951 16506 5977
rect 16422 5950 16506 5951
rect 16198 5754 16226 5759
rect 16198 5707 16226 5726
rect 16422 5642 16450 5950
rect 16478 5945 16506 5950
rect 16422 5609 16450 5614
rect 16478 5697 16506 5703
rect 16478 5671 16479 5697
rect 16505 5671 16506 5697
rect 15806 5530 15834 5535
rect 15806 1666 15834 5502
rect 15918 5249 15946 5255
rect 15918 5223 15919 5249
rect 15945 5223 15946 5249
rect 15918 5138 15946 5223
rect 15918 5105 15946 5110
rect 16310 5082 16338 5087
rect 15974 4858 16002 4863
rect 15974 2674 16002 4830
rect 16310 4802 16338 5054
rect 16310 4769 16338 4774
rect 16030 4466 16058 4471
rect 16030 3290 16058 4438
rect 16478 4214 16506 5671
rect 16534 5025 16562 6286
rect 16534 4999 16535 5025
rect 16561 4999 16562 5025
rect 16534 4993 16562 4999
rect 16646 6258 16674 6263
rect 16478 4186 16562 4214
rect 16030 3257 16058 3262
rect 15974 2641 16002 2646
rect 16142 2842 16170 2847
rect 15974 2114 16002 2119
rect 15974 2067 16002 2086
rect 15918 1834 15946 1839
rect 15918 1787 15946 1806
rect 15806 1633 15834 1638
rect 15750 1577 15778 1582
rect 15974 1386 16002 1391
rect 15974 1339 16002 1358
rect 15862 1274 15890 1279
rect 15806 658 15834 663
rect 15806 601 15834 630
rect 15806 575 15807 601
rect 15833 575 15834 601
rect 15806 569 15834 575
rect 15862 490 15890 1246
rect 16086 490 16114 495
rect 15638 457 15666 462
rect 15806 462 15890 490
rect 16030 489 16114 490
rect 16030 463 16087 489
rect 16113 463 16114 489
rect 16030 462 16114 463
rect 15806 56 15834 462
rect 16030 56 16058 462
rect 16086 457 16114 462
rect 16142 378 16170 2814
rect 16422 2562 16450 2567
rect 16254 2114 16282 2119
rect 16254 2067 16282 2086
rect 16198 1890 16226 1895
rect 16198 1843 16226 1862
rect 16422 1610 16450 2534
rect 16478 2450 16506 2455
rect 16478 2169 16506 2422
rect 16534 2226 16562 4186
rect 16534 2193 16562 2198
rect 16590 2450 16618 2455
rect 16478 2143 16479 2169
rect 16505 2143 16506 2169
rect 16478 2137 16506 2143
rect 16478 1834 16506 1839
rect 16590 1834 16618 2422
rect 16646 2394 16674 6230
rect 16702 5754 16730 6790
rect 17318 6762 17346 6767
rect 16758 6482 16786 6487
rect 16758 6435 16786 6454
rect 16814 6370 16842 6375
rect 16758 6034 16786 6039
rect 16758 5987 16786 6006
rect 16814 5922 16842 6342
rect 17318 6089 17346 6734
rect 17318 6063 17319 6089
rect 17345 6063 17346 6089
rect 17318 6057 17346 6063
rect 17486 6482 17514 6487
rect 16702 5721 16730 5726
rect 16758 5894 16842 5922
rect 17206 6034 17234 6039
rect 16758 5642 16786 5894
rect 16702 5614 16786 5642
rect 16702 4858 16730 5614
rect 16758 5306 16786 5311
rect 16758 4970 16786 5278
rect 16758 4937 16786 4942
rect 16870 5082 16898 5087
rect 16758 4858 16786 4863
rect 16702 4857 16786 4858
rect 16702 4831 16759 4857
rect 16785 4831 16786 4857
rect 16702 4830 16786 4831
rect 16758 4825 16786 4830
rect 16870 4746 16898 5054
rect 16814 4718 16898 4746
rect 16758 4354 16786 4359
rect 16758 3570 16786 4326
rect 16814 4130 16842 4718
rect 16926 4522 16954 4527
rect 16926 4354 16954 4494
rect 16982 4410 17010 4415
rect 16982 4363 17010 4382
rect 16926 4321 16954 4326
rect 16814 4097 16842 4102
rect 16870 4298 16898 4303
rect 16814 3570 16842 3575
rect 16758 3542 16814 3570
rect 16814 3537 16842 3542
rect 16758 3458 16786 3463
rect 16870 3458 16898 4270
rect 16786 3430 16898 3458
rect 16758 3425 16786 3430
rect 16646 2361 16674 2366
rect 16702 3402 16730 3407
rect 16702 2170 16730 3374
rect 16758 3010 16786 3015
rect 16758 2506 16786 2982
rect 16982 2674 17010 2679
rect 16982 2627 17010 2646
rect 17206 2674 17234 6006
rect 17262 4522 17290 4527
rect 17262 4475 17290 4494
rect 17486 3793 17514 6454
rect 17766 6425 17794 7014
rect 18438 6538 18466 6543
rect 18942 6538 18970 7056
rect 20398 7042 20426 7056
rect 20398 7009 20426 7014
rect 20622 7042 20650 7047
rect 18942 6510 19194 6538
rect 18270 6482 18298 6487
rect 18270 6435 18298 6454
rect 17766 6399 17767 6425
rect 17793 6399 17794 6425
rect 17766 6393 17794 6399
rect 17598 6033 17626 6039
rect 17598 6007 17599 6033
rect 17625 6007 17626 6033
rect 17598 5922 17626 6007
rect 17598 5889 17626 5894
rect 18382 5698 18410 5703
rect 18382 4970 18410 5670
rect 18438 5474 18466 6510
rect 19166 6201 19194 6510
rect 19166 6175 19167 6201
rect 19193 6175 19194 6201
rect 19166 6169 19194 6175
rect 19222 6482 19250 6487
rect 18606 6146 18634 6151
rect 18606 6089 18634 6118
rect 18606 6063 18607 6089
rect 18633 6063 18634 6089
rect 18606 6057 18634 6063
rect 18886 6034 18914 6039
rect 18886 5987 18914 6006
rect 18774 5978 18802 5983
rect 18438 5441 18466 5446
rect 18494 5866 18522 5871
rect 18494 5305 18522 5838
rect 18718 5586 18746 5591
rect 18718 5361 18746 5558
rect 18718 5335 18719 5361
rect 18745 5335 18746 5361
rect 18718 5329 18746 5335
rect 18494 5279 18495 5305
rect 18521 5279 18522 5305
rect 18494 5273 18522 5279
rect 18382 4937 18410 4942
rect 18718 5026 18746 5031
rect 18718 4969 18746 4998
rect 18718 4943 18719 4969
rect 18745 4943 18746 4969
rect 18718 4937 18746 4943
rect 18494 4913 18522 4919
rect 18494 4887 18495 4913
rect 18521 4887 18522 4913
rect 18270 4746 18298 4751
rect 17486 3767 17487 3793
rect 17513 3767 17514 3793
rect 17486 3761 17514 3767
rect 17542 4354 17570 4359
rect 17542 2953 17570 4326
rect 17766 3906 17794 3911
rect 17766 3737 17794 3878
rect 17766 3711 17767 3737
rect 17793 3711 17794 3737
rect 17766 3705 17794 3711
rect 18214 3625 18242 3631
rect 18214 3599 18215 3625
rect 18241 3599 18242 3625
rect 17542 2927 17543 2953
rect 17569 2927 17570 2953
rect 17542 2921 17570 2927
rect 17766 3514 17794 3519
rect 17206 2641 17234 2646
rect 16758 2473 16786 2478
rect 17206 2505 17234 2511
rect 17206 2479 17207 2505
rect 17233 2479 17234 2505
rect 16702 2137 16730 2142
rect 16478 1833 16618 1834
rect 16478 1807 16479 1833
rect 16505 1807 16618 1833
rect 16478 1806 16618 1807
rect 16758 2113 16786 2119
rect 16758 2087 16759 2113
rect 16785 2087 16786 2113
rect 16478 1801 16506 1806
rect 16422 1577 16450 1582
rect 16198 1274 16226 1279
rect 16198 1227 16226 1246
rect 16366 1050 16394 1055
rect 16366 1003 16394 1022
rect 16758 1050 16786 2087
rect 16814 1442 16842 1447
rect 16814 1385 16842 1414
rect 16814 1359 16815 1385
rect 16841 1359 16842 1385
rect 16814 1353 16842 1359
rect 16758 1017 16786 1022
rect 17038 1329 17066 1335
rect 17038 1303 17039 1329
rect 17065 1303 17066 1329
rect 16142 345 16170 350
rect 16198 882 16226 887
rect 16646 882 16674 887
rect 16198 266 16226 854
rect 16198 233 16226 238
rect 16254 881 16674 882
rect 16254 855 16647 881
rect 16673 855 16674 881
rect 16254 854 16674 855
rect 16254 56 16282 854
rect 16646 849 16674 854
rect 16758 882 16786 887
rect 16702 658 16730 663
rect 16478 657 16730 658
rect 16478 631 16703 657
rect 16729 631 16730 657
rect 16478 630 16730 631
rect 16478 56 16506 630
rect 16702 625 16730 630
rect 16758 434 16786 854
rect 17038 602 17066 1303
rect 17150 1218 17178 1223
rect 17150 1049 17178 1190
rect 17150 1023 17151 1049
rect 17177 1023 17178 1049
rect 17150 1017 17178 1023
rect 17150 658 17178 663
rect 17094 602 17122 607
rect 17038 601 17122 602
rect 17038 575 17095 601
rect 17121 575 17122 601
rect 17038 574 17122 575
rect 17094 569 17122 574
rect 16702 406 16786 434
rect 16926 490 16954 495
rect 16702 56 16730 406
rect 16926 56 16954 462
rect 17150 56 17178 630
rect 17206 602 17234 2479
rect 17262 2114 17290 2119
rect 17262 1385 17290 2086
rect 17766 1890 17794 3486
rect 18158 3402 18186 3407
rect 18158 3178 18186 3374
rect 18158 3145 18186 3150
rect 17822 2898 17850 2903
rect 17822 2897 18186 2898
rect 17822 2871 17823 2897
rect 17849 2871 18186 2897
rect 17822 2870 18186 2871
rect 17822 2865 17850 2870
rect 17934 1890 17962 1895
rect 17766 1889 17962 1890
rect 17766 1863 17935 1889
rect 17961 1863 17962 1889
rect 17766 1862 17962 1863
rect 17934 1857 17962 1862
rect 17262 1359 17263 1385
rect 17289 1359 17290 1385
rect 17262 1353 17290 1359
rect 18158 1385 18186 2870
rect 18214 2730 18242 3599
rect 18214 2697 18242 2702
rect 18214 1722 18242 1727
rect 18214 1675 18242 1694
rect 18158 1359 18159 1385
rect 18185 1359 18186 1385
rect 18158 1353 18186 1359
rect 18270 1386 18298 4718
rect 18494 4466 18522 4887
rect 18494 4433 18522 4438
rect 18438 4354 18466 4359
rect 18438 4074 18466 4326
rect 18438 4041 18466 4046
rect 18494 3682 18522 3687
rect 18494 3681 18746 3682
rect 18494 3655 18495 3681
rect 18521 3655 18746 3681
rect 18494 3654 18746 3655
rect 18494 3649 18522 3654
rect 18382 3570 18410 3575
rect 18382 3178 18410 3542
rect 18382 3145 18410 3150
rect 18438 3234 18466 3239
rect 18270 1353 18298 1358
rect 18326 2226 18354 2231
rect 17654 1329 17682 1335
rect 17654 1303 17655 1329
rect 17681 1303 17682 1329
rect 17598 1106 17626 1111
rect 17206 569 17234 574
rect 17374 994 17402 999
rect 17374 56 17402 966
rect 17430 882 17458 887
rect 17430 835 17458 854
rect 17598 714 17626 1078
rect 17598 681 17626 686
rect 17654 658 17682 1303
rect 17934 1050 17962 1055
rect 17934 1003 17962 1022
rect 18214 994 18242 999
rect 18214 937 18242 966
rect 18214 911 18215 937
rect 18241 911 18242 937
rect 18214 905 18242 911
rect 18046 882 18074 887
rect 17654 625 17682 630
rect 17822 658 17850 663
rect 17654 546 17682 551
rect 17654 499 17682 518
rect 17598 434 17626 439
rect 17598 56 17626 406
rect 17822 56 17850 630
rect 17934 490 17962 495
rect 17934 443 17962 462
rect 18046 56 18074 854
rect 18270 826 18298 831
rect 18270 56 18298 798
rect 18326 154 18354 2198
rect 18438 2170 18466 3206
rect 18438 2137 18466 2142
rect 18494 2730 18522 2735
rect 18382 1946 18410 1951
rect 18382 1833 18410 1918
rect 18382 1807 18383 1833
rect 18409 1807 18410 1833
rect 18382 1801 18410 1807
rect 18438 1890 18466 1895
rect 18438 1554 18466 1862
rect 18438 1521 18466 1526
rect 18494 1442 18522 2702
rect 18494 1409 18522 1414
rect 18662 1665 18690 1671
rect 18662 1639 18663 1665
rect 18689 1639 18690 1665
rect 18550 1329 18578 1335
rect 18550 1303 18551 1329
rect 18577 1303 18578 1329
rect 18382 714 18410 719
rect 18382 322 18410 686
rect 18550 658 18578 1303
rect 18662 826 18690 1639
rect 18718 1049 18746 3654
rect 18774 1610 18802 5950
rect 19054 5922 19082 5927
rect 18886 4298 18914 4303
rect 18886 4241 18914 4270
rect 18886 4215 18887 4241
rect 18913 4215 18914 4241
rect 18886 4209 18914 4215
rect 18830 2170 18858 2175
rect 18830 2123 18858 2142
rect 18774 1577 18802 1582
rect 18942 1386 18970 1391
rect 18942 1339 18970 1358
rect 18718 1023 18719 1049
rect 18745 1023 18746 1049
rect 18718 1017 18746 1023
rect 18774 1274 18802 1279
rect 18662 793 18690 798
rect 18550 625 18578 630
rect 18438 602 18466 607
rect 18438 555 18466 574
rect 18382 289 18410 294
rect 18494 546 18522 551
rect 18326 121 18354 126
rect 18494 56 18522 518
rect 18718 490 18746 495
rect 18718 443 18746 462
rect 18774 378 18802 1246
rect 19054 1162 19082 5894
rect 19166 4410 19194 4415
rect 19166 4185 19194 4382
rect 19166 4159 19167 4185
rect 19193 4159 19194 4185
rect 19166 4153 19194 4159
rect 19166 2618 19194 2623
rect 19166 2571 19194 2590
rect 19110 2114 19138 2119
rect 19110 2067 19138 2086
rect 19166 1778 19194 1783
rect 19166 1731 19194 1750
rect 19222 1386 19250 6454
rect 20622 6425 20650 7014
rect 21854 7042 21882 7056
rect 21854 7009 21882 7014
rect 22078 7042 22106 7047
rect 21126 6482 21154 6487
rect 21126 6481 21266 6482
rect 21126 6455 21127 6481
rect 21153 6455 21266 6481
rect 21126 6454 21266 6455
rect 21126 6449 21154 6454
rect 20622 6399 20623 6425
rect 20649 6399 20650 6425
rect 20622 6393 20650 6399
rect 20846 6090 20874 6095
rect 20846 6043 20874 6062
rect 21126 6090 21154 6095
rect 21126 6043 21154 6062
rect 19670 6033 19698 6039
rect 19670 6007 19671 6033
rect 19697 6007 19698 6033
rect 19446 5697 19474 5703
rect 19446 5671 19447 5697
rect 19473 5671 19474 5697
rect 19446 5082 19474 5671
rect 19446 5049 19474 5054
rect 19558 4802 19586 4807
rect 19446 4466 19474 4471
rect 19446 2617 19474 4438
rect 19446 2591 19447 2617
rect 19473 2591 19474 2617
rect 19446 2585 19474 2591
rect 19222 1353 19250 1358
rect 19446 1721 19474 1727
rect 19446 1695 19447 1721
rect 19473 1695 19474 1721
rect 19222 1274 19250 1279
rect 19222 1227 19250 1246
rect 19054 1129 19082 1134
rect 18998 882 19026 887
rect 18998 835 19026 854
rect 19166 882 19194 887
rect 18718 350 18802 378
rect 18942 490 18970 495
rect 18718 56 18746 350
rect 18942 56 18970 462
rect 19166 56 19194 854
rect 19446 434 19474 1695
rect 19446 401 19474 406
rect 19502 993 19530 999
rect 19502 967 19503 993
rect 19529 967 19530 993
rect 19502 378 19530 967
rect 19558 601 19586 4774
rect 19670 4242 19698 6007
rect 20678 6034 20706 6039
rect 20678 6033 20762 6034
rect 20678 6007 20679 6033
rect 20705 6007 20762 6033
rect 20678 6006 20762 6007
rect 20678 6001 20706 6006
rect 20398 5978 20426 5983
rect 20398 5931 20426 5950
rect 19726 5642 19754 5647
rect 19726 5595 19754 5614
rect 20286 4802 20314 4807
rect 20118 4690 20146 4695
rect 19670 4209 19698 4214
rect 20006 4409 20034 4415
rect 20006 4383 20007 4409
rect 20033 4383 20034 4409
rect 20006 2730 20034 4383
rect 20118 3346 20146 4662
rect 20286 4577 20314 4774
rect 20286 4551 20287 4577
rect 20313 4551 20314 4577
rect 20286 4545 20314 4551
rect 20566 4354 20594 4359
rect 20118 3313 20146 3318
rect 20342 3850 20370 3855
rect 20006 2697 20034 2702
rect 20342 2170 20370 3822
rect 20566 3737 20594 4326
rect 20566 3711 20567 3737
rect 20593 3711 20594 3737
rect 20566 3705 20594 3711
rect 20678 3850 20706 3855
rect 20398 3178 20426 3183
rect 20398 2953 20426 3150
rect 20678 3009 20706 3822
rect 20678 2983 20679 3009
rect 20705 2983 20706 3009
rect 20678 2977 20706 2983
rect 20398 2927 20399 2953
rect 20425 2927 20426 2953
rect 20398 2921 20426 2927
rect 20734 2338 20762 6006
rect 20958 5978 20986 5983
rect 20958 5754 20986 5950
rect 20958 5721 20986 5726
rect 20958 4186 20986 4191
rect 20902 3794 20930 3799
rect 20846 3681 20874 3687
rect 20846 3655 20847 3681
rect 20873 3655 20874 3681
rect 20790 3626 20818 3631
rect 20790 3290 20818 3598
rect 20790 3257 20818 3262
rect 20846 3010 20874 3655
rect 20846 2977 20874 2982
rect 20902 2394 20930 3766
rect 20958 2506 20986 4158
rect 21070 4186 21098 4191
rect 21070 3906 21098 4158
rect 21070 3873 21098 3878
rect 20958 2473 20986 2478
rect 20902 2361 20930 2366
rect 20734 2305 20762 2310
rect 20342 2137 20370 2142
rect 20454 2113 20482 2119
rect 20454 2087 20455 2113
rect 20481 2087 20482 2113
rect 20174 2057 20202 2063
rect 20174 2031 20175 2057
rect 20201 2031 20202 2057
rect 20174 2002 20202 2031
rect 20174 1969 20202 1974
rect 19726 1722 19754 1727
rect 19726 1385 19754 1694
rect 19726 1359 19727 1385
rect 19753 1359 19754 1385
rect 19726 1353 19754 1359
rect 19894 1722 19922 1727
rect 19558 575 19559 601
rect 19585 575 19586 601
rect 19558 569 19586 575
rect 19614 1106 19642 1111
rect 19502 345 19530 350
rect 19390 322 19418 327
rect 19390 56 19418 294
rect 19614 56 19642 1078
rect 19782 994 19810 999
rect 19782 947 19810 966
rect 19838 546 19866 551
rect 19838 489 19866 518
rect 19838 463 19839 489
rect 19865 463 19866 489
rect 19838 457 19866 463
rect 19894 378 19922 1694
rect 20230 1722 20258 1741
rect 20230 1689 20258 1694
rect 20342 1498 20370 1503
rect 20006 1273 20034 1279
rect 20006 1247 20007 1273
rect 20033 1247 20034 1273
rect 20006 882 20034 1247
rect 20174 1274 20202 1279
rect 20118 994 20146 999
rect 20118 947 20146 966
rect 20006 849 20034 854
rect 19838 350 19922 378
rect 20062 658 20090 663
rect 19838 56 19866 350
rect 20062 56 20090 630
rect 20174 266 20202 1246
rect 20174 233 20202 238
rect 20230 994 20258 999
rect 20230 210 20258 966
rect 20342 601 20370 1470
rect 20454 1386 20482 2087
rect 20510 2114 20538 2119
rect 20510 1498 20538 2086
rect 20734 2114 20762 2119
rect 20734 1833 20762 2086
rect 21070 2114 21098 2119
rect 21070 2067 21098 2086
rect 20790 2058 20818 2063
rect 20790 2011 20818 2030
rect 20734 1807 20735 1833
rect 20761 1807 20762 1833
rect 20734 1801 20762 1807
rect 21014 1721 21042 1727
rect 21014 1695 21015 1721
rect 21041 1695 21042 1721
rect 21014 1694 21042 1695
rect 20510 1465 20538 1470
rect 20734 1666 21042 1694
rect 20510 1386 20538 1391
rect 20454 1385 20538 1386
rect 20454 1359 20511 1385
rect 20537 1359 20538 1385
rect 20454 1358 20538 1359
rect 20510 1353 20538 1358
rect 20342 575 20343 601
rect 20369 575 20370 601
rect 20342 569 20370 575
rect 20398 881 20426 887
rect 20398 855 20399 881
rect 20425 855 20426 881
rect 20230 177 20258 182
rect 20286 546 20314 551
rect 20286 56 20314 518
rect 20398 322 20426 855
rect 20398 289 20426 294
rect 20510 826 20538 831
rect 20510 56 20538 798
rect 20622 490 20650 495
rect 20622 443 20650 462
rect 20734 56 20762 1666
rect 21238 1442 21266 6454
rect 22078 6425 22106 7014
rect 23310 7042 23338 7056
rect 23310 7009 23338 7014
rect 23534 7042 23562 7047
rect 22232 6678 22364 6683
rect 22260 6650 22284 6678
rect 22312 6650 22336 6678
rect 22232 6645 22364 6650
rect 22582 6482 22610 6487
rect 22582 6481 22666 6482
rect 22582 6455 22583 6481
rect 22609 6455 22666 6481
rect 22582 6454 22666 6455
rect 22582 6449 22610 6454
rect 22078 6399 22079 6425
rect 22105 6399 22106 6425
rect 22078 6393 22106 6399
rect 21902 6286 22034 6291
rect 21930 6258 21954 6286
rect 21982 6258 22006 6286
rect 21902 6253 22034 6258
rect 22232 5894 22364 5899
rect 22260 5866 22284 5894
rect 22312 5866 22336 5894
rect 22232 5861 22364 5866
rect 21742 5697 21770 5703
rect 21742 5671 21743 5697
rect 21769 5671 21770 5697
rect 21742 5530 21770 5671
rect 21742 5497 21770 5502
rect 21798 5698 21826 5703
rect 21518 5474 21546 5479
rect 21462 2562 21490 2567
rect 21462 1777 21490 2534
rect 21518 2169 21546 5446
rect 21798 4970 21826 5670
rect 22022 5642 22050 5647
rect 22022 5641 22106 5642
rect 22022 5615 22023 5641
rect 22049 5615 22106 5641
rect 22022 5614 22106 5615
rect 22022 5609 22050 5614
rect 21902 5502 22034 5507
rect 21930 5474 21954 5502
rect 21982 5474 22006 5502
rect 21902 5469 22034 5474
rect 21798 4937 21826 4942
rect 22078 4858 22106 5614
rect 22232 5110 22364 5115
rect 22260 5082 22284 5110
rect 22312 5082 22336 5110
rect 22232 5077 22364 5082
rect 22078 4825 22106 4830
rect 22414 4802 22442 4807
rect 21902 4718 22034 4723
rect 21930 4690 21954 4718
rect 21982 4690 22006 4718
rect 21902 4685 22034 4690
rect 21966 4634 21994 4639
rect 21966 4578 21994 4606
rect 22414 4634 22442 4774
rect 22414 4601 22442 4606
rect 22190 4578 22218 4583
rect 21966 4550 22190 4578
rect 22190 4545 22218 4550
rect 22232 4326 22364 4331
rect 22260 4298 22284 4326
rect 22312 4298 22336 4326
rect 22232 4293 22364 4298
rect 22414 4242 22442 4247
rect 21902 3934 22034 3939
rect 21930 3906 21954 3934
rect 21982 3906 22006 3934
rect 21902 3901 22034 3906
rect 22232 3542 22364 3547
rect 22260 3514 22284 3542
rect 22312 3514 22336 3542
rect 22232 3509 22364 3514
rect 21686 3402 21714 3407
rect 21630 2617 21658 2623
rect 21630 2591 21631 2617
rect 21657 2591 21658 2617
rect 21630 2506 21658 2591
rect 21630 2473 21658 2478
rect 21518 2143 21519 2169
rect 21545 2143 21546 2169
rect 21518 2137 21546 2143
rect 21686 2058 21714 3374
rect 22414 3178 22442 4214
rect 21902 3150 22034 3155
rect 21930 3122 21954 3150
rect 21982 3122 22006 3150
rect 22414 3145 22442 3150
rect 22526 3234 22554 3239
rect 21902 3117 22034 3122
rect 22526 2953 22554 3206
rect 22526 2927 22527 2953
rect 22553 2927 22554 2953
rect 22526 2921 22554 2927
rect 22582 3122 22610 3127
rect 22134 2786 22162 2791
rect 22134 2674 22162 2758
rect 22232 2758 22364 2763
rect 22260 2730 22284 2758
rect 22312 2730 22336 2758
rect 22232 2725 22364 2730
rect 22190 2674 22218 2679
rect 22134 2673 22218 2674
rect 22134 2647 22191 2673
rect 22217 2647 22218 2673
rect 22134 2646 22218 2647
rect 22190 2641 22218 2646
rect 21798 2561 21826 2567
rect 21798 2535 21799 2561
rect 21825 2535 21826 2561
rect 21686 2025 21714 2030
rect 21742 2225 21770 2231
rect 21742 2199 21743 2225
rect 21769 2199 21770 2225
rect 21462 1751 21463 1777
rect 21489 1751 21490 1777
rect 21462 1745 21490 1751
rect 21238 1409 21266 1414
rect 21406 1722 21434 1727
rect 21294 1330 21322 1335
rect 21294 1283 21322 1302
rect 20790 1273 20818 1279
rect 20790 1247 20791 1273
rect 20817 1247 20818 1273
rect 20790 658 20818 1247
rect 21182 1106 21210 1111
rect 21182 1059 21210 1078
rect 20902 1050 20930 1055
rect 20902 1003 20930 1022
rect 20790 625 20818 630
rect 20958 658 20986 663
rect 20958 56 20986 630
rect 21182 490 21210 495
rect 21182 56 21210 462
rect 21406 56 21434 1694
rect 21574 1329 21602 1335
rect 21574 1303 21575 1329
rect 21601 1303 21602 1329
rect 21574 601 21602 1303
rect 21574 575 21575 601
rect 21601 575 21602 601
rect 21574 569 21602 575
rect 21630 1330 21658 1335
rect 21630 56 21658 1302
rect 21742 993 21770 2199
rect 21798 2226 21826 2535
rect 22470 2562 22498 2567
rect 22470 2515 22498 2534
rect 21902 2366 22034 2371
rect 21930 2338 21954 2366
rect 21982 2338 22006 2366
rect 21902 2333 22034 2338
rect 21798 2193 21826 2198
rect 22232 1974 22364 1979
rect 22260 1946 22284 1974
rect 22312 1946 22336 1974
rect 22232 1941 22364 1946
rect 22302 1778 22330 1783
rect 21798 1722 21826 1741
rect 22302 1731 22330 1750
rect 21798 1689 21826 1694
rect 21902 1582 22034 1587
rect 21930 1554 21954 1582
rect 21982 1554 22006 1582
rect 21902 1549 22034 1554
rect 22582 1385 22610 3094
rect 22638 2394 22666 6454
rect 23534 6425 23562 7014
rect 24094 6874 24122 6879
rect 23534 6399 23535 6425
rect 23561 6399 23562 6425
rect 23534 6393 23562 6399
rect 24038 6481 24066 6487
rect 24038 6455 24039 6481
rect 24065 6455 24066 6481
rect 24038 6146 24066 6455
rect 24038 6113 24066 6118
rect 23534 5642 23562 5647
rect 23534 3570 23562 5614
rect 23534 3537 23562 3542
rect 22694 3402 22722 3407
rect 22694 3290 22722 3374
rect 22694 3257 22722 3262
rect 23422 3066 23450 3071
rect 23422 2953 23450 3038
rect 23422 2927 23423 2953
rect 23449 2927 23450 2953
rect 23422 2921 23450 2927
rect 22806 2897 22834 2903
rect 22806 2871 22807 2897
rect 22833 2871 22834 2897
rect 22638 2361 22666 2366
rect 22694 2674 22722 2679
rect 22582 1359 22583 1385
rect 22609 1359 22610 1385
rect 22582 1353 22610 1359
rect 22638 2226 22666 2231
rect 22302 1330 22330 1335
rect 22302 1283 22330 1302
rect 22470 1330 22498 1335
rect 22232 1190 22364 1195
rect 22260 1162 22284 1190
rect 22312 1162 22336 1190
rect 22232 1157 22364 1162
rect 21742 967 21743 993
rect 21769 967 21770 993
rect 21742 961 21770 967
rect 22414 1050 22442 1055
rect 21966 882 21994 901
rect 21966 849 21994 854
rect 21902 798 22034 803
rect 21930 770 21954 798
rect 21982 770 22006 798
rect 21902 765 22034 770
rect 22078 770 22106 775
rect 21854 546 21882 551
rect 21854 499 21882 518
rect 21854 210 21882 215
rect 21854 56 21882 182
rect 22078 56 22106 742
rect 22358 658 22386 663
rect 22358 611 22386 630
rect 22232 406 22364 411
rect 22260 378 22284 406
rect 22312 378 22336 406
rect 22232 373 22364 378
rect 22302 322 22330 327
rect 22302 56 22330 294
rect 22414 98 22442 1022
rect 22470 714 22498 1302
rect 22470 681 22498 686
rect 22582 994 22610 999
rect 22582 714 22610 966
rect 22582 681 22610 686
rect 22638 490 22666 2198
rect 22694 1050 22722 2646
rect 22694 1017 22722 1022
rect 22750 1721 22778 1727
rect 22750 1695 22751 1721
rect 22777 1695 22778 1721
rect 22694 937 22722 943
rect 22694 911 22695 937
rect 22721 911 22722 937
rect 22694 546 22722 911
rect 22694 513 22722 518
rect 22638 457 22666 462
rect 22750 322 22778 1695
rect 22806 601 22834 2871
rect 23702 2897 23730 2903
rect 23702 2871 23703 2897
rect 23729 2871 23730 2897
rect 23478 2562 23506 2567
rect 23086 1946 23114 1951
rect 23086 1833 23114 1918
rect 23086 1807 23087 1833
rect 23113 1807 23114 1833
rect 23086 1801 23114 1807
rect 23254 1722 23282 1727
rect 22974 1441 23002 1447
rect 22974 1415 22975 1441
rect 23001 1415 23002 1441
rect 22974 770 23002 1415
rect 23086 1050 23114 1055
rect 23086 1003 23114 1022
rect 23254 1049 23282 1694
rect 23478 1385 23506 2534
rect 23478 1359 23479 1385
rect 23505 1359 23506 1385
rect 23478 1353 23506 1359
rect 23590 2225 23618 2231
rect 23590 2199 23591 2225
rect 23617 2199 23618 2225
rect 23254 1023 23255 1049
rect 23281 1023 23282 1049
rect 23254 1017 23282 1023
rect 23478 1162 23506 1167
rect 23422 994 23450 999
rect 22974 737 23002 742
rect 23198 826 23226 831
rect 22806 575 22807 601
rect 22833 575 22834 601
rect 22806 569 22834 575
rect 22974 658 23002 663
rect 22750 289 22778 294
rect 22414 65 22442 70
rect 22526 154 22554 159
rect 22526 56 22554 126
rect 22750 98 22778 103
rect 22750 56 22778 70
rect 22974 56 23002 630
rect 23198 56 23226 798
rect 23422 56 23450 966
rect 23478 993 23506 1134
rect 23478 967 23479 993
rect 23505 967 23506 993
rect 23478 961 23506 967
rect 23590 826 23618 2199
rect 23646 1329 23674 1335
rect 23646 1303 23647 1329
rect 23673 1303 23674 1329
rect 23646 1274 23674 1303
rect 23646 1241 23674 1246
rect 23702 1050 23730 2871
rect 23982 2786 24010 2791
rect 23926 2114 23954 2119
rect 23926 2067 23954 2086
rect 23702 1017 23730 1022
rect 23926 1273 23954 1279
rect 23926 1247 23927 1273
rect 23953 1247 23954 1273
rect 23590 793 23618 798
rect 23646 882 23674 887
rect 23590 545 23618 551
rect 23590 519 23591 545
rect 23617 519 23618 545
rect 23590 210 23618 519
rect 23590 177 23618 182
rect 23646 56 23674 854
rect 23870 770 23898 775
rect 23870 56 23898 742
rect 23926 658 23954 1247
rect 23926 625 23954 630
rect 23982 601 24010 2758
rect 24094 2225 24122 6846
rect 24766 6202 24794 7056
rect 26222 7042 26250 7056
rect 26222 7009 26250 7014
rect 26390 7042 26418 7047
rect 25662 6594 25690 6599
rect 25606 6426 25634 6431
rect 24990 6202 25018 6207
rect 24766 6201 25018 6202
rect 24766 6175 24991 6201
rect 25017 6175 25018 6201
rect 24766 6174 25018 6175
rect 24990 6169 25018 6174
rect 25494 6034 25522 6039
rect 25494 5987 25522 6006
rect 25438 5866 25466 5871
rect 24878 3402 24906 3407
rect 24486 3346 24514 3351
rect 24486 3299 24514 3318
rect 24710 3289 24738 3295
rect 24710 3263 24711 3289
rect 24737 3263 24738 3289
rect 24318 2618 24346 2623
rect 24318 2506 24346 2590
rect 24318 2473 24346 2478
rect 24094 2199 24095 2225
rect 24121 2199 24122 2225
rect 24094 2193 24122 2199
rect 24038 2170 24066 2175
rect 24038 1833 24066 2142
rect 24318 2169 24346 2175
rect 24318 2143 24319 2169
rect 24345 2143 24346 2169
rect 24038 1807 24039 1833
rect 24065 1807 24066 1833
rect 24038 1801 24066 1807
rect 24206 2058 24234 2063
rect 24038 993 24066 999
rect 24038 967 24039 993
rect 24065 967 24066 993
rect 24038 938 24066 967
rect 24038 905 24066 910
rect 23982 575 23983 601
rect 24009 575 24010 601
rect 23982 569 24010 575
rect 24206 546 24234 2030
rect 24318 1722 24346 2143
rect 24710 1778 24738 3263
rect 24822 1890 24850 1895
rect 24822 1833 24850 1862
rect 24822 1807 24823 1833
rect 24849 1807 24850 1833
rect 24822 1801 24850 1807
rect 24710 1745 24738 1750
rect 24318 1689 24346 1694
rect 24374 1721 24402 1727
rect 24374 1695 24375 1721
rect 24401 1695 24402 1721
rect 24206 513 24234 518
rect 24318 938 24346 943
rect 24094 266 24122 271
rect 24094 56 24122 238
rect 24318 56 24346 910
rect 24374 770 24402 1695
rect 24486 1385 24514 1391
rect 24486 1359 24487 1385
rect 24513 1359 24514 1385
rect 24374 737 24402 742
rect 24430 937 24458 943
rect 24430 911 24431 937
rect 24457 911 24458 937
rect 24374 545 24402 551
rect 24374 519 24375 545
rect 24401 519 24402 545
rect 24374 154 24402 519
rect 24374 121 24402 126
rect 24430 98 24458 911
rect 24486 602 24514 1359
rect 24710 1273 24738 1279
rect 24710 1247 24711 1273
rect 24737 1247 24738 1273
rect 24710 994 24738 1247
rect 24710 961 24738 966
rect 24766 1218 24794 1223
rect 24486 569 24514 574
rect 24542 770 24570 775
rect 24430 65 24458 70
rect 24542 56 24570 742
rect 24766 714 24794 1190
rect 24878 993 24906 3374
rect 25102 2954 25130 2959
rect 25102 2169 25130 2926
rect 25438 2953 25466 5838
rect 25438 2927 25439 2953
rect 25465 2927 25466 2953
rect 25438 2921 25466 2927
rect 25494 5698 25522 5703
rect 25102 2143 25103 2169
rect 25129 2143 25130 2169
rect 25102 2137 25130 2143
rect 25326 2282 25354 2287
rect 25270 1721 25298 1727
rect 25270 1695 25271 1721
rect 25297 1695 25298 1721
rect 25214 1386 25242 1391
rect 25214 1339 25242 1358
rect 24878 967 24879 993
rect 24905 967 24906 993
rect 24878 961 24906 967
rect 25214 937 25242 943
rect 25214 911 25215 937
rect 25241 911 25242 937
rect 25214 882 25242 911
rect 25214 849 25242 854
rect 24766 681 24794 686
rect 24990 826 25018 831
rect 24766 602 24794 607
rect 24766 555 24794 574
rect 24766 210 24794 215
rect 24766 56 24794 182
rect 24990 56 25018 798
rect 25270 770 25298 1695
rect 25326 1386 25354 2254
rect 25326 1353 25354 1358
rect 25382 2057 25410 2063
rect 25382 2031 25383 2057
rect 25409 2031 25410 2057
rect 25382 826 25410 2031
rect 25382 793 25410 798
rect 25438 2058 25466 2063
rect 25270 737 25298 742
rect 25438 714 25466 2030
rect 25494 1694 25522 5670
rect 25550 3010 25578 3015
rect 25550 2394 25578 2982
rect 25550 2361 25578 2366
rect 25606 1833 25634 6398
rect 25662 5082 25690 6566
rect 26390 6425 26418 7014
rect 27678 7042 27706 7056
rect 27678 7009 27706 7014
rect 27902 7042 27930 7047
rect 26390 6399 26391 6425
rect 26417 6399 26418 6425
rect 26390 6393 26418 6399
rect 26894 6481 26922 6487
rect 26894 6455 26895 6481
rect 26921 6455 26922 6481
rect 26502 6202 26530 6207
rect 25998 5698 26026 5703
rect 25662 5049 25690 5054
rect 25886 5362 25914 5367
rect 25774 4186 25802 4191
rect 25606 1807 25607 1833
rect 25633 1807 25634 1833
rect 25606 1801 25634 1807
rect 25662 3794 25690 3799
rect 25662 1694 25690 3766
rect 25718 2897 25746 2903
rect 25718 2871 25719 2897
rect 25745 2871 25746 2897
rect 25718 2618 25746 2871
rect 25718 2585 25746 2590
rect 25494 1666 25578 1694
rect 25550 1633 25578 1638
rect 25606 1666 25690 1694
rect 25718 2506 25746 2511
rect 25550 1498 25578 1503
rect 25494 1273 25522 1279
rect 25494 1247 25495 1273
rect 25521 1247 25522 1273
rect 25494 882 25522 1247
rect 25494 849 25522 854
rect 25550 826 25578 1470
rect 25550 793 25578 798
rect 25438 681 25466 686
rect 25382 602 25410 607
rect 25606 602 25634 1666
rect 25382 601 25634 602
rect 25382 575 25383 601
rect 25409 575 25634 601
rect 25382 574 25634 575
rect 25662 1162 25690 1167
rect 25382 569 25410 574
rect 25438 490 25466 495
rect 25214 378 25242 383
rect 25214 56 25242 350
rect 25438 56 25466 462
rect 25550 489 25578 495
rect 25550 463 25551 489
rect 25577 463 25578 489
rect 25550 266 25578 463
rect 25550 233 25578 238
rect 25662 56 25690 1134
rect 25718 993 25746 2478
rect 25774 1610 25802 4158
rect 25886 2506 25914 5334
rect 25942 5138 25970 5143
rect 25942 3290 25970 5110
rect 25998 4690 26026 5670
rect 25998 4657 26026 4662
rect 26278 5082 26306 5087
rect 25942 3257 25970 3262
rect 26166 4578 26194 4583
rect 25886 2473 25914 2478
rect 26110 3178 26138 3183
rect 25886 1777 25914 1783
rect 25886 1751 25887 1777
rect 25913 1751 25914 1777
rect 25774 1577 25802 1582
rect 25830 1722 25858 1727
rect 25718 967 25719 993
rect 25745 967 25746 993
rect 25718 961 25746 967
rect 25830 770 25858 1694
rect 25886 1694 25914 1751
rect 25886 1666 26082 1694
rect 25886 938 25914 943
rect 25886 891 25914 910
rect 25830 742 25914 770
rect 25886 56 25914 742
rect 26054 658 26082 1666
rect 26110 1441 26138 3150
rect 26110 1415 26111 1441
rect 26137 1415 26138 1441
rect 26110 1409 26138 1415
rect 26054 630 26138 658
rect 26110 56 26138 630
rect 26166 601 26194 4550
rect 26166 575 26167 601
rect 26193 575 26194 601
rect 26166 569 26194 575
rect 26222 2338 26250 2343
rect 26222 546 26250 2310
rect 26222 513 26250 518
rect 26278 378 26306 5054
rect 26502 1694 26530 6174
rect 26838 6090 26866 6095
rect 26558 5922 26586 5927
rect 26558 5026 26586 5894
rect 26558 4993 26586 4998
rect 26726 5810 26754 5815
rect 26726 2338 26754 5782
rect 26838 3234 26866 6062
rect 26894 5138 26922 6455
rect 27902 6425 27930 7014
rect 29134 7042 29162 7056
rect 29134 7009 29162 7014
rect 29358 7042 29386 7047
rect 28406 6482 28434 6487
rect 28406 6435 28434 6454
rect 27902 6399 27903 6425
rect 27929 6399 27930 6425
rect 27902 6393 27930 6399
rect 29358 6425 29386 7014
rect 30590 6594 30618 7056
rect 31318 6986 31346 6991
rect 30590 6561 30618 6566
rect 31150 6762 31178 6767
rect 31094 6538 31122 6543
rect 29358 6399 29359 6425
rect 29385 6399 29386 6425
rect 29358 6393 29386 6399
rect 29750 6481 29778 6487
rect 29750 6455 29751 6481
rect 29777 6455 29778 6481
rect 29526 6314 29554 6319
rect 29526 6201 29554 6286
rect 29526 6175 29527 6201
rect 29553 6175 29554 6201
rect 29526 6169 29554 6175
rect 28462 6146 28490 6151
rect 27566 6034 27594 6039
rect 27566 5987 27594 6006
rect 27734 6034 27762 6039
rect 26894 5105 26922 5110
rect 27678 5866 27706 5871
rect 27678 4186 27706 5838
rect 27734 5306 27762 6006
rect 27734 5273 27762 5278
rect 27846 5977 27874 5983
rect 27846 5951 27847 5977
rect 27873 5951 27874 5977
rect 27846 5082 27874 5951
rect 27846 5049 27874 5054
rect 27678 4158 27762 4186
rect 27678 3738 27706 3743
rect 26838 3201 26866 3206
rect 27622 3570 27650 3575
rect 27062 2897 27090 2903
rect 27062 2871 27063 2897
rect 27089 2871 27090 2897
rect 26782 2842 26810 2847
rect 26782 2795 26810 2814
rect 27062 2786 27090 2871
rect 27062 2753 27090 2758
rect 27398 2674 27426 2679
rect 27398 2627 27426 2646
rect 27622 2618 27650 3542
rect 27678 3346 27706 3710
rect 27678 3313 27706 3318
rect 27622 2585 27650 2590
rect 27678 2562 27706 2567
rect 27678 2515 27706 2534
rect 26726 2305 26754 2310
rect 26950 2506 26978 2511
rect 26502 1666 26586 1694
rect 26446 1330 26474 1335
rect 26390 1273 26418 1279
rect 26390 1247 26391 1273
rect 26417 1247 26418 1273
rect 26390 1162 26418 1247
rect 26390 1129 26418 1134
rect 26446 993 26474 1302
rect 26446 967 26447 993
rect 26473 967 26474 993
rect 26446 961 26474 967
rect 26446 545 26474 551
rect 26446 519 26447 545
rect 26473 519 26474 545
rect 26278 350 26362 378
rect 26334 56 26362 350
rect 26446 210 26474 519
rect 26446 177 26474 182
rect 26558 56 26586 1666
rect 26726 1442 26754 1447
rect 26726 1395 26754 1414
rect 26950 1162 26978 2478
rect 27734 2170 27762 4158
rect 27734 2137 27762 2142
rect 27790 3234 27818 3239
rect 27790 1834 27818 3206
rect 28070 2394 28098 2399
rect 27790 1801 27818 1806
rect 27958 2002 27986 2007
rect 27958 1833 27986 1974
rect 27958 1807 27959 1833
rect 27985 1807 27986 1833
rect 27958 1801 27986 1807
rect 27230 1666 27258 1671
rect 27006 1274 27034 1279
rect 27006 1227 27034 1246
rect 26950 1134 27034 1162
rect 26670 881 26698 887
rect 26670 855 26671 881
rect 26697 855 26698 881
rect 26670 378 26698 855
rect 26670 345 26698 350
rect 26782 490 26810 495
rect 26782 56 26810 462
rect 27006 56 27034 1134
rect 27230 56 27258 1638
rect 28070 1666 28098 2366
rect 28462 1833 28490 6118
rect 29022 6034 29050 6039
rect 29022 5987 29050 6006
rect 29358 5697 29386 5703
rect 29358 5671 29359 5697
rect 29385 5671 29386 5697
rect 29022 5082 29050 5087
rect 28462 1807 28463 1833
rect 28489 1807 28490 1833
rect 28462 1801 28490 1807
rect 28518 2114 28546 2119
rect 28238 1778 28266 1783
rect 28238 1731 28266 1750
rect 28070 1633 28098 1638
rect 27678 1610 27706 1615
rect 27454 322 27482 327
rect 27454 56 27482 294
rect 27678 56 27706 1582
rect 28350 1274 28378 1279
rect 28126 1162 28154 1167
rect 27902 882 27930 887
rect 27902 56 27930 854
rect 28126 56 28154 1134
rect 28350 56 28378 1246
rect 28518 1050 28546 2086
rect 28518 1017 28546 1022
rect 28574 1778 28602 1783
rect 28574 56 28602 1750
rect 28742 1777 28770 1783
rect 28742 1751 28743 1777
rect 28769 1751 28770 1777
rect 28742 1694 28770 1751
rect 28742 1666 28826 1694
rect 28798 56 28826 1666
rect 29022 56 29050 5054
rect 29358 4522 29386 5671
rect 29358 4489 29386 4494
rect 29582 5138 29610 5143
rect 29414 4018 29442 4023
rect 29414 3737 29442 3990
rect 29414 3711 29415 3737
rect 29441 3711 29442 3737
rect 29414 3705 29442 3711
rect 29582 2225 29610 5110
rect 29582 2199 29583 2225
rect 29609 2199 29610 2225
rect 29582 2193 29610 2199
rect 29638 3681 29666 3687
rect 29638 3655 29639 3681
rect 29665 3655 29666 3681
rect 29414 2169 29442 2175
rect 29414 2143 29415 2169
rect 29441 2143 29442 2169
rect 29414 1498 29442 2143
rect 29638 1890 29666 3655
rect 29638 1857 29666 1862
rect 29750 1694 29778 6455
rect 30086 6481 30114 6487
rect 30086 6455 30087 6481
rect 30113 6455 30114 6481
rect 30086 5922 30114 6455
rect 30814 6482 30842 6487
rect 30254 6370 30282 6375
rect 30254 6089 30282 6342
rect 30254 6063 30255 6089
rect 30281 6063 30282 6089
rect 30254 6057 30282 6063
rect 30590 6369 30618 6375
rect 30590 6343 30591 6369
rect 30617 6343 30618 6369
rect 30590 6090 30618 6343
rect 30590 6057 30618 6062
rect 30758 6145 30786 6151
rect 30758 6119 30759 6145
rect 30785 6119 30786 6145
rect 30086 5889 30114 5894
rect 30758 5922 30786 6119
rect 30758 5889 30786 5894
rect 29862 5754 29890 5759
rect 29862 5641 29890 5726
rect 30142 5698 30170 5703
rect 30142 5651 30170 5670
rect 29862 5615 29863 5641
rect 29889 5615 29890 5641
rect 29862 5609 29890 5615
rect 30646 5642 30674 5647
rect 30646 5595 30674 5614
rect 30254 5249 30282 5255
rect 30254 5223 30255 5249
rect 30281 5223 30282 5249
rect 30254 5194 30282 5223
rect 30254 5161 30282 5166
rect 30646 5249 30674 5255
rect 30646 5223 30647 5249
rect 30673 5223 30674 5249
rect 30646 5194 30674 5223
rect 30646 5161 30674 5166
rect 30534 4970 30562 4975
rect 30534 4923 30562 4942
rect 30142 4914 30170 4919
rect 30142 4867 30170 4886
rect 30254 4802 30282 4807
rect 30254 4521 30282 4774
rect 30758 4634 30786 4639
rect 30758 4587 30786 4606
rect 30254 4495 30255 4521
rect 30281 4495 30282 4521
rect 30254 4489 30282 4495
rect 30478 4130 30506 4135
rect 30478 4083 30506 4102
rect 30702 4073 30730 4079
rect 30702 4047 30703 4073
rect 30729 4047 30730 4073
rect 30254 3682 30282 3687
rect 30254 3635 30282 3654
rect 30142 3345 30170 3351
rect 30142 3319 30143 3345
rect 30169 3319 30170 3345
rect 30142 3290 30170 3319
rect 30142 3257 30170 3262
rect 30646 3233 30674 3239
rect 30646 3207 30647 3233
rect 30673 3207 30674 3233
rect 30646 2954 30674 3207
rect 30646 2921 30674 2926
rect 30590 2841 30618 2847
rect 30590 2815 30591 2841
rect 30617 2815 30618 2841
rect 30142 2730 30170 2735
rect 30142 2617 30170 2702
rect 30142 2591 30143 2617
rect 30169 2591 30170 2617
rect 30142 2585 30170 2591
rect 30534 2562 30562 2567
rect 30534 2515 30562 2534
rect 30254 2170 30282 2175
rect 30254 2123 30282 2142
rect 30142 1834 30170 1839
rect 30142 1787 30170 1806
rect 29302 1470 29442 1498
rect 29526 1666 29778 1694
rect 29190 1162 29218 1167
rect 29190 1049 29218 1134
rect 29190 1023 29191 1049
rect 29217 1023 29218 1049
rect 29190 1017 29218 1023
rect 29302 826 29330 1470
rect 29358 1330 29386 1335
rect 29526 1330 29554 1666
rect 30254 1386 30282 1391
rect 30254 1339 30282 1358
rect 29358 1329 29554 1330
rect 29358 1303 29359 1329
rect 29385 1303 29554 1329
rect 29358 1302 29554 1303
rect 29358 1297 29386 1302
rect 29638 1274 29666 1279
rect 29638 1273 29722 1274
rect 29638 1247 29639 1273
rect 29665 1247 29722 1273
rect 29638 1246 29722 1247
rect 29638 1241 29666 1246
rect 29582 1218 29610 1223
rect 29582 1106 29610 1190
rect 29638 1106 29666 1111
rect 29582 1105 29666 1106
rect 29582 1079 29639 1105
rect 29665 1079 29666 1105
rect 29582 1078 29666 1079
rect 29638 1073 29666 1078
rect 29246 798 29330 826
rect 29470 993 29498 999
rect 29470 967 29471 993
rect 29497 967 29498 993
rect 29246 56 29274 798
rect 29302 714 29330 719
rect 29302 601 29330 686
rect 29302 575 29303 601
rect 29329 575 29330 601
rect 29302 569 29330 575
rect 29470 490 29498 967
rect 29470 457 29498 462
rect 29526 770 29554 775
rect 29526 378 29554 742
rect 29470 350 29554 378
rect 29470 56 29498 350
rect 29694 56 29722 1246
rect 29918 1050 29946 1055
rect 29918 1003 29946 1022
rect 30142 993 30170 999
rect 30142 967 30143 993
rect 30169 967 30170 993
rect 30142 826 30170 967
rect 30142 793 30170 798
rect 30590 770 30618 2815
rect 30646 2113 30674 2119
rect 30646 2087 30647 2113
rect 30673 2087 30674 2113
rect 30646 1834 30674 2087
rect 30646 1801 30674 1806
rect 30646 1722 30674 1741
rect 30646 1689 30674 1694
rect 30646 1330 30674 1335
rect 30646 1283 30674 1302
rect 30646 882 30674 887
rect 30646 835 30674 854
rect 30590 737 30618 742
rect 29806 657 29834 663
rect 29806 631 29807 657
rect 29833 631 29834 657
rect 29806 266 29834 631
rect 30590 657 30618 663
rect 30590 631 30591 657
rect 30617 631 30618 657
rect 30086 545 30114 551
rect 30086 519 30087 545
rect 30113 519 30114 545
rect 29806 233 29834 238
rect 29918 490 29946 495
rect 29918 56 29946 462
rect 30086 434 30114 519
rect 30590 490 30618 631
rect 30702 602 30730 4047
rect 30758 3793 30786 3799
rect 30758 3767 30759 3793
rect 30785 3767 30786 3793
rect 30758 3402 30786 3767
rect 30758 3369 30786 3374
rect 30814 3009 30842 6454
rect 30982 6481 31010 6487
rect 30982 6455 30983 6481
rect 31009 6455 31010 6481
rect 30926 5697 30954 5703
rect 30926 5671 30927 5697
rect 30953 5671 30954 5697
rect 30926 5418 30954 5671
rect 30926 5385 30954 5390
rect 30926 4913 30954 4919
rect 30926 4887 30927 4913
rect 30953 4887 30954 4913
rect 30926 4858 30954 4887
rect 30926 4825 30954 4830
rect 30926 4129 30954 4135
rect 30926 4103 30927 4129
rect 30953 4103 30954 4129
rect 30926 4074 30954 4103
rect 30926 4041 30954 4046
rect 30926 3346 30954 3351
rect 30926 3299 30954 3318
rect 30814 2983 30815 3009
rect 30841 2983 30842 3009
rect 30814 2977 30842 2983
rect 30926 2618 30954 2623
rect 30926 2571 30954 2590
rect 30926 2338 30954 2343
rect 30926 1833 30954 2310
rect 30926 1807 30927 1833
rect 30953 1807 30954 1833
rect 30926 1801 30954 1807
rect 30926 1666 30954 1671
rect 30926 1049 30954 1638
rect 30982 1162 31010 6455
rect 31038 6033 31066 6039
rect 31038 6007 31039 6033
rect 31065 6007 31066 6033
rect 31038 5138 31066 6007
rect 31094 5754 31122 6510
rect 31094 5721 31122 5726
rect 31094 5305 31122 5311
rect 31094 5279 31095 5305
rect 31121 5279 31122 5305
rect 31094 5250 31122 5279
rect 31094 5217 31122 5222
rect 31038 5110 31122 5138
rect 31094 4690 31122 5110
rect 31150 4970 31178 6734
rect 31262 6594 31290 6599
rect 31262 6547 31290 6566
rect 31150 4937 31178 4942
rect 31094 4657 31122 4662
rect 31318 4634 31346 6958
rect 31542 6145 31570 6151
rect 31542 6119 31543 6145
rect 31569 6119 31570 6145
rect 31374 5641 31402 5647
rect 31374 5615 31375 5641
rect 31401 5615 31402 5641
rect 31374 4970 31402 5615
rect 31542 5418 31570 6119
rect 31542 5385 31570 5390
rect 31374 4937 31402 4942
rect 31430 5249 31458 5255
rect 31430 5223 31431 5249
rect 31457 5223 31458 5249
rect 31318 4601 31346 4606
rect 31374 4857 31402 4863
rect 31374 4831 31375 4857
rect 31401 4831 31402 4857
rect 31094 4521 31122 4527
rect 31094 4495 31095 4521
rect 31121 4495 31122 4521
rect 31094 4410 31122 4495
rect 31374 4522 31402 4831
rect 31430 4746 31458 5223
rect 31430 4713 31458 4718
rect 31374 4489 31402 4494
rect 31094 4377 31122 4382
rect 31430 4465 31458 4471
rect 31430 4439 31431 4465
rect 31457 4439 31458 4465
rect 31430 4298 31458 4439
rect 31430 4265 31458 4270
rect 31542 4074 31570 4079
rect 31430 4017 31458 4023
rect 31430 3991 31431 4017
rect 31457 3991 31458 4017
rect 31094 3962 31122 3967
rect 31094 3737 31122 3934
rect 31430 3850 31458 3991
rect 31430 3817 31458 3822
rect 31542 3849 31570 4046
rect 31542 3823 31543 3849
rect 31569 3823 31570 3849
rect 31542 3817 31570 3823
rect 31094 3711 31095 3737
rect 31121 3711 31122 3737
rect 31094 3705 31122 3711
rect 31430 3626 31458 3631
rect 31430 3289 31458 3598
rect 31430 3263 31431 3289
rect 31457 3263 31458 3289
rect 31430 3257 31458 3263
rect 31542 3178 31570 3183
rect 31542 3065 31570 3150
rect 31542 3039 31543 3065
rect 31569 3039 31570 3065
rect 31542 3033 31570 3039
rect 31094 2953 31122 2959
rect 31094 2927 31095 2953
rect 31121 2927 31122 2953
rect 31094 2898 31122 2927
rect 31094 2865 31122 2870
rect 31318 2730 31346 2735
rect 31318 2617 31346 2702
rect 31318 2591 31319 2617
rect 31345 2591 31346 2617
rect 31318 2585 31346 2591
rect 31262 2562 31290 2567
rect 31094 2450 31122 2455
rect 31094 2169 31122 2422
rect 31262 2282 31290 2534
rect 31262 2249 31290 2254
rect 31542 2506 31570 2511
rect 31542 2281 31570 2478
rect 31542 2255 31543 2281
rect 31569 2255 31570 2281
rect 31542 2249 31570 2255
rect 31094 2143 31095 2169
rect 31121 2143 31122 2169
rect 31094 2137 31122 2143
rect 31430 2058 31458 2063
rect 31318 1722 31346 1727
rect 30982 1129 31010 1134
rect 31094 1385 31122 1391
rect 31094 1359 31095 1385
rect 31121 1359 31122 1385
rect 31094 1106 31122 1359
rect 31318 1386 31346 1694
rect 31430 1721 31458 2030
rect 31430 1695 31431 1721
rect 31457 1695 31458 1721
rect 31430 1689 31458 1695
rect 31542 1610 31570 1615
rect 31542 1497 31570 1582
rect 31542 1471 31543 1497
rect 31569 1471 31570 1497
rect 31542 1465 31570 1471
rect 31318 1353 31346 1358
rect 31094 1073 31122 1078
rect 31374 1330 31402 1335
rect 30926 1023 30927 1049
rect 30953 1023 30954 1049
rect 30926 1017 30954 1023
rect 30702 569 30730 574
rect 31094 601 31122 607
rect 31094 575 31095 601
rect 31121 575 31122 601
rect 31094 546 31122 575
rect 31094 513 31122 518
rect 30590 457 30618 462
rect 30086 401 30114 406
rect 2128 0 2184 56
rect 2352 0 2408 56
rect 2576 0 2632 56
rect 2800 0 2856 56
rect 3024 0 3080 56
rect 3248 0 3304 56
rect 3472 0 3528 56
rect 3696 0 3752 56
rect 3920 0 3976 56
rect 4144 0 4200 56
rect 4368 0 4424 56
rect 4592 0 4648 56
rect 4816 0 4872 56
rect 5040 0 5096 56
rect 5264 0 5320 56
rect 5488 0 5544 56
rect 5712 0 5768 56
rect 5936 0 5992 56
rect 6160 0 6216 56
rect 6384 0 6440 56
rect 6608 0 6664 56
rect 6832 0 6888 56
rect 7056 0 7112 56
rect 7280 0 7336 56
rect 7504 0 7560 56
rect 7728 0 7784 56
rect 7952 0 8008 56
rect 8176 0 8232 56
rect 8400 0 8456 56
rect 8624 0 8680 56
rect 8848 0 8904 56
rect 9072 0 9128 56
rect 9296 0 9352 56
rect 9520 0 9576 56
rect 9744 0 9800 56
rect 9968 0 10024 56
rect 10192 0 10248 56
rect 10416 0 10472 56
rect 10640 0 10696 56
rect 10864 0 10920 56
rect 11088 0 11144 56
rect 11312 0 11368 56
rect 11536 0 11592 56
rect 11760 0 11816 56
rect 11984 0 12040 56
rect 12208 0 12264 56
rect 12432 0 12488 56
rect 12656 0 12712 56
rect 12880 0 12936 56
rect 13104 0 13160 56
rect 13328 0 13384 56
rect 13552 0 13608 56
rect 13776 0 13832 56
rect 14000 0 14056 56
rect 14224 0 14280 56
rect 14448 0 14504 56
rect 14672 0 14728 56
rect 14896 0 14952 56
rect 15120 0 15176 56
rect 15344 0 15400 56
rect 15568 0 15624 56
rect 15792 0 15848 56
rect 16016 0 16072 56
rect 16240 0 16296 56
rect 16464 0 16520 56
rect 16688 0 16744 56
rect 16912 0 16968 56
rect 17136 0 17192 56
rect 17360 0 17416 56
rect 17584 0 17640 56
rect 17808 0 17864 56
rect 18032 0 18088 56
rect 18256 0 18312 56
rect 18480 0 18536 56
rect 18704 0 18760 56
rect 18928 0 18984 56
rect 19152 0 19208 56
rect 19376 0 19432 56
rect 19600 0 19656 56
rect 19824 0 19880 56
rect 20048 0 20104 56
rect 20272 0 20328 56
rect 20496 0 20552 56
rect 20720 0 20776 56
rect 20944 0 21000 56
rect 21168 0 21224 56
rect 21392 0 21448 56
rect 21616 0 21672 56
rect 21840 0 21896 56
rect 22064 0 22120 56
rect 22288 0 22344 56
rect 22512 0 22568 56
rect 22736 0 22792 56
rect 22960 0 23016 56
rect 23184 0 23240 56
rect 23408 0 23464 56
rect 23632 0 23688 56
rect 23856 0 23912 56
rect 24080 0 24136 56
rect 24304 0 24360 56
rect 24528 0 24584 56
rect 24752 0 24808 56
rect 24976 0 25032 56
rect 25200 0 25256 56
rect 25424 0 25480 56
rect 25648 0 25704 56
rect 25872 0 25928 56
rect 26096 0 26152 56
rect 26320 0 26376 56
rect 26544 0 26600 56
rect 26768 0 26824 56
rect 26992 0 27048 56
rect 27216 0 27272 56
rect 27440 0 27496 56
rect 27664 0 27720 56
rect 27888 0 27944 56
rect 28112 0 28168 56
rect 28336 0 28392 56
rect 28560 0 28616 56
rect 28784 0 28840 56
rect 29008 0 29064 56
rect 29232 0 29288 56
rect 29456 0 29512 56
rect 29680 0 29736 56
rect 29904 0 29960 56
rect 31374 42 31402 1302
rect 31430 1162 31458 1167
rect 31430 937 31458 1134
rect 31430 911 31431 937
rect 31457 911 31458 937
rect 31430 905 31458 911
rect 31542 938 31570 943
rect 31542 713 31570 910
rect 31542 687 31543 713
rect 31569 687 31570 713
rect 31542 681 31570 687
rect 31374 9 31402 14
<< via2 >>
rect 910 6958 938 6986
rect 798 6734 826 6762
rect 2926 7014 2954 7042
rect 3150 7014 3178 7042
rect 2232 6677 2260 6678
rect 2232 6651 2233 6677
rect 2233 6651 2259 6677
rect 2259 6651 2260 6677
rect 2232 6650 2260 6651
rect 2284 6677 2312 6678
rect 2284 6651 2285 6677
rect 2285 6651 2311 6677
rect 2311 6651 2312 6677
rect 2284 6650 2312 6651
rect 2336 6677 2364 6678
rect 2336 6651 2337 6677
rect 2337 6651 2363 6677
rect 2363 6651 2364 6677
rect 2336 6650 2364 6651
rect 1750 6481 1778 6482
rect 1750 6455 1751 6481
rect 1751 6455 1777 6481
rect 1777 6455 1778 6481
rect 1750 6454 1778 6455
rect 4382 7014 4410 7042
rect 4606 7014 4634 7042
rect 3822 6734 3850 6762
rect 3654 6342 3682 6370
rect 1902 6285 1930 6286
rect 1902 6259 1903 6285
rect 1903 6259 1929 6285
rect 1929 6259 1930 6285
rect 1902 6258 1930 6259
rect 1954 6285 1982 6286
rect 1954 6259 1955 6285
rect 1955 6259 1981 6285
rect 1981 6259 1982 6285
rect 1954 6258 1982 6259
rect 2006 6285 2034 6286
rect 2006 6259 2007 6285
rect 2007 6259 2033 6285
rect 2033 6259 2034 6285
rect 2006 6258 2034 6259
rect 2232 5893 2260 5894
rect 2232 5867 2233 5893
rect 2233 5867 2259 5893
rect 2259 5867 2260 5893
rect 2232 5866 2260 5867
rect 2284 5893 2312 5894
rect 2284 5867 2285 5893
rect 2285 5867 2311 5893
rect 2311 5867 2312 5893
rect 2284 5866 2312 5867
rect 2336 5893 2364 5894
rect 2336 5867 2337 5893
rect 2337 5867 2363 5893
rect 2363 5867 2364 5893
rect 2336 5866 2364 5867
rect 910 5782 938 5810
rect 798 5670 826 5698
rect 1902 5501 1930 5502
rect 1902 5475 1903 5501
rect 1903 5475 1929 5501
rect 1929 5475 1930 5501
rect 1902 5474 1930 5475
rect 1954 5501 1982 5502
rect 1954 5475 1955 5501
rect 1955 5475 1981 5501
rect 1981 5475 1982 5501
rect 1954 5474 1982 5475
rect 2006 5501 2034 5502
rect 2006 5475 2007 5501
rect 2007 5475 2033 5501
rect 2033 5475 2034 5501
rect 2006 5474 2034 5475
rect 2814 5278 2842 5306
rect 2232 5109 2260 5110
rect 2232 5083 2233 5109
rect 2233 5083 2259 5109
rect 2259 5083 2260 5109
rect 2232 5082 2260 5083
rect 2284 5109 2312 5110
rect 2284 5083 2285 5109
rect 2285 5083 2311 5109
rect 2311 5083 2312 5109
rect 2284 5082 2312 5083
rect 2336 5109 2364 5110
rect 2336 5083 2337 5109
rect 2337 5083 2363 5109
rect 2363 5083 2364 5109
rect 2336 5082 2364 5083
rect 1902 4717 1930 4718
rect 1902 4691 1903 4717
rect 1903 4691 1929 4717
rect 1929 4691 1930 4717
rect 1902 4690 1930 4691
rect 1954 4717 1982 4718
rect 1954 4691 1955 4717
rect 1955 4691 1981 4717
rect 1981 4691 1982 4717
rect 1954 4690 1982 4691
rect 2006 4717 2034 4718
rect 2006 4691 2007 4717
rect 2007 4691 2033 4717
rect 2033 4691 2034 4717
rect 2006 4690 2034 4691
rect 966 4465 994 4466
rect 966 4439 967 4465
rect 967 4439 993 4465
rect 993 4439 994 4465
rect 966 4438 994 4439
rect 1246 4409 1274 4410
rect 1246 4383 1247 4409
rect 1247 4383 1273 4409
rect 1273 4383 1274 4409
rect 1246 4382 1274 4383
rect 2232 4325 2260 4326
rect 2232 4299 2233 4325
rect 2233 4299 2259 4325
rect 2259 4299 2260 4325
rect 2232 4298 2260 4299
rect 2284 4325 2312 4326
rect 2284 4299 2285 4325
rect 2285 4299 2311 4325
rect 2311 4299 2312 4325
rect 2284 4298 2312 4299
rect 2336 4325 2364 4326
rect 2336 4299 2337 4325
rect 2337 4299 2363 4325
rect 2363 4299 2364 4325
rect 2336 4298 2364 4299
rect 1526 3990 1554 4018
rect 350 3038 378 3066
rect 1902 3933 1930 3934
rect 1902 3907 1903 3933
rect 1903 3907 1929 3933
rect 1929 3907 1930 3933
rect 1902 3906 1930 3907
rect 1954 3933 1982 3934
rect 1954 3907 1955 3933
rect 1955 3907 1981 3933
rect 1981 3907 1982 3933
rect 1954 3906 1982 3907
rect 2006 3933 2034 3934
rect 2006 3907 2007 3933
rect 2007 3907 2033 3933
rect 2033 3907 2034 3933
rect 2006 3906 2034 3907
rect 1526 2702 1554 2730
rect 1638 3766 1666 3794
rect 910 2617 938 2618
rect 910 2591 911 2617
rect 911 2591 937 2617
rect 937 2591 938 2617
rect 910 2590 938 2591
rect 1190 2561 1218 2562
rect 1190 2535 1191 2561
rect 1191 2535 1217 2561
rect 1217 2535 1218 2561
rect 1190 2534 1218 2535
rect 1022 2142 1050 2170
rect 350 1358 378 1386
rect 854 1750 882 1778
rect 910 1329 938 1330
rect 910 1303 911 1329
rect 911 1303 937 1329
rect 937 1303 938 1329
rect 910 1302 938 1303
rect 854 910 882 938
rect 966 937 994 938
rect 966 911 967 937
rect 967 911 993 937
rect 993 911 994 937
rect 966 910 994 911
rect 1190 1273 1218 1274
rect 1190 1247 1191 1273
rect 1191 1247 1217 1273
rect 1217 1247 1218 1273
rect 1190 1246 1218 1247
rect 2232 3541 2260 3542
rect 2232 3515 2233 3541
rect 2233 3515 2259 3541
rect 2259 3515 2260 3541
rect 2232 3514 2260 3515
rect 2284 3541 2312 3542
rect 2284 3515 2285 3541
rect 2285 3515 2311 3541
rect 2311 3515 2312 3541
rect 2284 3514 2312 3515
rect 2336 3541 2364 3542
rect 2336 3515 2337 3541
rect 2337 3515 2363 3541
rect 2363 3515 2364 3541
rect 2336 3514 2364 3515
rect 1902 3149 1930 3150
rect 1902 3123 1903 3149
rect 1903 3123 1929 3149
rect 1929 3123 1930 3149
rect 1902 3122 1930 3123
rect 1954 3149 1982 3150
rect 1954 3123 1955 3149
rect 1955 3123 1981 3149
rect 1981 3123 1982 3149
rect 1954 3122 1982 3123
rect 2006 3149 2034 3150
rect 2006 3123 2007 3149
rect 2007 3123 2033 3149
rect 2033 3123 2034 3149
rect 2006 3122 2034 3123
rect 2646 2870 2674 2898
rect 2422 2814 2450 2842
rect 2232 2757 2260 2758
rect 2232 2731 2233 2757
rect 2233 2731 2259 2757
rect 2259 2731 2260 2757
rect 2232 2730 2260 2731
rect 2284 2757 2312 2758
rect 2284 2731 2285 2757
rect 2285 2731 2311 2757
rect 2311 2731 2312 2757
rect 2284 2730 2312 2731
rect 2336 2757 2364 2758
rect 2336 2731 2337 2757
rect 2337 2731 2363 2757
rect 2363 2731 2364 2757
rect 2336 2730 2364 2731
rect 2534 2422 2562 2450
rect 1902 2365 1930 2366
rect 1902 2339 1903 2365
rect 1903 2339 1929 2365
rect 1929 2339 1930 2365
rect 1902 2338 1930 2339
rect 1954 2365 1982 2366
rect 1954 2339 1955 2365
rect 1955 2339 1981 2365
rect 1981 2339 1982 2365
rect 1954 2338 1982 2339
rect 2006 2365 2034 2366
rect 2006 2339 2007 2365
rect 2007 2339 2033 2365
rect 2033 2339 2034 2365
rect 2006 2338 2034 2339
rect 2086 2086 2114 2114
rect 1902 1581 1930 1582
rect 1902 1555 1903 1581
rect 1903 1555 1929 1581
rect 1929 1555 1930 1581
rect 1902 1554 1930 1555
rect 1954 1581 1982 1582
rect 1954 1555 1955 1581
rect 1955 1555 1981 1581
rect 1981 1555 1982 1581
rect 1954 1554 1982 1555
rect 2006 1581 2034 1582
rect 2006 1555 2007 1581
rect 2007 1555 2033 1581
rect 2033 1555 2034 1581
rect 2006 1554 2034 1555
rect 1638 1134 1666 1162
rect 1022 854 1050 882
rect 1902 797 1930 798
rect 1902 771 1903 797
rect 1903 771 1929 797
rect 1929 771 1930 797
rect 1902 770 1930 771
rect 1954 797 1982 798
rect 1954 771 1955 797
rect 1955 771 1981 797
rect 1981 771 1982 797
rect 1954 770 1982 771
rect 2006 797 2034 798
rect 2006 771 2007 797
rect 2007 771 2033 797
rect 2033 771 2034 797
rect 2006 770 2034 771
rect 2232 1973 2260 1974
rect 2232 1947 2233 1973
rect 2233 1947 2259 1973
rect 2259 1947 2260 1973
rect 2232 1946 2260 1947
rect 2284 1973 2312 1974
rect 2284 1947 2285 1973
rect 2285 1947 2311 1973
rect 2311 1947 2312 1973
rect 2284 1946 2312 1947
rect 2336 1973 2364 1974
rect 2336 1947 2337 1973
rect 2337 1947 2363 1973
rect 2363 1947 2364 1973
rect 2336 1946 2364 1947
rect 2814 2030 2842 2058
rect 2926 3542 2954 3570
rect 2534 1470 2562 1498
rect 2534 1358 2562 1386
rect 2232 1189 2260 1190
rect 2232 1163 2233 1189
rect 2233 1163 2259 1189
rect 2259 1163 2260 1189
rect 2232 1162 2260 1163
rect 2284 1189 2312 1190
rect 2284 1163 2285 1189
rect 2285 1163 2311 1189
rect 2311 1163 2312 1189
rect 2284 1162 2312 1163
rect 2336 1189 2364 1190
rect 2336 1163 2337 1189
rect 2337 1163 2363 1189
rect 2363 1163 2364 1189
rect 2336 1162 2364 1163
rect 2366 1078 2394 1106
rect 2086 462 2114 490
rect 2232 405 2260 406
rect 2232 379 2233 405
rect 2233 379 2259 405
rect 2259 379 2260 405
rect 2232 378 2260 379
rect 2284 405 2312 406
rect 2284 379 2285 405
rect 2285 379 2311 405
rect 2311 379 2312 405
rect 2284 378 2312 379
rect 2336 405 2364 406
rect 2336 379 2337 405
rect 2337 379 2363 405
rect 2363 379 2364 405
rect 2336 378 2364 379
rect 2366 294 2394 322
rect 1190 126 1218 154
rect 2142 182 2170 210
rect 2534 238 2562 266
rect 2590 798 2618 826
rect 2646 574 2674 602
rect 5110 6846 5138 6874
rect 7294 7014 7322 7042
rect 7518 7014 7546 7042
rect 6734 6622 6762 6650
rect 5838 6510 5866 6538
rect 6454 6537 6482 6538
rect 6454 6511 6455 6537
rect 6455 6511 6481 6537
rect 6481 6511 6482 6537
rect 6454 6510 6482 6511
rect 5838 6174 5866 6202
rect 5446 5894 5474 5922
rect 4214 5110 4242 5138
rect 4158 4913 4186 4914
rect 4158 4887 4159 4913
rect 4159 4887 4185 4913
rect 4185 4887 4186 4913
rect 4158 4886 4186 4887
rect 3934 4857 3962 4858
rect 3934 4831 3935 4857
rect 3935 4831 3961 4857
rect 3961 4831 3962 4857
rect 3934 4830 3962 4831
rect 4214 3990 4242 4018
rect 4270 4718 4298 4746
rect 3822 2422 3850 2450
rect 3934 3318 3962 3346
rect 3486 1862 3514 1890
rect 3262 1526 3290 1554
rect 2926 294 2954 322
rect 3038 294 3066 322
rect 2814 238 2842 266
rect 3710 1806 3738 1834
rect 4438 3737 4466 3738
rect 4438 3711 4439 3737
rect 4439 3711 4465 3737
rect 4465 3711 4466 3737
rect 4438 3710 4466 3711
rect 4718 3486 4746 3514
rect 4830 3374 4858 3402
rect 4270 3038 4298 3066
rect 4606 3094 4634 3122
rect 4438 2617 4466 2618
rect 4438 2591 4439 2617
rect 4439 2591 4465 2617
rect 4465 2591 4466 2617
rect 4438 2590 4466 2591
rect 4158 2030 4186 2058
rect 4382 1134 4410 1162
rect 4718 182 4746 210
rect 5278 2646 5306 2674
rect 4998 2534 5026 2562
rect 4998 1190 5026 1218
rect 5054 742 5082 770
rect 5838 5782 5866 5810
rect 6510 6118 6538 6146
rect 6118 3878 6146 3906
rect 5446 2254 5474 2282
rect 5726 1974 5754 2002
rect 5502 406 5530 434
rect 6454 3345 6482 3346
rect 6454 3319 6455 3345
rect 6455 3319 6481 3345
rect 6481 3319 6482 3345
rect 6454 3318 6482 3319
rect 6454 2926 6482 2954
rect 6006 2478 6034 2506
rect 5950 2198 5978 2226
rect 5838 798 5866 826
rect 6454 2254 6482 2282
rect 6678 4998 6706 5026
rect 6510 1638 6538 1666
rect 6622 3934 6650 3962
rect 6286 742 6314 770
rect 6398 910 6426 938
rect 6174 686 6202 714
rect 7014 6566 7042 6594
rect 6902 6510 6930 6538
rect 6846 6398 6874 6426
rect 6790 6286 6818 6314
rect 6790 5838 6818 5866
rect 6734 4774 6762 4802
rect 7294 6566 7322 6594
rect 7238 6537 7266 6538
rect 7238 6511 7239 6537
rect 7239 6511 7265 6537
rect 7265 6511 7266 6537
rect 7238 6510 7266 6511
rect 8750 7014 8778 7042
rect 9142 7014 9170 7042
rect 7742 6678 7770 6706
rect 7350 6510 7378 6538
rect 7238 5558 7266 5586
rect 7238 4942 7266 4970
rect 7462 6454 7490 6482
rect 7462 4998 7490 5026
rect 7686 5110 7714 5138
rect 7686 4942 7714 4970
rect 7406 4774 7434 4802
rect 7014 4270 7042 4298
rect 7126 4438 7154 4466
rect 6846 3766 6874 3794
rect 6678 3430 6706 3458
rect 6734 3654 6762 3682
rect 6678 3262 6706 3290
rect 6734 3038 6762 3066
rect 6734 2870 6762 2898
rect 6734 2142 6762 2170
rect 6790 1246 6818 1274
rect 6678 1022 6706 1050
rect 7070 2758 7098 2786
rect 6846 798 6874 826
rect 6958 1414 6986 1442
rect 6790 630 6818 658
rect 6678 518 6706 546
rect 6846 462 6874 490
rect 6958 350 6986 378
rect 7238 3822 7266 3850
rect 7350 4326 7378 4354
rect 7126 2702 7154 2730
rect 7238 3206 7266 3234
rect 7126 1694 7154 1722
rect 7126 1358 7154 1386
rect 7182 1582 7210 1610
rect 7070 1302 7098 1330
rect 7014 238 7042 266
rect 7070 798 7098 826
rect 7350 2702 7378 2730
rect 7462 4606 7490 4634
rect 7462 4438 7490 4466
rect 7462 4326 7490 4354
rect 7462 4214 7490 4242
rect 7518 4102 7546 4130
rect 7574 4438 7602 4466
rect 7518 3822 7546 3850
rect 7518 3710 7546 3738
rect 7462 3598 7490 3626
rect 7406 2646 7434 2674
rect 7686 3374 7714 3402
rect 7518 2590 7546 2618
rect 7406 2366 7434 2394
rect 7238 1358 7266 1386
rect 7350 1246 7378 1274
rect 7350 686 7378 714
rect 7294 518 7322 546
rect 7406 406 7434 434
rect 7462 1190 7490 1218
rect 7182 294 7210 322
rect 7294 350 7322 378
rect 7462 294 7490 322
rect 7518 854 7546 882
rect 10206 7014 10234 7042
rect 10598 7014 10626 7042
rect 10262 6622 10290 6650
rect 9926 6454 9954 6482
rect 8750 6174 8778 6202
rect 8358 6062 8386 6090
rect 8246 5726 8274 5754
rect 8022 4494 8050 4522
rect 7910 1750 7938 1778
rect 8246 3318 8274 3346
rect 8302 4830 8330 4858
rect 8078 3038 8106 3066
rect 9086 5334 9114 5362
rect 10038 5166 10066 5194
rect 9086 4886 9114 4914
rect 9982 5054 10010 5082
rect 8358 4718 8386 4746
rect 8862 4718 8890 4746
rect 8358 4606 8386 4634
rect 8862 4214 8890 4242
rect 10206 5054 10234 5082
rect 10038 4214 10066 4242
rect 9982 3934 10010 3962
rect 8358 3654 8386 3682
rect 9758 3542 9786 3570
rect 9198 3486 9226 3514
rect 8862 3206 8890 3234
rect 8470 2198 8498 2226
rect 8302 1078 8330 1106
rect 8414 1918 8442 1946
rect 8078 966 8106 994
rect 8190 966 8218 994
rect 8022 798 8050 826
rect 7966 686 7994 714
rect 8414 798 8442 826
rect 8638 126 8666 154
rect 9086 2590 9114 2618
rect 8974 2057 9002 2058
rect 8974 2031 8975 2057
rect 8975 2031 9001 2057
rect 9001 2031 9002 2057
rect 8974 2030 9002 2031
rect 9086 1414 9114 1442
rect 9142 1918 9170 1946
rect 9870 3430 9898 3458
rect 9870 2814 9898 2842
rect 9926 2926 9954 2954
rect 9758 2702 9786 2730
rect 9198 1302 9226 1330
rect 9142 966 9170 994
rect 9310 630 9338 658
rect 9086 406 9114 434
rect 9422 630 9450 658
rect 9534 294 9562 322
rect 9982 2254 10010 2282
rect 9982 1190 10010 1218
rect 10990 6902 11018 6930
rect 10318 6481 10346 6482
rect 10318 6455 10319 6481
rect 10319 6455 10345 6481
rect 10345 6455 10346 6481
rect 10318 6454 10346 6455
rect 10598 6342 10626 6370
rect 10598 5558 10626 5586
rect 10934 5670 10962 5698
rect 10934 5446 10962 5474
rect 10318 4550 10346 4578
rect 10430 4550 10458 4578
rect 10654 4494 10682 4522
rect 10430 4438 10458 4466
rect 10542 4438 10570 4466
rect 10654 4326 10682 4354
rect 10934 4494 10962 4522
rect 10598 4270 10626 4298
rect 10822 4158 10850 4186
rect 10598 4046 10626 4074
rect 10542 3990 10570 4018
rect 10430 3598 10458 3626
rect 10262 3318 10290 3346
rect 10374 2926 10402 2954
rect 10318 2617 10346 2618
rect 10318 2591 10319 2617
rect 10319 2591 10345 2617
rect 10345 2591 10346 2617
rect 10318 2590 10346 2591
rect 10486 2758 10514 2786
rect 10374 2198 10402 2226
rect 10430 2254 10458 2282
rect 10038 966 10066 994
rect 10094 686 10122 714
rect 10206 686 10234 714
rect 10094 294 10122 322
rect 10206 574 10234 602
rect 10374 462 10402 490
rect 10486 2198 10514 2226
rect 10598 3878 10626 3906
rect 10598 3710 10626 3738
rect 10654 3822 10682 3850
rect 10598 2814 10626 2842
rect 12614 6790 12642 6818
rect 11662 6510 11690 6538
rect 12054 6678 12082 6706
rect 11046 6454 11074 6482
rect 11942 6481 11970 6482
rect 11942 6455 11943 6481
rect 11943 6455 11969 6481
rect 11969 6455 11970 6481
rect 11942 6454 11970 6455
rect 12232 6677 12260 6678
rect 12232 6651 12233 6677
rect 12233 6651 12259 6677
rect 12259 6651 12260 6677
rect 12232 6650 12260 6651
rect 12284 6677 12312 6678
rect 12284 6651 12285 6677
rect 12285 6651 12311 6677
rect 12311 6651 12312 6677
rect 12284 6650 12312 6651
rect 12336 6677 12364 6678
rect 12336 6651 12337 6677
rect 12337 6651 12363 6677
rect 12363 6651 12364 6677
rect 12336 6650 12364 6651
rect 12222 6510 12250 6538
rect 12054 6454 12082 6482
rect 11718 6286 11746 6314
rect 11158 5334 11186 5362
rect 11102 5110 11130 5138
rect 11902 6285 11930 6286
rect 11902 6259 11903 6285
rect 11903 6259 11929 6285
rect 11929 6259 11930 6285
rect 11902 6258 11930 6259
rect 11954 6285 11982 6286
rect 11954 6259 11955 6285
rect 11955 6259 11981 6285
rect 11981 6259 11982 6285
rect 11954 6258 11982 6259
rect 12006 6285 12034 6286
rect 12006 6259 12007 6285
rect 12007 6259 12033 6285
rect 12033 6259 12034 6285
rect 12006 6258 12034 6259
rect 12110 6286 12138 6314
rect 11774 6006 11802 6034
rect 11774 5838 11802 5866
rect 11718 5558 11746 5586
rect 11902 5501 11930 5502
rect 11902 5475 11903 5501
rect 11903 5475 11929 5501
rect 11929 5475 11930 5501
rect 11902 5474 11930 5475
rect 11954 5501 11982 5502
rect 11954 5475 11955 5501
rect 11955 5475 11981 5501
rect 11981 5475 11982 5501
rect 11954 5474 11982 5475
rect 12006 5501 12034 5502
rect 12006 5475 12007 5501
rect 12007 5475 12033 5501
rect 12033 5475 12034 5501
rect 12006 5474 12034 5475
rect 11326 5334 11354 5362
rect 11158 4998 11186 5026
rect 12232 5893 12260 5894
rect 12232 5867 12233 5893
rect 12233 5867 12259 5893
rect 12259 5867 12260 5893
rect 12232 5866 12260 5867
rect 12284 5893 12312 5894
rect 12284 5867 12285 5893
rect 12285 5867 12311 5893
rect 12311 5867 12312 5893
rect 12284 5866 12312 5867
rect 12336 5893 12364 5894
rect 12336 5867 12337 5893
rect 12337 5867 12363 5893
rect 12363 5867 12364 5893
rect 12336 5866 12364 5867
rect 12166 5726 12194 5754
rect 12278 5753 12306 5754
rect 12278 5727 12279 5753
rect 12279 5727 12305 5753
rect 12305 5727 12306 5753
rect 12278 5726 12306 5727
rect 12166 5446 12194 5474
rect 12446 5670 12474 5698
rect 12222 5222 12250 5250
rect 12166 5110 12194 5138
rect 12558 5697 12586 5698
rect 12558 5671 12559 5697
rect 12559 5671 12585 5697
rect 12585 5671 12586 5697
rect 12558 5670 12586 5671
rect 14574 7014 14602 7042
rect 14798 7014 14826 7042
rect 13566 6958 13594 6986
rect 12726 6230 12754 6258
rect 12726 5894 12754 5922
rect 13454 5950 13482 5978
rect 12950 5726 12978 5754
rect 13342 5838 13370 5866
rect 12782 5614 12810 5642
rect 12614 5390 12642 5418
rect 12232 5109 12260 5110
rect 12232 5083 12233 5109
rect 12233 5083 12259 5109
rect 12259 5083 12260 5109
rect 12232 5082 12260 5083
rect 12284 5109 12312 5110
rect 12284 5083 12285 5109
rect 12285 5083 12311 5109
rect 12311 5083 12312 5109
rect 12284 5082 12312 5083
rect 12336 5109 12364 5110
rect 12336 5083 12337 5109
rect 12337 5083 12363 5109
rect 12363 5083 12364 5109
rect 12446 5110 12474 5138
rect 12336 5082 12364 5083
rect 12558 4998 12586 5026
rect 12334 4942 12362 4970
rect 12110 4774 12138 4802
rect 12278 4774 12306 4802
rect 11102 4718 11130 4746
rect 11902 4717 11930 4718
rect 11902 4691 11903 4717
rect 11903 4691 11929 4717
rect 11929 4691 11930 4717
rect 11902 4690 11930 4691
rect 11954 4717 11982 4718
rect 11954 4691 11955 4717
rect 11955 4691 11981 4717
rect 11981 4691 11982 4717
rect 11954 4690 11982 4691
rect 12006 4717 12034 4718
rect 12006 4691 12007 4717
rect 12007 4691 12033 4717
rect 12033 4691 12034 4717
rect 12006 4690 12034 4691
rect 11662 4606 11690 4634
rect 12334 4606 12362 4634
rect 12278 4550 12306 4578
rect 12278 4438 12306 4466
rect 12446 4438 12474 4466
rect 12166 4326 12194 4354
rect 12232 4325 12260 4326
rect 11942 3990 11970 4018
rect 12110 4270 12138 4298
rect 12232 4299 12233 4325
rect 12233 4299 12259 4325
rect 12259 4299 12260 4325
rect 12232 4298 12260 4299
rect 12284 4325 12312 4326
rect 12284 4299 12285 4325
rect 12285 4299 12311 4325
rect 12311 4299 12312 4325
rect 12284 4298 12312 4299
rect 12336 4325 12364 4326
rect 12336 4299 12337 4325
rect 12337 4299 12363 4325
rect 12363 4299 12364 4325
rect 12336 4298 12364 4299
rect 11902 3933 11930 3934
rect 11902 3907 11903 3933
rect 11903 3907 11929 3933
rect 11929 3907 11930 3933
rect 11902 3906 11930 3907
rect 11954 3933 11982 3934
rect 11954 3907 11955 3933
rect 11955 3907 11981 3933
rect 11981 3907 11982 3933
rect 11954 3906 11982 3907
rect 12006 3933 12034 3934
rect 12006 3907 12007 3933
rect 12007 3907 12033 3933
rect 12033 3907 12034 3933
rect 12006 3906 12034 3907
rect 10990 3542 11018 3570
rect 11830 3486 11858 3514
rect 10710 3374 10738 3402
rect 11774 3374 11802 3402
rect 11550 3262 11578 3290
rect 11326 3150 11354 3178
rect 10934 2870 10962 2898
rect 10934 2646 10962 2674
rect 11158 2590 11186 2618
rect 10654 2310 10682 2338
rect 10542 1134 10570 1162
rect 10430 406 10458 434
rect 10430 126 10458 154
rect 10934 2142 10962 2170
rect 10766 1638 10794 1666
rect 10766 1414 10794 1442
rect 10822 1049 10850 1050
rect 10822 1023 10823 1049
rect 10823 1023 10849 1049
rect 10849 1023 10850 1049
rect 10822 1022 10850 1023
rect 10822 350 10850 378
rect 10878 742 10906 770
rect 10710 126 10738 154
rect 11046 630 11074 658
rect 11102 1750 11130 1778
rect 11494 2113 11522 2114
rect 11494 2087 11495 2113
rect 11495 2087 11521 2113
rect 11521 2087 11522 2113
rect 11494 2086 11522 2087
rect 11158 1078 11186 1106
rect 11214 1750 11242 1778
rect 11214 910 11242 938
rect 11326 574 11354 602
rect 11606 1078 11634 1106
rect 11662 574 11690 602
rect 12502 4158 12530 4186
rect 12614 4214 12642 4242
rect 12446 3766 12474 3794
rect 12232 3541 12260 3542
rect 12232 3515 12233 3541
rect 12233 3515 12259 3541
rect 12259 3515 12260 3541
rect 12232 3514 12260 3515
rect 12284 3541 12312 3542
rect 12284 3515 12285 3541
rect 12285 3515 12311 3541
rect 12311 3515 12312 3541
rect 12284 3514 12312 3515
rect 12336 3541 12364 3542
rect 12336 3515 12337 3541
rect 12337 3515 12363 3541
rect 12363 3515 12364 3541
rect 12336 3514 12364 3515
rect 12110 3262 12138 3290
rect 12782 4969 12810 4970
rect 12782 4943 12783 4969
rect 12783 4943 12809 4969
rect 12809 4943 12810 4969
rect 12782 4942 12810 4943
rect 13062 4886 13090 4914
rect 12838 4662 12866 4690
rect 12726 4270 12754 4298
rect 12726 3822 12754 3850
rect 12782 4102 12810 4130
rect 12670 3430 12698 3458
rect 12726 3542 12754 3570
rect 11902 3149 11930 3150
rect 11902 3123 11903 3149
rect 11903 3123 11929 3149
rect 11929 3123 11930 3149
rect 11902 3122 11930 3123
rect 11954 3149 11982 3150
rect 11954 3123 11955 3149
rect 11955 3123 11981 3149
rect 11981 3123 11982 3149
rect 11954 3122 11982 3123
rect 12006 3149 12034 3150
rect 12006 3123 12007 3149
rect 12007 3123 12033 3149
rect 12033 3123 12034 3149
rect 12614 3150 12642 3178
rect 12670 3206 12698 3234
rect 12006 3122 12034 3123
rect 12614 3038 12642 3066
rect 12232 2757 12260 2758
rect 11830 2646 11858 2674
rect 12166 2702 12194 2730
rect 12232 2731 12233 2757
rect 12233 2731 12259 2757
rect 12259 2731 12260 2757
rect 12232 2730 12260 2731
rect 12284 2757 12312 2758
rect 12284 2731 12285 2757
rect 12285 2731 12311 2757
rect 12311 2731 12312 2757
rect 12284 2730 12312 2731
rect 12336 2757 12364 2758
rect 12336 2731 12337 2757
rect 12337 2731 12363 2757
rect 12363 2731 12364 2757
rect 12336 2730 12364 2731
rect 12446 2702 12474 2730
rect 11902 2365 11930 2366
rect 11902 2339 11903 2365
rect 11903 2339 11929 2365
rect 11929 2339 11930 2365
rect 11902 2338 11930 2339
rect 11954 2365 11982 2366
rect 11954 2339 11955 2365
rect 11955 2339 11981 2365
rect 11981 2339 11982 2365
rect 11954 2338 11982 2339
rect 12006 2365 12034 2366
rect 12006 2339 12007 2365
rect 12007 2339 12033 2365
rect 12033 2339 12034 2365
rect 12614 2366 12642 2394
rect 12006 2338 12034 2339
rect 12232 1973 12260 1974
rect 12232 1947 12233 1973
rect 12233 1947 12259 1973
rect 12259 1947 12260 1973
rect 12232 1946 12260 1947
rect 12284 1973 12312 1974
rect 12284 1947 12285 1973
rect 12285 1947 12311 1973
rect 12311 1947 12312 1973
rect 12284 1946 12312 1947
rect 12336 1973 12364 1974
rect 12336 1947 12337 1973
rect 12337 1947 12363 1973
rect 12363 1947 12364 1973
rect 12336 1946 12364 1947
rect 12614 1806 12642 1834
rect 11902 1581 11930 1582
rect 11902 1555 11903 1581
rect 11903 1555 11929 1581
rect 11929 1555 11930 1581
rect 11902 1554 11930 1555
rect 11954 1581 11982 1582
rect 11954 1555 11955 1581
rect 11955 1555 11981 1581
rect 11981 1555 11982 1581
rect 11954 1554 11982 1555
rect 12006 1581 12034 1582
rect 12006 1555 12007 1581
rect 12007 1555 12033 1581
rect 12033 1555 12034 1581
rect 12006 1554 12034 1555
rect 12166 1526 12194 1554
rect 13454 5782 13482 5810
rect 13454 5502 13482 5530
rect 13342 4326 13370 4354
rect 13398 5166 13426 5194
rect 13006 4214 13034 4242
rect 12838 3374 12866 3402
rect 12894 3990 12922 4018
rect 12894 2926 12922 2954
rect 12726 2254 12754 2282
rect 12782 2758 12810 2786
rect 12558 1526 12586 1554
rect 12166 1190 12194 1218
rect 12232 1189 12260 1190
rect 12232 1163 12233 1189
rect 12233 1163 12259 1189
rect 12259 1163 12260 1189
rect 12232 1162 12260 1163
rect 12284 1189 12312 1190
rect 12284 1163 12285 1189
rect 12285 1163 12311 1189
rect 12311 1163 12312 1189
rect 12284 1162 12312 1163
rect 12336 1189 12364 1190
rect 12336 1163 12337 1189
rect 12337 1163 12363 1189
rect 12363 1163 12364 1189
rect 12336 1162 12364 1163
rect 12390 937 12418 938
rect 12390 911 12391 937
rect 12391 911 12417 937
rect 12417 911 12418 937
rect 12390 910 12418 911
rect 11902 797 11930 798
rect 11902 771 11903 797
rect 11903 771 11929 797
rect 11929 771 11930 797
rect 11902 770 11930 771
rect 11954 797 11982 798
rect 11954 771 11955 797
rect 11955 771 11981 797
rect 11981 771 11982 797
rect 11954 770 11982 771
rect 12006 797 12034 798
rect 12006 771 12007 797
rect 12007 771 12033 797
rect 12033 771 12034 797
rect 12006 770 12034 771
rect 11998 630 12026 658
rect 12446 462 12474 490
rect 12232 405 12260 406
rect 12232 379 12233 405
rect 12233 379 12259 405
rect 12259 379 12260 405
rect 12232 378 12260 379
rect 12284 405 12312 406
rect 12284 379 12285 405
rect 12285 379 12311 405
rect 12311 379 12312 405
rect 12284 378 12312 379
rect 12336 405 12364 406
rect 12336 379 12337 405
rect 12337 379 12363 405
rect 12363 379 12364 405
rect 12336 378 12364 379
rect 12222 238 12250 266
rect 12894 1750 12922 1778
rect 16030 7014 16058 7042
rect 16254 7014 16282 7042
rect 15750 6790 15778 6818
rect 14294 6342 14322 6370
rect 13566 5502 13594 5530
rect 13790 6230 13818 6258
rect 13454 4998 13482 5026
rect 13398 4158 13426 4186
rect 13678 4102 13706 4130
rect 13398 3934 13426 3962
rect 13062 3793 13090 3794
rect 13062 3767 13063 3793
rect 13063 3767 13089 3793
rect 13089 3767 13090 3793
rect 13062 3766 13090 3767
rect 13342 3430 13370 3458
rect 13342 3318 13370 3346
rect 13118 3262 13146 3290
rect 14238 6006 14266 6034
rect 14238 5614 14266 5642
rect 14126 5446 14154 5474
rect 14014 4774 14042 4802
rect 13790 3654 13818 3682
rect 13846 3990 13874 4018
rect 13734 2590 13762 2618
rect 13454 2534 13482 2562
rect 13454 2030 13482 2058
rect 13510 2198 13538 2226
rect 13006 1414 13034 1442
rect 13174 1582 13202 1610
rect 12838 1358 12866 1386
rect 12782 854 12810 882
rect 13118 574 13146 602
rect 12894 518 12922 546
rect 13286 1470 13314 1498
rect 13678 1862 13706 1890
rect 13958 3681 13986 3682
rect 13958 3655 13959 3681
rect 13959 3655 13985 3681
rect 13985 3655 13986 3681
rect 13958 3654 13986 3655
rect 14014 3094 14042 3122
rect 14070 4494 14098 4522
rect 14238 5222 14266 5250
rect 14182 4606 14210 4634
rect 14798 5894 14826 5922
rect 14686 5278 14714 5306
rect 14518 4577 14546 4578
rect 14518 4551 14519 4577
rect 14519 4551 14545 4577
rect 14545 4551 14546 4577
rect 14518 4550 14546 4551
rect 14182 4102 14210 4130
rect 14126 3878 14154 3906
rect 14070 2590 14098 2618
rect 14126 3710 14154 3738
rect 14014 2254 14042 2282
rect 13846 1582 13874 1610
rect 13510 1470 13538 1498
rect 14294 3486 14322 3514
rect 14182 3038 14210 3066
rect 14966 5782 14994 5810
rect 15302 5726 15330 5754
rect 15694 5390 15722 5418
rect 14966 5222 14994 5250
rect 14854 5166 14882 5194
rect 14910 4214 14938 4242
rect 15638 5193 15666 5194
rect 15638 5167 15639 5193
rect 15639 5167 15665 5193
rect 15665 5167 15666 5193
rect 15638 5166 15666 5167
rect 15190 5110 15218 5138
rect 15134 4494 15162 4522
rect 15134 4046 15162 4074
rect 14966 3766 14994 3794
rect 15078 3822 15106 3850
rect 15022 3737 15050 3738
rect 15022 3711 15023 3737
rect 15023 3711 15049 3737
rect 15049 3711 15050 3737
rect 15022 3710 15050 3711
rect 14910 3374 14938 3402
rect 14854 3206 14882 3234
rect 14798 3038 14826 3066
rect 15582 3374 15610 3402
rect 15358 3345 15386 3346
rect 15358 3319 15359 3345
rect 15359 3319 15385 3345
rect 15385 3319 15386 3345
rect 15358 3318 15386 3319
rect 15190 3206 15218 3234
rect 14294 1918 14322 1946
rect 14350 2814 14378 2842
rect 14182 1582 14210 1610
rect 14294 1806 14322 1834
rect 14294 1414 14322 1442
rect 13902 1358 13930 1386
rect 14742 2366 14770 2394
rect 14686 1862 14714 1890
rect 13678 1273 13706 1274
rect 13678 1247 13679 1273
rect 13679 1247 13705 1273
rect 13705 1247 13706 1273
rect 13678 1246 13706 1247
rect 13846 1246 13874 1274
rect 13454 1134 13482 1162
rect 13342 545 13370 546
rect 13342 519 13343 545
rect 13343 519 13369 545
rect 13369 519 13370 545
rect 13342 518 13370 519
rect 12894 406 12922 434
rect 13734 993 13762 994
rect 13734 967 13735 993
rect 13735 967 13761 993
rect 13761 967 13762 993
rect 13734 966 13762 967
rect 13566 630 13594 658
rect 13790 518 13818 546
rect 13454 182 13482 210
rect 13566 350 13594 378
rect 13342 126 13370 154
rect 13958 1190 13986 1218
rect 14070 1078 14098 1106
rect 13846 294 13874 322
rect 14014 462 14042 490
rect 14406 462 14434 490
rect 14686 1134 14714 1162
rect 14518 1049 14546 1050
rect 14518 1023 14519 1049
rect 14519 1023 14545 1049
rect 14545 1023 14546 1049
rect 14518 1022 14546 1023
rect 14742 686 14770 714
rect 14854 601 14882 602
rect 14854 575 14855 601
rect 14855 575 14881 601
rect 14881 575 14882 601
rect 14854 574 14882 575
rect 15078 2870 15106 2898
rect 15526 1750 15554 1778
rect 15190 1694 15218 1722
rect 15078 1526 15106 1554
rect 15134 1329 15162 1330
rect 15134 1303 15135 1329
rect 15135 1303 15161 1329
rect 15161 1303 15162 1329
rect 15134 1302 15162 1303
rect 15470 1022 15498 1050
rect 15638 1582 15666 1610
rect 15022 406 15050 434
rect 17486 7014 17514 7042
rect 17766 7014 17794 7042
rect 16702 6790 16730 6818
rect 16534 6286 16562 6314
rect 16198 5753 16226 5754
rect 16198 5727 16199 5753
rect 16199 5727 16225 5753
rect 16225 5727 16226 5753
rect 16198 5726 16226 5727
rect 16422 5614 16450 5642
rect 15806 5502 15834 5530
rect 15918 5110 15946 5138
rect 16310 5054 16338 5082
rect 15974 4830 16002 4858
rect 16310 4774 16338 4802
rect 16030 4438 16058 4466
rect 16646 6230 16674 6258
rect 16030 3262 16058 3290
rect 15974 2646 16002 2674
rect 16142 2814 16170 2842
rect 15974 2113 16002 2114
rect 15974 2087 15975 2113
rect 15975 2087 16001 2113
rect 16001 2087 16002 2113
rect 15974 2086 16002 2087
rect 15918 1833 15946 1834
rect 15918 1807 15919 1833
rect 15919 1807 15945 1833
rect 15945 1807 15946 1833
rect 15918 1806 15946 1807
rect 15806 1638 15834 1666
rect 15750 1582 15778 1610
rect 15974 1385 16002 1386
rect 15974 1359 15975 1385
rect 15975 1359 16001 1385
rect 16001 1359 16002 1385
rect 15974 1358 16002 1359
rect 15862 1246 15890 1274
rect 15806 630 15834 658
rect 15638 462 15666 490
rect 16422 2534 16450 2562
rect 16254 2113 16282 2114
rect 16254 2087 16255 2113
rect 16255 2087 16281 2113
rect 16281 2087 16282 2113
rect 16254 2086 16282 2087
rect 16198 1889 16226 1890
rect 16198 1863 16199 1889
rect 16199 1863 16225 1889
rect 16225 1863 16226 1889
rect 16198 1862 16226 1863
rect 16478 2422 16506 2450
rect 16534 2198 16562 2226
rect 16590 2422 16618 2450
rect 17318 6734 17346 6762
rect 16758 6481 16786 6482
rect 16758 6455 16759 6481
rect 16759 6455 16785 6481
rect 16785 6455 16786 6481
rect 16758 6454 16786 6455
rect 16814 6342 16842 6370
rect 16758 6033 16786 6034
rect 16758 6007 16759 6033
rect 16759 6007 16785 6033
rect 16785 6007 16786 6033
rect 16758 6006 16786 6007
rect 17486 6454 17514 6482
rect 16702 5726 16730 5754
rect 17206 6006 17234 6034
rect 16758 5278 16786 5306
rect 16758 4942 16786 4970
rect 16870 5054 16898 5082
rect 16758 4326 16786 4354
rect 16926 4494 16954 4522
rect 16982 4409 17010 4410
rect 16982 4383 16983 4409
rect 16983 4383 17009 4409
rect 17009 4383 17010 4409
rect 16982 4382 17010 4383
rect 16926 4326 16954 4354
rect 16814 4102 16842 4130
rect 16870 4270 16898 4298
rect 16814 3542 16842 3570
rect 16758 3430 16786 3458
rect 16646 2366 16674 2394
rect 16702 3374 16730 3402
rect 16758 2982 16786 3010
rect 16982 2673 17010 2674
rect 16982 2647 16983 2673
rect 16983 2647 17009 2673
rect 17009 2647 17010 2673
rect 16982 2646 17010 2647
rect 17262 4521 17290 4522
rect 17262 4495 17263 4521
rect 17263 4495 17289 4521
rect 17289 4495 17290 4521
rect 17262 4494 17290 4495
rect 18438 6510 18466 6538
rect 20398 7014 20426 7042
rect 20622 7014 20650 7042
rect 18270 6481 18298 6482
rect 18270 6455 18271 6481
rect 18271 6455 18297 6481
rect 18297 6455 18298 6481
rect 18270 6454 18298 6455
rect 17598 5894 17626 5922
rect 18382 5670 18410 5698
rect 19222 6454 19250 6482
rect 18606 6118 18634 6146
rect 18886 6033 18914 6034
rect 18886 6007 18887 6033
rect 18887 6007 18913 6033
rect 18913 6007 18914 6033
rect 18886 6006 18914 6007
rect 18774 5950 18802 5978
rect 18438 5446 18466 5474
rect 18494 5838 18522 5866
rect 18718 5558 18746 5586
rect 18382 4942 18410 4970
rect 18718 4998 18746 5026
rect 18270 4718 18298 4746
rect 17542 4326 17570 4354
rect 17766 3878 17794 3906
rect 17766 3486 17794 3514
rect 17206 2646 17234 2674
rect 16758 2478 16786 2506
rect 16702 2142 16730 2170
rect 16422 1582 16450 1610
rect 16198 1273 16226 1274
rect 16198 1247 16199 1273
rect 16199 1247 16225 1273
rect 16225 1247 16226 1273
rect 16198 1246 16226 1247
rect 16366 1049 16394 1050
rect 16366 1023 16367 1049
rect 16367 1023 16393 1049
rect 16393 1023 16394 1049
rect 16366 1022 16394 1023
rect 16814 1414 16842 1442
rect 16758 1022 16786 1050
rect 16142 350 16170 378
rect 16198 854 16226 882
rect 16198 238 16226 266
rect 16758 854 16786 882
rect 17150 1190 17178 1218
rect 17150 630 17178 658
rect 16926 462 16954 490
rect 17262 2086 17290 2114
rect 18158 3374 18186 3402
rect 18158 3150 18186 3178
rect 18214 2702 18242 2730
rect 18214 1721 18242 1722
rect 18214 1695 18215 1721
rect 18215 1695 18241 1721
rect 18241 1695 18242 1721
rect 18214 1694 18242 1695
rect 18494 4438 18522 4466
rect 18438 4326 18466 4354
rect 18438 4046 18466 4074
rect 18382 3542 18410 3570
rect 18382 3150 18410 3178
rect 18438 3206 18466 3234
rect 18270 1358 18298 1386
rect 18326 2198 18354 2226
rect 17598 1078 17626 1106
rect 17206 574 17234 602
rect 17374 966 17402 994
rect 17430 881 17458 882
rect 17430 855 17431 881
rect 17431 855 17457 881
rect 17457 855 17458 881
rect 17430 854 17458 855
rect 17598 686 17626 714
rect 17934 1049 17962 1050
rect 17934 1023 17935 1049
rect 17935 1023 17961 1049
rect 17961 1023 17962 1049
rect 17934 1022 17962 1023
rect 18214 966 18242 994
rect 18046 854 18074 882
rect 17654 630 17682 658
rect 17822 630 17850 658
rect 17654 545 17682 546
rect 17654 519 17655 545
rect 17655 519 17681 545
rect 17681 519 17682 545
rect 17654 518 17682 519
rect 17598 406 17626 434
rect 17934 489 17962 490
rect 17934 463 17935 489
rect 17935 463 17961 489
rect 17961 463 17962 489
rect 17934 462 17962 463
rect 18270 798 18298 826
rect 18438 2142 18466 2170
rect 18494 2702 18522 2730
rect 18382 1918 18410 1946
rect 18438 1862 18466 1890
rect 18438 1526 18466 1554
rect 18494 1414 18522 1442
rect 18382 686 18410 714
rect 19054 5894 19082 5922
rect 18886 4270 18914 4298
rect 18830 2169 18858 2170
rect 18830 2143 18831 2169
rect 18831 2143 18857 2169
rect 18857 2143 18858 2169
rect 18830 2142 18858 2143
rect 18774 1582 18802 1610
rect 18942 1385 18970 1386
rect 18942 1359 18943 1385
rect 18943 1359 18969 1385
rect 18969 1359 18970 1385
rect 18942 1358 18970 1359
rect 18774 1246 18802 1274
rect 18662 798 18690 826
rect 18550 630 18578 658
rect 18438 601 18466 602
rect 18438 575 18439 601
rect 18439 575 18465 601
rect 18465 575 18466 601
rect 18438 574 18466 575
rect 18382 294 18410 322
rect 18494 518 18522 546
rect 18326 126 18354 154
rect 18718 489 18746 490
rect 18718 463 18719 489
rect 18719 463 18745 489
rect 18745 463 18746 489
rect 18718 462 18746 463
rect 19166 4382 19194 4410
rect 19166 2617 19194 2618
rect 19166 2591 19167 2617
rect 19167 2591 19193 2617
rect 19193 2591 19194 2617
rect 19166 2590 19194 2591
rect 19110 2113 19138 2114
rect 19110 2087 19111 2113
rect 19111 2087 19137 2113
rect 19137 2087 19138 2113
rect 19110 2086 19138 2087
rect 19166 1777 19194 1778
rect 19166 1751 19167 1777
rect 19167 1751 19193 1777
rect 19193 1751 19194 1777
rect 19166 1750 19194 1751
rect 21854 7014 21882 7042
rect 22078 7014 22106 7042
rect 20846 6089 20874 6090
rect 20846 6063 20847 6089
rect 20847 6063 20873 6089
rect 20873 6063 20874 6089
rect 20846 6062 20874 6063
rect 21126 6089 21154 6090
rect 21126 6063 21127 6089
rect 21127 6063 21153 6089
rect 21153 6063 21154 6089
rect 21126 6062 21154 6063
rect 19446 5054 19474 5082
rect 19558 4774 19586 4802
rect 19446 4438 19474 4466
rect 19222 1358 19250 1386
rect 19222 1273 19250 1274
rect 19222 1247 19223 1273
rect 19223 1247 19249 1273
rect 19249 1247 19250 1273
rect 19222 1246 19250 1247
rect 19054 1134 19082 1162
rect 18998 881 19026 882
rect 18998 855 18999 881
rect 18999 855 19025 881
rect 19025 855 19026 881
rect 18998 854 19026 855
rect 19166 854 19194 882
rect 18942 462 18970 490
rect 19446 406 19474 434
rect 20398 5977 20426 5978
rect 20398 5951 20399 5977
rect 20399 5951 20425 5977
rect 20425 5951 20426 5977
rect 20398 5950 20426 5951
rect 19726 5641 19754 5642
rect 19726 5615 19727 5641
rect 19727 5615 19753 5641
rect 19753 5615 19754 5641
rect 19726 5614 19754 5615
rect 20286 4774 20314 4802
rect 20118 4662 20146 4690
rect 19670 4214 19698 4242
rect 20566 4326 20594 4354
rect 20118 3318 20146 3346
rect 20342 3822 20370 3850
rect 20006 2702 20034 2730
rect 20678 3822 20706 3850
rect 20398 3150 20426 3178
rect 20958 5950 20986 5978
rect 20958 5726 20986 5754
rect 20958 4158 20986 4186
rect 20902 3766 20930 3794
rect 20790 3598 20818 3626
rect 20790 3262 20818 3290
rect 20846 2982 20874 3010
rect 21070 4158 21098 4186
rect 21070 3878 21098 3906
rect 20958 2478 20986 2506
rect 20902 2366 20930 2394
rect 20734 2310 20762 2338
rect 20342 2142 20370 2170
rect 20174 1974 20202 2002
rect 19726 1694 19754 1722
rect 19894 1694 19922 1722
rect 19614 1078 19642 1106
rect 19502 350 19530 378
rect 19390 294 19418 322
rect 19782 993 19810 994
rect 19782 967 19783 993
rect 19783 967 19809 993
rect 19809 967 19810 993
rect 19782 966 19810 967
rect 19838 518 19866 546
rect 20230 1721 20258 1722
rect 20230 1695 20231 1721
rect 20231 1695 20257 1721
rect 20257 1695 20258 1721
rect 20230 1694 20258 1695
rect 20342 1470 20370 1498
rect 20174 1246 20202 1274
rect 20118 993 20146 994
rect 20118 967 20119 993
rect 20119 967 20145 993
rect 20145 967 20146 993
rect 20118 966 20146 967
rect 20006 854 20034 882
rect 20062 630 20090 658
rect 20174 238 20202 266
rect 20230 966 20258 994
rect 20510 2086 20538 2114
rect 20734 2086 20762 2114
rect 21070 2113 21098 2114
rect 21070 2087 21071 2113
rect 21071 2087 21097 2113
rect 21097 2087 21098 2113
rect 21070 2086 21098 2087
rect 20790 2057 20818 2058
rect 20790 2031 20791 2057
rect 20791 2031 20817 2057
rect 20817 2031 20818 2057
rect 20790 2030 20818 2031
rect 20510 1470 20538 1498
rect 20230 182 20258 210
rect 20286 518 20314 546
rect 20398 294 20426 322
rect 20510 798 20538 826
rect 20622 489 20650 490
rect 20622 463 20623 489
rect 20623 463 20649 489
rect 20649 463 20650 489
rect 20622 462 20650 463
rect 23310 7014 23338 7042
rect 23534 7014 23562 7042
rect 22232 6677 22260 6678
rect 22232 6651 22233 6677
rect 22233 6651 22259 6677
rect 22259 6651 22260 6677
rect 22232 6650 22260 6651
rect 22284 6677 22312 6678
rect 22284 6651 22285 6677
rect 22285 6651 22311 6677
rect 22311 6651 22312 6677
rect 22284 6650 22312 6651
rect 22336 6677 22364 6678
rect 22336 6651 22337 6677
rect 22337 6651 22363 6677
rect 22363 6651 22364 6677
rect 22336 6650 22364 6651
rect 21902 6285 21930 6286
rect 21902 6259 21903 6285
rect 21903 6259 21929 6285
rect 21929 6259 21930 6285
rect 21902 6258 21930 6259
rect 21954 6285 21982 6286
rect 21954 6259 21955 6285
rect 21955 6259 21981 6285
rect 21981 6259 21982 6285
rect 21954 6258 21982 6259
rect 22006 6285 22034 6286
rect 22006 6259 22007 6285
rect 22007 6259 22033 6285
rect 22033 6259 22034 6285
rect 22006 6258 22034 6259
rect 22232 5893 22260 5894
rect 22232 5867 22233 5893
rect 22233 5867 22259 5893
rect 22259 5867 22260 5893
rect 22232 5866 22260 5867
rect 22284 5893 22312 5894
rect 22284 5867 22285 5893
rect 22285 5867 22311 5893
rect 22311 5867 22312 5893
rect 22284 5866 22312 5867
rect 22336 5893 22364 5894
rect 22336 5867 22337 5893
rect 22337 5867 22363 5893
rect 22363 5867 22364 5893
rect 22336 5866 22364 5867
rect 21742 5502 21770 5530
rect 21798 5670 21826 5698
rect 21518 5446 21546 5474
rect 21462 2534 21490 2562
rect 21902 5501 21930 5502
rect 21902 5475 21903 5501
rect 21903 5475 21929 5501
rect 21929 5475 21930 5501
rect 21902 5474 21930 5475
rect 21954 5501 21982 5502
rect 21954 5475 21955 5501
rect 21955 5475 21981 5501
rect 21981 5475 21982 5501
rect 21954 5474 21982 5475
rect 22006 5501 22034 5502
rect 22006 5475 22007 5501
rect 22007 5475 22033 5501
rect 22033 5475 22034 5501
rect 22006 5474 22034 5475
rect 21798 4942 21826 4970
rect 22232 5109 22260 5110
rect 22232 5083 22233 5109
rect 22233 5083 22259 5109
rect 22259 5083 22260 5109
rect 22232 5082 22260 5083
rect 22284 5109 22312 5110
rect 22284 5083 22285 5109
rect 22285 5083 22311 5109
rect 22311 5083 22312 5109
rect 22284 5082 22312 5083
rect 22336 5109 22364 5110
rect 22336 5083 22337 5109
rect 22337 5083 22363 5109
rect 22363 5083 22364 5109
rect 22336 5082 22364 5083
rect 22078 4830 22106 4858
rect 22414 4774 22442 4802
rect 21902 4717 21930 4718
rect 21902 4691 21903 4717
rect 21903 4691 21929 4717
rect 21929 4691 21930 4717
rect 21902 4690 21930 4691
rect 21954 4717 21982 4718
rect 21954 4691 21955 4717
rect 21955 4691 21981 4717
rect 21981 4691 21982 4717
rect 21954 4690 21982 4691
rect 22006 4717 22034 4718
rect 22006 4691 22007 4717
rect 22007 4691 22033 4717
rect 22033 4691 22034 4717
rect 22006 4690 22034 4691
rect 21966 4606 21994 4634
rect 22414 4606 22442 4634
rect 22190 4550 22218 4578
rect 22232 4325 22260 4326
rect 22232 4299 22233 4325
rect 22233 4299 22259 4325
rect 22259 4299 22260 4325
rect 22232 4298 22260 4299
rect 22284 4325 22312 4326
rect 22284 4299 22285 4325
rect 22285 4299 22311 4325
rect 22311 4299 22312 4325
rect 22284 4298 22312 4299
rect 22336 4325 22364 4326
rect 22336 4299 22337 4325
rect 22337 4299 22363 4325
rect 22363 4299 22364 4325
rect 22336 4298 22364 4299
rect 22414 4214 22442 4242
rect 21902 3933 21930 3934
rect 21902 3907 21903 3933
rect 21903 3907 21929 3933
rect 21929 3907 21930 3933
rect 21902 3906 21930 3907
rect 21954 3933 21982 3934
rect 21954 3907 21955 3933
rect 21955 3907 21981 3933
rect 21981 3907 21982 3933
rect 21954 3906 21982 3907
rect 22006 3933 22034 3934
rect 22006 3907 22007 3933
rect 22007 3907 22033 3933
rect 22033 3907 22034 3933
rect 22006 3906 22034 3907
rect 22232 3541 22260 3542
rect 22232 3515 22233 3541
rect 22233 3515 22259 3541
rect 22259 3515 22260 3541
rect 22232 3514 22260 3515
rect 22284 3541 22312 3542
rect 22284 3515 22285 3541
rect 22285 3515 22311 3541
rect 22311 3515 22312 3541
rect 22284 3514 22312 3515
rect 22336 3541 22364 3542
rect 22336 3515 22337 3541
rect 22337 3515 22363 3541
rect 22363 3515 22364 3541
rect 22336 3514 22364 3515
rect 21686 3374 21714 3402
rect 21630 2478 21658 2506
rect 21902 3149 21930 3150
rect 21902 3123 21903 3149
rect 21903 3123 21929 3149
rect 21929 3123 21930 3149
rect 21902 3122 21930 3123
rect 21954 3149 21982 3150
rect 21954 3123 21955 3149
rect 21955 3123 21981 3149
rect 21981 3123 21982 3149
rect 21954 3122 21982 3123
rect 22006 3149 22034 3150
rect 22006 3123 22007 3149
rect 22007 3123 22033 3149
rect 22033 3123 22034 3149
rect 22414 3150 22442 3178
rect 22526 3206 22554 3234
rect 22006 3122 22034 3123
rect 22582 3094 22610 3122
rect 22134 2758 22162 2786
rect 22232 2757 22260 2758
rect 22232 2731 22233 2757
rect 22233 2731 22259 2757
rect 22259 2731 22260 2757
rect 22232 2730 22260 2731
rect 22284 2757 22312 2758
rect 22284 2731 22285 2757
rect 22285 2731 22311 2757
rect 22311 2731 22312 2757
rect 22284 2730 22312 2731
rect 22336 2757 22364 2758
rect 22336 2731 22337 2757
rect 22337 2731 22363 2757
rect 22363 2731 22364 2757
rect 22336 2730 22364 2731
rect 21686 2030 21714 2058
rect 21238 1414 21266 1442
rect 21406 1694 21434 1722
rect 21294 1329 21322 1330
rect 21294 1303 21295 1329
rect 21295 1303 21321 1329
rect 21321 1303 21322 1329
rect 21294 1302 21322 1303
rect 21182 1105 21210 1106
rect 21182 1079 21183 1105
rect 21183 1079 21209 1105
rect 21209 1079 21210 1105
rect 21182 1078 21210 1079
rect 20902 1049 20930 1050
rect 20902 1023 20903 1049
rect 20903 1023 20929 1049
rect 20929 1023 20930 1049
rect 20902 1022 20930 1023
rect 20790 630 20818 658
rect 20958 630 20986 658
rect 21182 462 21210 490
rect 21630 1302 21658 1330
rect 22470 2561 22498 2562
rect 22470 2535 22471 2561
rect 22471 2535 22497 2561
rect 22497 2535 22498 2561
rect 22470 2534 22498 2535
rect 21902 2365 21930 2366
rect 21902 2339 21903 2365
rect 21903 2339 21929 2365
rect 21929 2339 21930 2365
rect 21902 2338 21930 2339
rect 21954 2365 21982 2366
rect 21954 2339 21955 2365
rect 21955 2339 21981 2365
rect 21981 2339 21982 2365
rect 21954 2338 21982 2339
rect 22006 2365 22034 2366
rect 22006 2339 22007 2365
rect 22007 2339 22033 2365
rect 22033 2339 22034 2365
rect 22006 2338 22034 2339
rect 21798 2198 21826 2226
rect 22232 1973 22260 1974
rect 22232 1947 22233 1973
rect 22233 1947 22259 1973
rect 22259 1947 22260 1973
rect 22232 1946 22260 1947
rect 22284 1973 22312 1974
rect 22284 1947 22285 1973
rect 22285 1947 22311 1973
rect 22311 1947 22312 1973
rect 22284 1946 22312 1947
rect 22336 1973 22364 1974
rect 22336 1947 22337 1973
rect 22337 1947 22363 1973
rect 22363 1947 22364 1973
rect 22336 1946 22364 1947
rect 22302 1777 22330 1778
rect 22302 1751 22303 1777
rect 22303 1751 22329 1777
rect 22329 1751 22330 1777
rect 22302 1750 22330 1751
rect 21798 1721 21826 1722
rect 21798 1695 21799 1721
rect 21799 1695 21825 1721
rect 21825 1695 21826 1721
rect 21798 1694 21826 1695
rect 21902 1581 21930 1582
rect 21902 1555 21903 1581
rect 21903 1555 21929 1581
rect 21929 1555 21930 1581
rect 21902 1554 21930 1555
rect 21954 1581 21982 1582
rect 21954 1555 21955 1581
rect 21955 1555 21981 1581
rect 21981 1555 21982 1581
rect 21954 1554 21982 1555
rect 22006 1581 22034 1582
rect 22006 1555 22007 1581
rect 22007 1555 22033 1581
rect 22033 1555 22034 1581
rect 22006 1554 22034 1555
rect 24094 6846 24122 6874
rect 24038 6118 24066 6146
rect 23534 5614 23562 5642
rect 23534 3542 23562 3570
rect 22694 3374 22722 3402
rect 22694 3262 22722 3290
rect 23422 3038 23450 3066
rect 22638 2366 22666 2394
rect 22694 2646 22722 2674
rect 22638 2198 22666 2226
rect 22302 1329 22330 1330
rect 22302 1303 22303 1329
rect 22303 1303 22329 1329
rect 22329 1303 22330 1329
rect 22302 1302 22330 1303
rect 22470 1302 22498 1330
rect 22232 1189 22260 1190
rect 22232 1163 22233 1189
rect 22233 1163 22259 1189
rect 22259 1163 22260 1189
rect 22232 1162 22260 1163
rect 22284 1189 22312 1190
rect 22284 1163 22285 1189
rect 22285 1163 22311 1189
rect 22311 1163 22312 1189
rect 22284 1162 22312 1163
rect 22336 1189 22364 1190
rect 22336 1163 22337 1189
rect 22337 1163 22363 1189
rect 22363 1163 22364 1189
rect 22336 1162 22364 1163
rect 22414 1022 22442 1050
rect 21966 881 21994 882
rect 21966 855 21967 881
rect 21967 855 21993 881
rect 21993 855 21994 881
rect 21966 854 21994 855
rect 21902 797 21930 798
rect 21902 771 21903 797
rect 21903 771 21929 797
rect 21929 771 21930 797
rect 21902 770 21930 771
rect 21954 797 21982 798
rect 21954 771 21955 797
rect 21955 771 21981 797
rect 21981 771 21982 797
rect 21954 770 21982 771
rect 22006 797 22034 798
rect 22006 771 22007 797
rect 22007 771 22033 797
rect 22033 771 22034 797
rect 22006 770 22034 771
rect 22078 742 22106 770
rect 21854 545 21882 546
rect 21854 519 21855 545
rect 21855 519 21881 545
rect 21881 519 21882 545
rect 21854 518 21882 519
rect 21854 182 21882 210
rect 22358 657 22386 658
rect 22358 631 22359 657
rect 22359 631 22385 657
rect 22385 631 22386 657
rect 22358 630 22386 631
rect 22232 405 22260 406
rect 22232 379 22233 405
rect 22233 379 22259 405
rect 22259 379 22260 405
rect 22232 378 22260 379
rect 22284 405 22312 406
rect 22284 379 22285 405
rect 22285 379 22311 405
rect 22311 379 22312 405
rect 22284 378 22312 379
rect 22336 405 22364 406
rect 22336 379 22337 405
rect 22337 379 22363 405
rect 22363 379 22364 405
rect 22336 378 22364 379
rect 22302 294 22330 322
rect 22470 686 22498 714
rect 22582 966 22610 994
rect 22582 686 22610 714
rect 22694 1022 22722 1050
rect 22694 518 22722 546
rect 22638 462 22666 490
rect 23478 2534 23506 2562
rect 23086 1918 23114 1946
rect 23254 1694 23282 1722
rect 23086 1049 23114 1050
rect 23086 1023 23087 1049
rect 23087 1023 23113 1049
rect 23113 1023 23114 1049
rect 23086 1022 23114 1023
rect 23478 1134 23506 1162
rect 23422 966 23450 994
rect 22974 742 23002 770
rect 23198 798 23226 826
rect 22974 630 23002 658
rect 22750 294 22778 322
rect 22414 70 22442 98
rect 22526 126 22554 154
rect 22750 70 22778 98
rect 23646 1246 23674 1274
rect 23982 2758 24010 2786
rect 23926 2113 23954 2114
rect 23926 2087 23927 2113
rect 23927 2087 23953 2113
rect 23953 2087 23954 2113
rect 23926 2086 23954 2087
rect 23702 1022 23730 1050
rect 23590 798 23618 826
rect 23646 854 23674 882
rect 23590 182 23618 210
rect 23870 742 23898 770
rect 23926 630 23954 658
rect 26222 7014 26250 7042
rect 26390 7014 26418 7042
rect 25662 6566 25690 6594
rect 25606 6398 25634 6426
rect 25494 6033 25522 6034
rect 25494 6007 25495 6033
rect 25495 6007 25521 6033
rect 25521 6007 25522 6033
rect 25494 6006 25522 6007
rect 25438 5838 25466 5866
rect 24878 3374 24906 3402
rect 24486 3345 24514 3346
rect 24486 3319 24487 3345
rect 24487 3319 24513 3345
rect 24513 3319 24514 3345
rect 24486 3318 24514 3319
rect 24318 2590 24346 2618
rect 24318 2478 24346 2506
rect 24038 2142 24066 2170
rect 24206 2030 24234 2058
rect 24038 910 24066 938
rect 24822 1862 24850 1890
rect 24710 1750 24738 1778
rect 24318 1694 24346 1722
rect 24206 518 24234 546
rect 24318 910 24346 938
rect 24094 238 24122 266
rect 24374 742 24402 770
rect 24374 126 24402 154
rect 24710 966 24738 994
rect 24766 1190 24794 1218
rect 24486 574 24514 602
rect 24542 742 24570 770
rect 24430 70 24458 98
rect 25102 2926 25130 2954
rect 25494 5670 25522 5698
rect 25326 2254 25354 2282
rect 25214 1385 25242 1386
rect 25214 1359 25215 1385
rect 25215 1359 25241 1385
rect 25241 1359 25242 1385
rect 25214 1358 25242 1359
rect 25214 854 25242 882
rect 24766 686 24794 714
rect 24990 798 25018 826
rect 24766 601 24794 602
rect 24766 575 24767 601
rect 24767 575 24793 601
rect 24793 575 24794 601
rect 24766 574 24794 575
rect 24766 182 24794 210
rect 25326 1358 25354 1386
rect 25382 798 25410 826
rect 25438 2030 25466 2058
rect 25270 742 25298 770
rect 25550 2982 25578 3010
rect 25550 2366 25578 2394
rect 27678 7014 27706 7042
rect 27902 7014 27930 7042
rect 26502 6174 26530 6202
rect 25998 5670 26026 5698
rect 25662 5054 25690 5082
rect 25886 5334 25914 5362
rect 25774 4158 25802 4186
rect 25662 3766 25690 3794
rect 25718 2590 25746 2618
rect 25550 1638 25578 1666
rect 25718 2478 25746 2506
rect 25550 1470 25578 1498
rect 25494 854 25522 882
rect 25550 798 25578 826
rect 25438 686 25466 714
rect 25662 1134 25690 1162
rect 25438 462 25466 490
rect 25214 350 25242 378
rect 25550 238 25578 266
rect 25942 5110 25970 5138
rect 25998 4662 26026 4690
rect 26278 5054 26306 5082
rect 25942 3262 25970 3290
rect 26166 4550 26194 4578
rect 25886 2478 25914 2506
rect 26110 3150 26138 3178
rect 25774 1582 25802 1610
rect 25830 1694 25858 1722
rect 25886 937 25914 938
rect 25886 911 25887 937
rect 25887 911 25913 937
rect 25913 911 25914 937
rect 25886 910 25914 911
rect 26222 2310 26250 2338
rect 26222 518 26250 546
rect 26838 6062 26866 6090
rect 26558 5894 26586 5922
rect 26558 4998 26586 5026
rect 26726 5782 26754 5810
rect 29134 7014 29162 7042
rect 29358 7014 29386 7042
rect 28406 6481 28434 6482
rect 28406 6455 28407 6481
rect 28407 6455 28433 6481
rect 28433 6455 28434 6481
rect 28406 6454 28434 6455
rect 31318 6958 31346 6986
rect 30590 6566 30618 6594
rect 31150 6734 31178 6762
rect 31094 6510 31122 6538
rect 29526 6286 29554 6314
rect 28462 6118 28490 6146
rect 27566 6033 27594 6034
rect 27566 6007 27567 6033
rect 27567 6007 27593 6033
rect 27593 6007 27594 6033
rect 27566 6006 27594 6007
rect 27734 6006 27762 6034
rect 26894 5110 26922 5138
rect 27678 5838 27706 5866
rect 27734 5278 27762 5306
rect 27846 5054 27874 5082
rect 27678 3710 27706 3738
rect 26838 3206 26866 3234
rect 27622 3542 27650 3570
rect 26782 2841 26810 2842
rect 26782 2815 26783 2841
rect 26783 2815 26809 2841
rect 26809 2815 26810 2841
rect 26782 2814 26810 2815
rect 27062 2758 27090 2786
rect 27398 2673 27426 2674
rect 27398 2647 27399 2673
rect 27399 2647 27425 2673
rect 27425 2647 27426 2673
rect 27398 2646 27426 2647
rect 27678 3318 27706 3346
rect 27622 2590 27650 2618
rect 27678 2561 27706 2562
rect 27678 2535 27679 2561
rect 27679 2535 27705 2561
rect 27705 2535 27706 2561
rect 27678 2534 27706 2535
rect 26726 2310 26754 2338
rect 26950 2478 26978 2506
rect 26446 1302 26474 1330
rect 26390 1134 26418 1162
rect 26446 182 26474 210
rect 26726 1441 26754 1442
rect 26726 1415 26727 1441
rect 26727 1415 26753 1441
rect 26753 1415 26754 1441
rect 26726 1414 26754 1415
rect 27734 2142 27762 2170
rect 27790 3206 27818 3234
rect 28070 2366 28098 2394
rect 27790 1806 27818 1834
rect 27958 1974 27986 2002
rect 27230 1638 27258 1666
rect 27006 1273 27034 1274
rect 27006 1247 27007 1273
rect 27007 1247 27033 1273
rect 27033 1247 27034 1273
rect 27006 1246 27034 1247
rect 26670 350 26698 378
rect 26782 462 26810 490
rect 29022 6033 29050 6034
rect 29022 6007 29023 6033
rect 29023 6007 29049 6033
rect 29049 6007 29050 6033
rect 29022 6006 29050 6007
rect 29022 5054 29050 5082
rect 28518 2086 28546 2114
rect 28238 1777 28266 1778
rect 28238 1751 28239 1777
rect 28239 1751 28265 1777
rect 28265 1751 28266 1777
rect 28238 1750 28266 1751
rect 28070 1638 28098 1666
rect 27678 1582 27706 1610
rect 27454 294 27482 322
rect 28350 1246 28378 1274
rect 28126 1134 28154 1162
rect 27902 854 27930 882
rect 28518 1022 28546 1050
rect 28574 1750 28602 1778
rect 29358 4494 29386 4522
rect 29582 5110 29610 5138
rect 29414 3990 29442 4018
rect 29638 1862 29666 1890
rect 30814 6454 30842 6482
rect 30254 6342 30282 6370
rect 30590 6062 30618 6090
rect 30086 5894 30114 5922
rect 30758 5894 30786 5922
rect 29862 5726 29890 5754
rect 30142 5697 30170 5698
rect 30142 5671 30143 5697
rect 30143 5671 30169 5697
rect 30169 5671 30170 5697
rect 30142 5670 30170 5671
rect 30646 5641 30674 5642
rect 30646 5615 30647 5641
rect 30647 5615 30673 5641
rect 30673 5615 30674 5641
rect 30646 5614 30674 5615
rect 30254 5166 30282 5194
rect 30646 5166 30674 5194
rect 30534 4969 30562 4970
rect 30534 4943 30535 4969
rect 30535 4943 30561 4969
rect 30561 4943 30562 4969
rect 30534 4942 30562 4943
rect 30142 4913 30170 4914
rect 30142 4887 30143 4913
rect 30143 4887 30169 4913
rect 30169 4887 30170 4913
rect 30142 4886 30170 4887
rect 30254 4774 30282 4802
rect 30758 4633 30786 4634
rect 30758 4607 30759 4633
rect 30759 4607 30785 4633
rect 30785 4607 30786 4633
rect 30758 4606 30786 4607
rect 30478 4129 30506 4130
rect 30478 4103 30479 4129
rect 30479 4103 30505 4129
rect 30505 4103 30506 4129
rect 30478 4102 30506 4103
rect 30254 3681 30282 3682
rect 30254 3655 30255 3681
rect 30255 3655 30281 3681
rect 30281 3655 30282 3681
rect 30254 3654 30282 3655
rect 30142 3262 30170 3290
rect 30646 2926 30674 2954
rect 30142 2702 30170 2730
rect 30534 2561 30562 2562
rect 30534 2535 30535 2561
rect 30535 2535 30561 2561
rect 30561 2535 30562 2561
rect 30534 2534 30562 2535
rect 30254 2169 30282 2170
rect 30254 2143 30255 2169
rect 30255 2143 30281 2169
rect 30281 2143 30282 2169
rect 30254 2142 30282 2143
rect 30142 1833 30170 1834
rect 30142 1807 30143 1833
rect 30143 1807 30169 1833
rect 30169 1807 30170 1833
rect 30142 1806 30170 1807
rect 29190 1134 29218 1162
rect 30254 1385 30282 1386
rect 30254 1359 30255 1385
rect 30255 1359 30281 1385
rect 30281 1359 30282 1385
rect 30254 1358 30282 1359
rect 29582 1190 29610 1218
rect 29302 686 29330 714
rect 29470 462 29498 490
rect 29526 742 29554 770
rect 29918 1049 29946 1050
rect 29918 1023 29919 1049
rect 29919 1023 29945 1049
rect 29945 1023 29946 1049
rect 29918 1022 29946 1023
rect 30142 798 30170 826
rect 30646 1806 30674 1834
rect 30646 1721 30674 1722
rect 30646 1695 30647 1721
rect 30647 1695 30673 1721
rect 30673 1695 30674 1721
rect 30646 1694 30674 1695
rect 30646 1329 30674 1330
rect 30646 1303 30647 1329
rect 30647 1303 30673 1329
rect 30673 1303 30674 1329
rect 30646 1302 30674 1303
rect 30646 881 30674 882
rect 30646 855 30647 881
rect 30647 855 30673 881
rect 30673 855 30674 881
rect 30646 854 30674 855
rect 30590 742 30618 770
rect 29806 238 29834 266
rect 29918 462 29946 490
rect 30758 3374 30786 3402
rect 30926 5390 30954 5418
rect 30926 4830 30954 4858
rect 30926 4046 30954 4074
rect 30926 3345 30954 3346
rect 30926 3319 30927 3345
rect 30927 3319 30953 3345
rect 30953 3319 30954 3345
rect 30926 3318 30954 3319
rect 30926 2617 30954 2618
rect 30926 2591 30927 2617
rect 30927 2591 30953 2617
rect 30953 2591 30954 2617
rect 30926 2590 30954 2591
rect 30926 2310 30954 2338
rect 30926 1638 30954 1666
rect 31094 5726 31122 5754
rect 31094 5222 31122 5250
rect 31262 6593 31290 6594
rect 31262 6567 31263 6593
rect 31263 6567 31289 6593
rect 31289 6567 31290 6593
rect 31262 6566 31290 6567
rect 31150 4942 31178 4970
rect 31094 4662 31122 4690
rect 31542 5390 31570 5418
rect 31374 4942 31402 4970
rect 31318 4606 31346 4634
rect 31430 4718 31458 4746
rect 31374 4494 31402 4522
rect 31094 4382 31122 4410
rect 31430 4270 31458 4298
rect 31542 4046 31570 4074
rect 31094 3934 31122 3962
rect 31430 3822 31458 3850
rect 31430 3598 31458 3626
rect 31542 3150 31570 3178
rect 31094 2870 31122 2898
rect 31318 2702 31346 2730
rect 31262 2534 31290 2562
rect 31094 2422 31122 2450
rect 31262 2254 31290 2282
rect 31542 2478 31570 2506
rect 31430 2030 31458 2058
rect 31318 1694 31346 1722
rect 30982 1134 31010 1162
rect 31542 1582 31570 1610
rect 31318 1358 31346 1386
rect 31094 1078 31122 1106
rect 31374 1302 31402 1330
rect 30702 574 30730 602
rect 31094 518 31122 546
rect 30590 462 30618 490
rect 30086 406 30114 434
rect 31430 1134 31458 1162
rect 31542 910 31570 938
rect 31374 14 31402 42
<< metal3 >>
rect 2921 7014 2926 7042
rect 2954 7014 3150 7042
rect 3178 7014 3183 7042
rect 4377 7014 4382 7042
rect 4410 7014 4606 7042
rect 4634 7014 4639 7042
rect 7289 7014 7294 7042
rect 7322 7014 7518 7042
rect 7546 7014 7551 7042
rect 8745 7014 8750 7042
rect 8778 7014 9142 7042
rect 9170 7014 9175 7042
rect 10201 7014 10206 7042
rect 10234 7014 10598 7042
rect 10626 7014 10631 7042
rect 14569 7014 14574 7042
rect 14602 7014 14798 7042
rect 14826 7014 14831 7042
rect 16025 7014 16030 7042
rect 16058 7014 16254 7042
rect 16282 7014 16287 7042
rect 17481 7014 17486 7042
rect 17514 7014 17766 7042
rect 17794 7014 17799 7042
rect 20393 7014 20398 7042
rect 20426 7014 20622 7042
rect 20650 7014 20655 7042
rect 21849 7014 21854 7042
rect 21882 7014 22078 7042
rect 22106 7014 22111 7042
rect 23305 7014 23310 7042
rect 23338 7014 23534 7042
rect 23562 7014 23567 7042
rect 26217 7014 26222 7042
rect 26250 7014 26390 7042
rect 26418 7014 26423 7042
rect 27673 7014 27678 7042
rect 27706 7014 27902 7042
rect 27930 7014 27935 7042
rect 29129 7014 29134 7042
rect 29162 7014 29358 7042
rect 29386 7014 29391 7042
rect 0 6986 56 7000
rect 32144 6986 32200 7000
rect 0 6958 910 6986
rect 938 6958 943 6986
rect 10481 6958 10486 6986
rect 10514 6958 13566 6986
rect 13594 6958 13599 6986
rect 31313 6958 31318 6986
rect 31346 6958 32200 6986
rect 0 6944 56 6958
rect 32144 6944 32200 6958
rect 10985 6902 10990 6930
rect 11018 6902 15862 6930
rect 15890 6902 15895 6930
rect 5105 6846 5110 6874
rect 5138 6846 24094 6874
rect 24122 6846 24127 6874
rect 2081 6790 2086 6818
rect 2114 6790 9086 6818
rect 9114 6790 9119 6818
rect 12609 6790 12614 6818
rect 12642 6790 15750 6818
rect 15778 6790 15783 6818
rect 15857 6790 15862 6818
rect 15890 6790 16702 6818
rect 16730 6790 16735 6818
rect 0 6762 56 6776
rect 32144 6762 32200 6776
rect 0 6734 798 6762
rect 826 6734 831 6762
rect 3817 6734 3822 6762
rect 3850 6734 17318 6762
rect 17346 6734 17351 6762
rect 31145 6734 31150 6762
rect 31178 6734 32200 6762
rect 0 6720 56 6734
rect 32144 6720 32200 6734
rect 7737 6678 7742 6706
rect 7770 6678 12054 6706
rect 12082 6678 12087 6706
rect 2227 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2369 6678
rect 12227 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12369 6678
rect 22227 6650 22232 6678
rect 22260 6650 22284 6678
rect 22312 6650 22336 6678
rect 22364 6650 22369 6678
rect 6729 6622 6734 6650
rect 6762 6622 10262 6650
rect 10290 6622 10295 6650
rect 4186 6566 7014 6594
rect 7042 6566 7047 6594
rect 7289 6566 7294 6594
rect 7322 6566 25662 6594
rect 25690 6566 25695 6594
rect 30585 6566 30590 6594
rect 30618 6566 31262 6594
rect 31290 6566 31295 6594
rect 0 6538 56 6552
rect 4186 6538 4214 6566
rect 32144 6538 32200 6552
rect 0 6510 4214 6538
rect 5833 6510 5838 6538
rect 5866 6510 6454 6538
rect 6482 6510 6487 6538
rect 6897 6510 6902 6538
rect 6930 6510 7238 6538
rect 7266 6510 7271 6538
rect 7345 6510 7350 6538
rect 7378 6510 8918 6538
rect 8946 6510 8951 6538
rect 11657 6510 11662 6538
rect 11690 6510 12222 6538
rect 12250 6510 12255 6538
rect 15946 6510 18438 6538
rect 18466 6510 18471 6538
rect 31089 6510 31094 6538
rect 31122 6510 32200 6538
rect 0 6496 56 6510
rect 15946 6482 15974 6510
rect 32144 6496 32200 6510
rect 1745 6454 1750 6482
rect 1778 6454 7462 6482
rect 7490 6454 7495 6482
rect 9921 6454 9926 6482
rect 9954 6454 10318 6482
rect 10346 6454 10351 6482
rect 11041 6454 11046 6482
rect 11074 6454 11942 6482
rect 11970 6454 11975 6482
rect 12049 6454 12054 6482
rect 12082 6454 15974 6482
rect 16753 6454 16758 6482
rect 16786 6454 17486 6482
rect 17514 6454 17519 6482
rect 18265 6454 18270 6482
rect 18298 6454 19222 6482
rect 19250 6454 19255 6482
rect 28401 6454 28406 6482
rect 28434 6454 30814 6482
rect 30842 6454 30847 6482
rect 6841 6398 6846 6426
rect 6874 6398 25606 6426
rect 25634 6398 25639 6426
rect 3649 6342 3654 6370
rect 3682 6342 10486 6370
rect 10514 6342 10519 6370
rect 10593 6342 10598 6370
rect 10626 6342 14294 6370
rect 14322 6342 14327 6370
rect 16809 6342 16814 6370
rect 16842 6342 30254 6370
rect 30282 6342 30287 6370
rect 0 6314 56 6328
rect 32144 6314 32200 6328
rect 0 6286 1834 6314
rect 6785 6286 6790 6314
rect 6818 6286 11718 6314
rect 11746 6286 11751 6314
rect 12105 6286 12110 6314
rect 12138 6286 16534 6314
rect 16562 6286 16567 6314
rect 29521 6286 29526 6314
rect 29554 6286 32200 6314
rect 0 6272 56 6286
rect 1806 6202 1834 6286
rect 1897 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2039 6286
rect 11897 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12039 6286
rect 21897 6258 21902 6286
rect 21930 6258 21954 6286
rect 21982 6258 22006 6286
rect 22034 6258 22039 6286
rect 32144 6272 32200 6286
rect 12105 6230 12110 6258
rect 12138 6230 12726 6258
rect 12754 6230 12759 6258
rect 13785 6230 13790 6258
rect 13818 6230 16646 6258
rect 16674 6230 16679 6258
rect 1806 6174 5838 6202
rect 5866 6174 5871 6202
rect 8745 6174 8750 6202
rect 8778 6174 26502 6202
rect 26530 6174 26535 6202
rect 6505 6118 6510 6146
rect 6538 6118 18606 6146
rect 18634 6118 18639 6146
rect 24033 6118 24038 6146
rect 24066 6118 28462 6146
rect 28490 6118 28495 6146
rect 0 6090 56 6104
rect 32144 6090 32200 6104
rect 0 6062 2086 6090
rect 2114 6062 2119 6090
rect 8353 6062 8358 6090
rect 8386 6062 20846 6090
rect 20874 6062 20879 6090
rect 21121 6062 21126 6090
rect 21154 6062 26838 6090
rect 26866 6062 26871 6090
rect 30585 6062 30590 6090
rect 30618 6062 32200 6090
rect 0 6048 56 6062
rect 32144 6048 32200 6062
rect 11769 6006 11774 6034
rect 11802 6006 14238 6034
rect 14266 6006 14271 6034
rect 16753 6006 16758 6034
rect 16786 6006 17206 6034
rect 17234 6006 17239 6034
rect 18881 6006 18886 6034
rect 18914 6006 25214 6034
rect 25489 6006 25494 6034
rect 25522 6006 27566 6034
rect 27594 6006 27599 6034
rect 27729 6006 27734 6034
rect 27762 6006 29022 6034
rect 29050 6006 29055 6034
rect 8913 5950 8918 5978
rect 8946 5950 12474 5978
rect 13449 5950 13454 5978
rect 13482 5950 17514 5978
rect 18769 5950 18774 5978
rect 18802 5950 20398 5978
rect 20426 5950 20431 5978
rect 20953 5950 20958 5978
rect 20986 5950 22722 5978
rect 5441 5894 5446 5922
rect 5474 5894 6930 5922
rect 10089 5894 10094 5922
rect 10122 5894 12110 5922
rect 12138 5894 12143 5922
rect 0 5866 56 5880
rect 2227 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2369 5894
rect 6902 5866 6930 5894
rect 12227 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12369 5894
rect 12446 5866 12474 5950
rect 12721 5894 12726 5922
rect 12754 5894 14798 5922
rect 14826 5894 14831 5922
rect 17486 5866 17514 5950
rect 17593 5894 17598 5922
rect 17626 5894 19054 5922
rect 19082 5894 19087 5922
rect 22227 5866 22232 5894
rect 22260 5866 22284 5894
rect 22312 5866 22336 5894
rect 22364 5866 22369 5894
rect 22694 5866 22722 5950
rect 25186 5922 25214 6006
rect 25186 5894 25578 5922
rect 26553 5894 26558 5922
rect 26586 5894 30086 5922
rect 30114 5894 30119 5922
rect 30753 5894 30758 5922
rect 30786 5894 31402 5922
rect 25550 5866 25578 5894
rect 31374 5866 31402 5894
rect 32144 5866 32200 5880
rect 0 5838 2086 5866
rect 2114 5838 2119 5866
rect 4186 5838 6790 5866
rect 6818 5838 6823 5866
rect 6902 5838 11774 5866
rect 11802 5838 11807 5866
rect 12446 5838 13342 5866
rect 13370 5838 13375 5866
rect 17486 5838 18494 5866
rect 18522 5838 18527 5866
rect 22694 5838 25438 5866
rect 25466 5838 25471 5866
rect 25550 5838 27678 5866
rect 27706 5838 27711 5866
rect 31374 5838 32200 5866
rect 0 5824 56 5838
rect 4186 5810 4214 5838
rect 32144 5824 32200 5838
rect 905 5782 910 5810
rect 938 5782 4214 5810
rect 5833 5782 5838 5810
rect 5866 5782 13454 5810
rect 13482 5782 13487 5810
rect 14961 5782 14966 5810
rect 14994 5782 26726 5810
rect 26754 5782 26759 5810
rect 8241 5726 8246 5754
rect 8274 5726 12166 5754
rect 12194 5726 12199 5754
rect 12273 5726 12278 5754
rect 12306 5726 12950 5754
rect 12978 5726 12983 5754
rect 15297 5726 15302 5754
rect 15330 5726 16198 5754
rect 16226 5726 16231 5754
rect 16697 5726 16702 5754
rect 16730 5726 20958 5754
rect 20986 5726 20991 5754
rect 29857 5726 29862 5754
rect 29890 5726 31094 5754
rect 31122 5726 31127 5754
rect 793 5670 798 5698
rect 826 5670 10178 5698
rect 10929 5670 10934 5698
rect 10962 5670 12446 5698
rect 12474 5670 12479 5698
rect 12553 5670 12558 5698
rect 12586 5670 18382 5698
rect 18410 5670 18415 5698
rect 21793 5670 21798 5698
rect 21826 5670 25494 5698
rect 25522 5670 25527 5698
rect 25993 5670 25998 5698
rect 26026 5670 30142 5698
rect 30170 5670 30175 5698
rect 0 5642 56 5656
rect 10150 5642 10178 5670
rect 32144 5642 32200 5656
rect 0 5614 7574 5642
rect 10150 5614 12782 5642
rect 12810 5614 12815 5642
rect 14233 5614 14238 5642
rect 14266 5614 16422 5642
rect 16450 5614 16455 5642
rect 19721 5614 19726 5642
rect 19754 5614 23534 5642
rect 23562 5614 23567 5642
rect 30641 5614 30646 5642
rect 30674 5614 32200 5642
rect 0 5600 56 5614
rect 7546 5586 7574 5614
rect 32144 5600 32200 5614
rect 2081 5558 2086 5586
rect 2114 5558 7238 5586
rect 7266 5558 7271 5586
rect 7546 5558 10598 5586
rect 10626 5558 10631 5586
rect 11713 5558 11718 5586
rect 11746 5558 15974 5586
rect 18713 5558 18718 5586
rect 18746 5558 22638 5586
rect 22666 5558 22671 5586
rect 15946 5530 15974 5558
rect 12105 5502 12110 5530
rect 12138 5502 13454 5530
rect 13482 5502 13487 5530
rect 13561 5502 13566 5530
rect 13594 5502 15806 5530
rect 15834 5502 15839 5530
rect 15946 5502 21742 5530
rect 21770 5502 21775 5530
rect 1897 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2039 5502
rect 11897 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12039 5502
rect 21897 5474 21902 5502
rect 21930 5474 21954 5502
rect 21982 5474 22006 5502
rect 22034 5474 22039 5502
rect 9137 5446 9142 5474
rect 9170 5446 10934 5474
rect 10962 5446 10967 5474
rect 12161 5446 12166 5474
rect 12194 5446 14126 5474
rect 14154 5446 14159 5474
rect 18433 5446 18438 5474
rect 18466 5446 21518 5474
rect 21546 5446 21551 5474
rect 0 5418 56 5432
rect 32144 5418 32200 5432
rect 0 5390 12614 5418
rect 12642 5390 12647 5418
rect 15689 5390 15694 5418
rect 15722 5390 30926 5418
rect 30954 5390 30959 5418
rect 31537 5390 31542 5418
rect 31570 5390 32200 5418
rect 0 5376 56 5390
rect 32144 5376 32200 5390
rect 9081 5334 9086 5362
rect 9114 5334 11158 5362
rect 11186 5334 11191 5362
rect 11321 5334 11326 5362
rect 11354 5334 25886 5362
rect 25914 5334 25919 5362
rect 2809 5278 2814 5306
rect 2842 5278 14686 5306
rect 14714 5278 14719 5306
rect 16753 5278 16758 5306
rect 16786 5278 22526 5306
rect 22554 5278 22559 5306
rect 22633 5278 22638 5306
rect 22666 5278 27734 5306
rect 27762 5278 27767 5306
rect 7121 5222 7126 5250
rect 7154 5222 12110 5250
rect 12138 5222 12143 5250
rect 12217 5222 12222 5250
rect 12250 5222 14238 5250
rect 14266 5222 14271 5250
rect 14961 5222 14966 5250
rect 14994 5222 31094 5250
rect 31122 5222 31127 5250
rect 0 5194 56 5208
rect 32144 5194 32200 5208
rect 0 5166 10038 5194
rect 10066 5166 10071 5194
rect 10990 5166 13398 5194
rect 13426 5166 13431 5194
rect 14849 5166 14854 5194
rect 14882 5166 15638 5194
rect 15666 5166 15671 5194
rect 15946 5166 22442 5194
rect 22521 5166 22526 5194
rect 22554 5166 30254 5194
rect 30282 5166 30287 5194
rect 30641 5166 30646 5194
rect 30674 5166 32200 5194
rect 0 5152 56 5166
rect 4209 5110 4214 5138
rect 4242 5110 7686 5138
rect 7714 5110 7719 5138
rect 2227 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2369 5110
rect 7350 5054 9982 5082
rect 10010 5054 10015 5082
rect 10201 5054 10206 5082
rect 10234 5054 10878 5082
rect 10906 5054 10911 5082
rect 7350 5026 7378 5054
rect 10990 5026 11018 5166
rect 11097 5110 11102 5138
rect 11130 5110 12166 5138
rect 12194 5110 12199 5138
rect 12441 5110 12446 5138
rect 12474 5110 15190 5138
rect 15218 5110 15223 5138
rect 15913 5110 15918 5138
rect 15946 5110 15974 5166
rect 22414 5138 22442 5166
rect 32144 5152 32200 5166
rect 22414 5110 25942 5138
rect 25970 5110 25975 5138
rect 26889 5110 26894 5138
rect 26922 5110 29582 5138
rect 29610 5110 29615 5138
rect 12227 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12369 5110
rect 22227 5082 22232 5110
rect 22260 5082 22284 5110
rect 22312 5082 22336 5110
rect 22364 5082 22369 5110
rect 12670 5054 16310 5082
rect 16338 5054 16343 5082
rect 16865 5054 16870 5082
rect 16898 5054 19446 5082
rect 19474 5054 19479 5082
rect 25657 5054 25662 5082
rect 25690 5054 26278 5082
rect 26306 5054 26311 5082
rect 27841 5054 27846 5082
rect 27874 5054 29022 5082
rect 29050 5054 29055 5082
rect 6673 4998 6678 5026
rect 6706 4998 7378 5026
rect 7457 4998 7462 5026
rect 7490 4998 11018 5026
rect 11153 4998 11158 5026
rect 11186 4998 12558 5026
rect 12586 4998 12591 5026
rect 0 4970 56 4984
rect 0 4942 7154 4970
rect 7233 4942 7238 4970
rect 7266 4942 7574 4970
rect 7602 4942 7607 4970
rect 7681 4942 7686 4970
rect 7714 4942 12334 4970
rect 12362 4942 12367 4970
rect 0 4928 56 4942
rect 7126 4914 7154 4942
rect 12670 4914 12698 5054
rect 13449 4998 13454 5026
rect 13482 4998 14686 5026
rect 14714 4998 14719 5026
rect 18713 4998 18718 5026
rect 18746 4998 26558 5026
rect 26586 4998 26591 5026
rect 32144 4970 32200 4984
rect 12777 4942 12782 4970
rect 12810 4942 16758 4970
rect 16786 4942 16791 4970
rect 18377 4942 18382 4970
rect 18410 4942 21798 4970
rect 21826 4942 21831 4970
rect 30529 4942 30534 4970
rect 30562 4942 31150 4970
rect 31178 4942 31183 4970
rect 31369 4942 31374 4970
rect 31402 4942 32200 4970
rect 32144 4928 32200 4942
rect 4153 4886 4158 4914
rect 4186 4886 6790 4914
rect 6818 4886 6823 4914
rect 7126 4886 9086 4914
rect 9114 4886 9119 4914
rect 9193 4886 9198 4914
rect 9226 4886 12698 4914
rect 13057 4886 13062 4914
rect 13090 4886 30142 4914
rect 30170 4886 30175 4914
rect 3929 4830 3934 4858
rect 3962 4830 8302 4858
rect 8330 4830 8335 4858
rect 10066 4830 15974 4858
rect 16002 4830 16007 4858
rect 22073 4830 22078 4858
rect 22106 4830 23618 4858
rect 24089 4830 24094 4858
rect 24122 4830 30926 4858
rect 30954 4830 30959 4858
rect 10066 4802 10094 4830
rect 23590 4802 23618 4830
rect 2081 4774 2086 4802
rect 2114 4774 6734 4802
rect 6762 4774 6767 4802
rect 7401 4774 7406 4802
rect 7434 4774 10094 4802
rect 11214 4774 12110 4802
rect 12138 4774 12143 4802
rect 12273 4774 12278 4802
rect 12306 4774 14014 4802
rect 14042 4774 14047 4802
rect 16305 4774 16310 4802
rect 16338 4774 19558 4802
rect 19586 4774 19591 4802
rect 20281 4774 20286 4802
rect 20314 4774 22414 4802
rect 22442 4774 22447 4802
rect 23590 4774 30254 4802
rect 30282 4774 30287 4802
rect 0 4746 56 4760
rect 0 4718 1834 4746
rect 4265 4718 4270 4746
rect 4298 4718 8358 4746
rect 8386 4718 8391 4746
rect 8857 4718 8862 4746
rect 8890 4718 11102 4746
rect 11130 4718 11135 4746
rect 0 4704 56 4718
rect 1806 4634 1834 4718
rect 1897 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2039 4718
rect 11214 4690 11242 4774
rect 32144 4746 32200 4760
rect 12110 4718 18270 4746
rect 18298 4718 18303 4746
rect 31425 4718 31430 4746
rect 31458 4718 32200 4746
rect 11897 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12039 4718
rect 7569 4662 7574 4690
rect 7602 4662 11242 4690
rect 1806 4606 7462 4634
rect 7490 4606 7495 4634
rect 8353 4606 8358 4634
rect 8386 4606 11662 4634
rect 11690 4606 11695 4634
rect 12110 4578 12138 4718
rect 21897 4690 21902 4718
rect 21930 4690 21954 4718
rect 21982 4690 22006 4718
rect 22034 4690 22039 4718
rect 32144 4704 32200 4718
rect 12833 4662 12838 4690
rect 12866 4662 15974 4690
rect 16753 4662 16758 4690
rect 16786 4662 20118 4690
rect 20146 4662 20151 4690
rect 22078 4662 25998 4690
rect 26026 4662 26031 4690
rect 28126 4662 31094 4690
rect 31122 4662 31127 4690
rect 15946 4634 15974 4662
rect 12329 4606 12334 4634
rect 12362 4606 14182 4634
rect 14210 4606 14215 4634
rect 15946 4606 21966 4634
rect 21994 4606 21999 4634
rect 22078 4578 22106 4662
rect 28126 4634 28154 4662
rect 22409 4606 22414 4634
rect 22442 4606 28154 4634
rect 30753 4606 30758 4634
rect 30786 4606 31318 4634
rect 31346 4606 31351 4634
rect 6785 4550 6790 4578
rect 6818 4550 10318 4578
rect 10346 4550 10351 4578
rect 10425 4550 10430 4578
rect 10458 4550 12138 4578
rect 12273 4550 12278 4578
rect 12306 4550 14210 4578
rect 14513 4550 14518 4578
rect 14546 4550 22106 4578
rect 22185 4550 22190 4578
rect 22218 4550 26166 4578
rect 26194 4550 26199 4578
rect 0 4522 56 4536
rect 14182 4522 14210 4550
rect 32144 4522 32200 4536
rect 0 4494 7518 4522
rect 7546 4494 7551 4522
rect 8017 4494 8022 4522
rect 8050 4494 10654 4522
rect 10682 4494 10687 4522
rect 10929 4494 10934 4522
rect 10962 4494 14070 4522
rect 14098 4494 14103 4522
rect 14182 4494 15134 4522
rect 15162 4494 15167 4522
rect 15946 4494 16926 4522
rect 16954 4494 16959 4522
rect 17257 4494 17262 4522
rect 17290 4494 29358 4522
rect 29386 4494 29391 4522
rect 31369 4494 31374 4522
rect 31402 4494 32200 4522
rect 0 4480 56 4494
rect 15946 4466 15974 4494
rect 32144 4480 32200 4494
rect 961 4438 966 4466
rect 994 4438 7042 4466
rect 7121 4438 7126 4466
rect 7154 4438 7462 4466
rect 7490 4438 7495 4466
rect 7569 4438 7574 4466
rect 7602 4438 10094 4466
rect 10122 4438 10127 4466
rect 10425 4438 10430 4466
rect 10458 4438 10463 4466
rect 10537 4438 10542 4466
rect 10570 4438 12278 4466
rect 12306 4438 12311 4466
rect 12441 4438 12446 4466
rect 12474 4438 15974 4466
rect 16025 4438 16030 4466
rect 16058 4438 18494 4466
rect 18522 4438 18527 4466
rect 19441 4438 19446 4466
rect 19474 4438 24094 4466
rect 24122 4438 24127 4466
rect 7014 4410 7042 4438
rect 1241 4382 1246 4410
rect 1274 4382 4214 4410
rect 7014 4382 9198 4410
rect 9226 4382 9231 4410
rect 4186 4354 4214 4382
rect 10430 4354 10458 4438
rect 4186 4326 7350 4354
rect 7378 4326 7383 4354
rect 7457 4326 7462 4354
rect 7490 4326 10458 4354
rect 10486 4382 16982 4410
rect 17010 4382 17015 4410
rect 19161 4382 19166 4410
rect 19194 4382 31094 4410
rect 31122 4382 31127 4410
rect 0 4298 56 4312
rect 2227 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2369 4326
rect 10486 4298 10514 4382
rect 10649 4326 10654 4354
rect 10682 4326 12166 4354
rect 12194 4326 12199 4354
rect 13337 4326 13342 4354
rect 13370 4326 16758 4354
rect 16786 4326 16791 4354
rect 16921 4326 16926 4354
rect 16954 4326 17542 4354
rect 17570 4326 17575 4354
rect 18433 4326 18438 4354
rect 18466 4326 20566 4354
rect 20594 4326 20599 4354
rect 12227 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12369 4326
rect 22227 4298 22232 4326
rect 22260 4298 22284 4326
rect 22312 4298 22336 4326
rect 22364 4298 22369 4326
rect 32144 4298 32200 4312
rect 0 4270 2086 4298
rect 2114 4270 2119 4298
rect 7009 4270 7014 4298
rect 7042 4270 10514 4298
rect 10593 4270 10598 4298
rect 10626 4270 12110 4298
rect 12138 4270 12143 4298
rect 12721 4270 12726 4298
rect 12754 4270 16758 4298
rect 16786 4270 16791 4298
rect 16865 4270 16870 4298
rect 16898 4270 18886 4298
rect 18914 4270 18919 4298
rect 31425 4270 31430 4298
rect 31458 4270 32200 4298
rect 0 4256 56 4270
rect 32144 4256 32200 4270
rect 7457 4214 7462 4242
rect 7490 4214 8862 4242
rect 8890 4214 8895 4242
rect 10033 4214 10038 4242
rect 10066 4214 10962 4242
rect 11041 4214 11046 4242
rect 11074 4214 12614 4242
rect 12642 4214 12647 4242
rect 13001 4214 13006 4242
rect 13034 4214 14910 4242
rect 14938 4214 14943 4242
rect 15078 4214 19306 4242
rect 19665 4214 19670 4242
rect 19698 4214 22414 4242
rect 22442 4214 22447 4242
rect 10934 4186 10962 4214
rect 15078 4186 15106 4214
rect 19278 4186 19306 4214
rect 7513 4158 7518 4186
rect 7546 4158 10822 4186
rect 10850 4158 10855 4186
rect 10934 4158 12502 4186
rect 12530 4158 12535 4186
rect 13393 4158 13398 4186
rect 13426 4158 15106 4186
rect 15969 4158 15974 4186
rect 16002 4158 16954 4186
rect 19278 4158 20958 4186
rect 20986 4158 20991 4186
rect 21065 4158 21070 4186
rect 21098 4158 25774 4186
rect 25802 4158 25807 4186
rect 16926 4130 16954 4158
rect 7513 4102 7518 4130
rect 7546 4102 12782 4130
rect 12810 4102 12815 4130
rect 13426 4102 13678 4130
rect 13706 4102 13711 4130
rect 14177 4102 14182 4130
rect 14210 4102 16814 4130
rect 16842 4102 16847 4130
rect 16926 4102 30478 4130
rect 30506 4102 30511 4130
rect 0 4074 56 4088
rect 13426 4074 13454 4102
rect 32144 4074 32200 4088
rect 0 4046 10598 4074
rect 10626 4046 10631 4074
rect 10710 4046 13454 4074
rect 15129 4046 15134 4074
rect 15162 4046 18438 4074
rect 18466 4046 18471 4074
rect 18886 4046 22274 4074
rect 22913 4046 22918 4074
rect 22946 4046 30926 4074
rect 30954 4046 30959 4074
rect 31537 4046 31542 4074
rect 31570 4046 32200 4074
rect 0 4032 56 4046
rect 1521 3990 1526 4018
rect 1554 3990 4214 4018
rect 4242 3990 4247 4018
rect 5609 3990 5614 4018
rect 5642 3990 10542 4018
rect 10570 3990 10575 4018
rect 10710 3962 10738 4046
rect 18886 4018 18914 4046
rect 22246 4018 22274 4046
rect 32144 4032 32200 4046
rect 11937 3990 11942 4018
rect 11970 3990 12894 4018
rect 12922 3990 12927 4018
rect 13841 3990 13846 4018
rect 13874 3990 18914 4018
rect 19306 3990 22162 4018
rect 22246 3990 29414 4018
rect 29442 3990 29447 4018
rect 19306 3962 19334 3990
rect 6617 3934 6622 3962
rect 6650 3934 8414 3962
rect 8442 3934 8447 3962
rect 9977 3934 9982 3962
rect 10010 3934 10738 3962
rect 13393 3934 13398 3962
rect 13426 3934 19334 3962
rect 22134 3962 22162 3990
rect 22134 3934 31094 3962
rect 31122 3934 31127 3962
rect 1897 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2039 3934
rect 11897 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12039 3934
rect 21897 3906 21902 3934
rect 21930 3906 21954 3934
rect 21982 3906 22006 3934
rect 22034 3906 22039 3934
rect 6113 3878 6118 3906
rect 6146 3878 10598 3906
rect 10626 3878 10631 3906
rect 14121 3878 14126 3906
rect 14154 3878 17570 3906
rect 17761 3878 17766 3906
rect 17794 3878 21070 3906
rect 21098 3878 21103 3906
rect 0 3850 56 3864
rect 0 3822 7238 3850
rect 7266 3822 7271 3850
rect 7513 3822 7518 3850
rect 7546 3822 10430 3850
rect 10458 3822 10463 3850
rect 10649 3822 10654 3850
rect 10682 3822 12726 3850
rect 12754 3822 12759 3850
rect 15073 3822 15078 3850
rect 15106 3822 15974 3850
rect 16002 3822 16007 3850
rect 0 3808 56 3822
rect 17542 3794 17570 3878
rect 32144 3850 32200 3864
rect 18494 3822 20342 3850
rect 20370 3822 20375 3850
rect 20673 3822 20678 3850
rect 20706 3822 22918 3850
rect 22946 3822 22951 3850
rect 31425 3822 31430 3850
rect 31458 3822 32200 3850
rect 18494 3794 18522 3822
rect 32144 3808 32200 3822
rect 1633 3766 1638 3794
rect 1666 3766 5614 3794
rect 5642 3766 5647 3794
rect 6841 3766 6846 3794
rect 6874 3766 12446 3794
rect 12474 3766 12479 3794
rect 13057 3766 13062 3794
rect 13090 3766 14966 3794
rect 14994 3766 14999 3794
rect 17542 3766 18522 3794
rect 20897 3766 20902 3794
rect 20930 3766 25662 3794
rect 25690 3766 25695 3794
rect 4433 3710 4438 3738
rect 4466 3710 7518 3738
rect 7546 3710 7551 3738
rect 10593 3710 10598 3738
rect 10626 3710 14126 3738
rect 14154 3710 14159 3738
rect 15017 3710 15022 3738
rect 15050 3710 27678 3738
rect 27706 3710 27711 3738
rect 6729 3654 6734 3682
rect 6762 3654 8358 3682
rect 8386 3654 8391 3682
rect 10425 3654 10430 3682
rect 10458 3654 13790 3682
rect 13818 3654 13823 3682
rect 13953 3654 13958 3682
rect 13986 3654 30254 3682
rect 30282 3654 30287 3682
rect 0 3626 56 3640
rect 32144 3626 32200 3640
rect 0 3598 7462 3626
rect 7490 3598 7495 3626
rect 8409 3598 8414 3626
rect 8442 3598 9898 3626
rect 10425 3598 10430 3626
rect 10458 3598 20790 3626
rect 20818 3598 20823 3626
rect 31425 3598 31430 3626
rect 31458 3598 32200 3626
rect 0 3584 56 3598
rect 9870 3570 9898 3598
rect 32144 3584 32200 3598
rect 2921 3542 2926 3570
rect 2954 3542 9758 3570
rect 9786 3542 9791 3570
rect 9870 3542 10990 3570
rect 11018 3542 11023 3570
rect 12721 3542 12726 3570
rect 12754 3542 14434 3570
rect 16809 3542 16814 3570
rect 16842 3542 18382 3570
rect 18410 3542 18415 3570
rect 23529 3542 23534 3570
rect 23562 3542 27622 3570
rect 27650 3542 27655 3570
rect 2227 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2369 3542
rect 12227 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12369 3542
rect 14406 3514 14434 3542
rect 22227 3514 22232 3542
rect 22260 3514 22284 3542
rect 22312 3514 22336 3542
rect 22364 3514 22369 3542
rect 4713 3486 4718 3514
rect 4746 3486 9198 3514
rect 9226 3486 9231 3514
rect 9366 3486 11830 3514
rect 11858 3486 11863 3514
rect 12446 3486 14294 3514
rect 14322 3486 14327 3514
rect 14406 3486 17766 3514
rect 17794 3486 17799 3514
rect 9366 3458 9394 3486
rect 12446 3458 12474 3486
rect 4186 3430 6678 3458
rect 6706 3430 6711 3458
rect 6790 3430 9394 3458
rect 9865 3430 9870 3458
rect 9898 3430 12474 3458
rect 12665 3430 12670 3458
rect 12698 3430 12978 3458
rect 13337 3430 13342 3458
rect 13370 3430 16758 3458
rect 16786 3430 16791 3458
rect 0 3402 56 3416
rect 4186 3402 4214 3430
rect 6790 3402 6818 3430
rect 12950 3402 12978 3430
rect 32144 3402 32200 3416
rect 0 3374 4214 3402
rect 4825 3374 4830 3402
rect 4858 3374 6818 3402
rect 7681 3374 7686 3402
rect 7714 3374 9282 3402
rect 10705 3374 10710 3402
rect 10738 3374 11774 3402
rect 11802 3374 11807 3402
rect 12105 3374 12110 3402
rect 12138 3374 12838 3402
rect 12866 3374 12871 3402
rect 12950 3374 13482 3402
rect 14905 3374 14910 3402
rect 14938 3374 15582 3402
rect 15610 3374 15615 3402
rect 16697 3374 16702 3402
rect 16730 3374 17682 3402
rect 18153 3374 18158 3402
rect 18186 3374 21686 3402
rect 21714 3374 21719 3402
rect 22689 3374 22694 3402
rect 22722 3374 24878 3402
rect 24906 3374 24911 3402
rect 30753 3374 30758 3402
rect 30786 3374 32200 3402
rect 0 3360 56 3374
rect 9254 3346 9282 3374
rect 13454 3346 13482 3374
rect 17654 3346 17682 3374
rect 32144 3360 32200 3374
rect 3929 3318 3934 3346
rect 3962 3318 6370 3346
rect 6449 3318 6454 3346
rect 6482 3318 8246 3346
rect 8274 3318 8279 3346
rect 9249 3318 9254 3346
rect 9282 3318 9287 3346
rect 10257 3318 10262 3346
rect 10290 3318 13342 3346
rect 13370 3318 13375 3346
rect 13454 3318 15358 3346
rect 15386 3318 15391 3346
rect 17654 3318 18914 3346
rect 20113 3318 20118 3346
rect 20146 3318 24486 3346
rect 24514 3318 24519 3346
rect 27673 3318 27678 3346
rect 27706 3318 30926 3346
rect 30954 3318 30959 3346
rect 6342 3234 6370 3318
rect 6673 3262 6678 3290
rect 6706 3262 11550 3290
rect 11578 3262 11583 3290
rect 12105 3262 12110 3290
rect 12138 3262 13118 3290
rect 13146 3262 13151 3290
rect 13225 3262 13230 3290
rect 13258 3262 16030 3290
rect 16058 3262 16063 3290
rect 18886 3234 18914 3318
rect 20785 3262 20790 3290
rect 20818 3262 22694 3290
rect 22722 3262 22727 3290
rect 25937 3262 25942 3290
rect 25970 3262 30142 3290
rect 30170 3262 30175 3290
rect 1806 3206 4242 3234
rect 6342 3206 7238 3234
rect 7266 3206 7271 3234
rect 8857 3206 8862 3234
rect 8890 3206 12138 3234
rect 12665 3206 12670 3234
rect 12698 3206 14854 3234
rect 14882 3206 14887 3234
rect 15185 3206 15190 3234
rect 15218 3206 18438 3234
rect 18466 3206 18471 3234
rect 18886 3206 22526 3234
rect 22554 3206 22559 3234
rect 26833 3206 26838 3234
rect 26866 3206 27790 3234
rect 27818 3206 27823 3234
rect 0 3178 56 3192
rect 1806 3178 1834 3206
rect 0 3150 1834 3178
rect 4214 3178 4242 3206
rect 4214 3150 4410 3178
rect 0 3136 56 3150
rect 1897 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2039 3150
rect 4382 3066 4410 3150
rect 7350 3150 11326 3178
rect 11354 3150 11359 3178
rect 7350 3122 7378 3150
rect 11897 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12039 3150
rect 12110 3122 12138 3206
rect 32144 3178 32200 3192
rect 12609 3150 12614 3178
rect 12642 3150 18158 3178
rect 18186 3150 18191 3178
rect 18377 3150 18382 3178
rect 18410 3150 20398 3178
rect 20426 3150 20431 3178
rect 22409 3150 22414 3178
rect 22442 3150 26110 3178
rect 26138 3150 26143 3178
rect 31537 3150 31542 3178
rect 31570 3150 32200 3178
rect 21897 3122 21902 3150
rect 21930 3122 21954 3150
rect 21982 3122 22006 3150
rect 22034 3122 22039 3150
rect 32144 3136 32200 3150
rect 4601 3094 4606 3122
rect 4634 3094 7378 3122
rect 9081 3094 9086 3122
rect 9114 3094 10038 3122
rect 10066 3094 10071 3122
rect 12110 3094 13454 3122
rect 14009 3094 14014 3122
rect 14042 3094 18914 3122
rect 22577 3094 22582 3122
rect 22610 3094 24430 3122
rect 24458 3094 24463 3122
rect 13426 3066 13454 3094
rect 18886 3066 18914 3094
rect 345 3038 350 3066
rect 378 3038 4270 3066
rect 4298 3038 4303 3066
rect 4382 3038 6734 3066
rect 6762 3038 6767 3066
rect 8073 3038 8078 3066
rect 8106 3038 12614 3066
rect 12642 3038 12647 3066
rect 13426 3038 14182 3066
rect 14210 3038 14215 3066
rect 14793 3038 14798 3066
rect 14826 3038 18858 3066
rect 18886 3038 23422 3066
rect 23450 3038 23455 3066
rect 6566 2982 7574 3010
rect 9249 2982 9254 3010
rect 9282 2982 16758 3010
rect 16786 2982 16791 3010
rect 0 2954 56 2968
rect 0 2926 6454 2954
rect 6482 2926 6487 2954
rect 0 2912 56 2926
rect 6566 2898 6594 2982
rect 7546 2954 7574 2982
rect 18830 2954 18858 3038
rect 20841 2982 20846 3010
rect 20874 2982 25550 3010
rect 25578 2982 25583 3010
rect 32144 2954 32200 2968
rect 7546 2926 9926 2954
rect 9954 2926 9959 2954
rect 10369 2926 10374 2954
rect 10402 2926 12670 2954
rect 12698 2926 12703 2954
rect 12889 2926 12894 2954
rect 12922 2926 15974 2954
rect 18830 2926 25102 2954
rect 25130 2926 25135 2954
rect 30641 2926 30646 2954
rect 30674 2926 32200 2954
rect 15946 2898 15974 2926
rect 32144 2912 32200 2926
rect 2641 2870 2646 2898
rect 2674 2870 6594 2898
rect 6729 2870 6734 2898
rect 6762 2870 9142 2898
rect 9170 2870 9175 2898
rect 10929 2870 10934 2898
rect 10962 2870 15078 2898
rect 15106 2870 15111 2898
rect 15946 2870 31094 2898
rect 31122 2870 31127 2898
rect 2417 2814 2422 2842
rect 2450 2814 9870 2842
rect 9898 2814 9903 2842
rect 10593 2814 10598 2842
rect 10626 2814 14350 2842
rect 14378 2814 14383 2842
rect 16137 2814 16142 2842
rect 16170 2814 26782 2842
rect 26810 2814 26815 2842
rect 7065 2758 7070 2786
rect 7098 2758 10486 2786
rect 10514 2758 10519 2786
rect 12777 2758 12782 2786
rect 12810 2758 22134 2786
rect 22162 2758 22167 2786
rect 23977 2758 23982 2786
rect 24010 2758 27062 2786
rect 27090 2758 27095 2786
rect 0 2730 56 2744
rect 2227 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2369 2758
rect 12227 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12369 2758
rect 22227 2730 22232 2758
rect 22260 2730 22284 2758
rect 22312 2730 22336 2758
rect 22364 2730 22369 2758
rect 32144 2730 32200 2744
rect 0 2702 1526 2730
rect 1554 2702 1559 2730
rect 4186 2702 7126 2730
rect 7154 2702 7159 2730
rect 7345 2702 7350 2730
rect 7378 2702 9758 2730
rect 9786 2702 9791 2730
rect 10089 2702 10094 2730
rect 10122 2702 12166 2730
rect 12194 2702 12199 2730
rect 12441 2702 12446 2730
rect 12474 2702 13230 2730
rect 13258 2702 13263 2730
rect 13426 2702 18214 2730
rect 18242 2702 18247 2730
rect 18489 2702 18494 2730
rect 18522 2702 20006 2730
rect 20034 2702 20039 2730
rect 22414 2702 30142 2730
rect 30170 2702 30175 2730
rect 31313 2702 31318 2730
rect 31346 2702 32200 2730
rect 0 2688 56 2702
rect 4186 2618 4214 2702
rect 13426 2674 13454 2702
rect 22414 2674 22442 2702
rect 32144 2688 32200 2702
rect 5273 2646 5278 2674
rect 5306 2646 7406 2674
rect 7434 2646 7439 2674
rect 7630 2646 10934 2674
rect 10962 2646 10967 2674
rect 11825 2646 11830 2674
rect 11858 2646 13454 2674
rect 15969 2646 15974 2674
rect 16002 2646 16982 2674
rect 17010 2646 17015 2674
rect 17201 2646 17206 2674
rect 17234 2646 22442 2674
rect 22689 2646 22694 2674
rect 22722 2646 27398 2674
rect 27426 2646 27431 2674
rect 905 2590 910 2618
rect 938 2590 4214 2618
rect 4433 2590 4438 2618
rect 4466 2590 7518 2618
rect 7546 2590 7551 2618
rect 7630 2562 7658 2646
rect 9081 2590 9086 2618
rect 9114 2590 10318 2618
rect 10346 2590 10351 2618
rect 11153 2590 11158 2618
rect 11186 2590 13734 2618
rect 13762 2590 13767 2618
rect 14065 2590 14070 2618
rect 14098 2590 19166 2618
rect 19194 2590 19199 2618
rect 19278 2590 24318 2618
rect 24346 2590 24351 2618
rect 24425 2590 24430 2618
rect 24458 2590 25718 2618
rect 25746 2590 25751 2618
rect 27617 2590 27622 2618
rect 27650 2590 30926 2618
rect 30954 2590 30959 2618
rect 19278 2562 19306 2590
rect 1185 2534 1190 2562
rect 1218 2534 4998 2562
rect 5026 2534 5031 2562
rect 6846 2534 7658 2562
rect 7686 2534 12586 2562
rect 12665 2534 12670 2562
rect 12698 2534 13454 2562
rect 13482 2534 13487 2562
rect 15078 2534 16422 2562
rect 16450 2534 16455 2562
rect 17654 2534 19306 2562
rect 21457 2534 21462 2562
rect 21490 2534 22470 2562
rect 22498 2534 22503 2562
rect 23473 2534 23478 2562
rect 23506 2534 27678 2562
rect 27706 2534 27711 2562
rect 30529 2534 30534 2562
rect 30562 2534 31262 2562
rect 31290 2534 31295 2562
rect 0 2506 56 2520
rect 6846 2506 6874 2534
rect 7686 2506 7714 2534
rect 0 2478 4214 2506
rect 6001 2478 6006 2506
rect 6034 2478 6874 2506
rect 7546 2478 7714 2506
rect 12558 2506 12586 2534
rect 15078 2506 15106 2534
rect 17654 2506 17682 2534
rect 32144 2506 32200 2520
rect 12558 2478 15106 2506
rect 16753 2478 16758 2506
rect 16786 2478 17682 2506
rect 20953 2478 20958 2506
rect 20986 2478 21630 2506
rect 21658 2478 21663 2506
rect 21793 2478 21798 2506
rect 21826 2478 22946 2506
rect 24313 2478 24318 2506
rect 24346 2478 25718 2506
rect 25746 2478 25751 2506
rect 25881 2478 25886 2506
rect 25914 2478 26950 2506
rect 26978 2478 26983 2506
rect 31537 2478 31542 2506
rect 31570 2478 32200 2506
rect 0 2464 56 2478
rect 4186 2450 4214 2478
rect 7546 2450 7574 2478
rect 22918 2450 22946 2478
rect 32144 2464 32200 2478
rect 2529 2422 2534 2450
rect 2562 2422 3822 2450
rect 3850 2422 3855 2450
rect 4186 2422 7574 2450
rect 10038 2422 16478 2450
rect 16506 2422 16511 2450
rect 16585 2422 16590 2450
rect 16618 2422 22274 2450
rect 22918 2422 31094 2450
rect 31122 2422 31127 2450
rect 10038 2394 10066 2422
rect 7401 2366 7406 2394
rect 7434 2366 10066 2394
rect 12609 2366 12614 2394
rect 12642 2366 14742 2394
rect 14770 2366 14775 2394
rect 16641 2366 16646 2394
rect 16674 2366 20902 2394
rect 20930 2366 20935 2394
rect 1897 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2039 2366
rect 11897 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12039 2366
rect 21897 2338 21902 2366
rect 21930 2338 21954 2366
rect 21982 2338 22006 2366
rect 22034 2338 22039 2366
rect 22246 2338 22274 2422
rect 22633 2366 22638 2394
rect 22666 2366 24990 2394
rect 25018 2366 25023 2394
rect 25545 2366 25550 2394
rect 25578 2366 28070 2394
rect 28098 2366 28103 2394
rect 7513 2310 7518 2338
rect 7546 2310 10654 2338
rect 10682 2310 10687 2338
rect 20729 2310 20734 2338
rect 20762 2310 21798 2338
rect 21826 2310 21831 2338
rect 22246 2310 26222 2338
rect 26250 2310 26255 2338
rect 26721 2310 26726 2338
rect 26754 2310 30926 2338
rect 30954 2310 30959 2338
rect 0 2282 56 2296
rect 32144 2282 32200 2296
rect 0 2254 5446 2282
rect 5474 2254 5479 2282
rect 6449 2254 6454 2282
rect 6482 2254 9982 2282
rect 10010 2254 10015 2282
rect 10425 2254 10430 2282
rect 10458 2254 12726 2282
rect 12754 2254 12759 2282
rect 14009 2254 14014 2282
rect 14042 2254 25326 2282
rect 25354 2254 25359 2282
rect 31257 2254 31262 2282
rect 31290 2254 32200 2282
rect 0 2240 56 2254
rect 32144 2240 32200 2254
rect 5945 2198 5950 2226
rect 5978 2198 7238 2226
rect 7266 2198 7271 2226
rect 8465 2198 8470 2226
rect 8498 2198 10374 2226
rect 10402 2198 10407 2226
rect 10481 2198 10486 2226
rect 10514 2198 13510 2226
rect 13538 2198 13543 2226
rect 16529 2198 16534 2226
rect 16562 2198 18326 2226
rect 18354 2198 18359 2226
rect 21793 2198 21798 2226
rect 21826 2198 22638 2226
rect 22666 2198 22671 2226
rect 1017 2142 1022 2170
rect 1050 2142 6734 2170
rect 6762 2142 6767 2170
rect 7126 2142 10822 2170
rect 10850 2142 10855 2170
rect 10929 2142 10934 2170
rect 10962 2142 16702 2170
rect 16730 2142 16735 2170
rect 18433 2142 18438 2170
rect 18466 2142 18830 2170
rect 18858 2142 18863 2170
rect 20337 2142 20342 2170
rect 20370 2142 24038 2170
rect 24066 2142 24071 2170
rect 27729 2142 27734 2170
rect 27762 2142 30254 2170
rect 30282 2142 30287 2170
rect 7126 2114 7154 2142
rect 2081 2086 2086 2114
rect 2114 2086 7154 2114
rect 7233 2086 7238 2114
rect 7266 2086 11494 2114
rect 11522 2086 11527 2114
rect 11606 2086 15974 2114
rect 16002 2086 16007 2114
rect 16249 2086 16254 2114
rect 16282 2086 17262 2114
rect 17290 2086 17295 2114
rect 19105 2086 19110 2114
rect 19138 2086 20510 2114
rect 20538 2086 20543 2114
rect 20729 2086 20734 2114
rect 20762 2086 21070 2114
rect 21098 2086 21103 2114
rect 23921 2086 23926 2114
rect 23954 2086 28518 2114
rect 28546 2086 28551 2114
rect 0 2058 56 2072
rect 0 2030 2814 2058
rect 2842 2030 2847 2058
rect 4153 2030 4158 2058
rect 4186 2030 8974 2058
rect 9002 2030 9007 2058
rect 0 2016 56 2030
rect 11606 2002 11634 2086
rect 32144 2058 32200 2072
rect 5721 1974 5726 2002
rect 5754 1974 11634 2002
rect 11662 2030 12474 2058
rect 13449 2030 13454 2058
rect 13482 2030 20790 2058
rect 20818 2030 20823 2058
rect 21681 2030 21686 2058
rect 21714 2030 24206 2058
rect 24234 2030 24239 2058
rect 24313 2030 24318 2058
rect 24346 2030 25438 2058
rect 25466 2030 25471 2058
rect 31425 2030 31430 2058
rect 31458 2030 32200 2058
rect 2227 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2369 1974
rect 11662 1946 11690 2030
rect 12446 2002 12474 2030
rect 32144 2016 32200 2030
rect 12446 1974 20174 2002
rect 20202 1974 20207 2002
rect 24985 1974 24990 2002
rect 25018 1974 27958 2002
rect 27986 1974 27991 2002
rect 12227 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12369 1974
rect 22227 1946 22232 1974
rect 22260 1946 22284 1974
rect 22312 1946 22336 1974
rect 22364 1946 22369 1974
rect 7121 1918 7126 1946
rect 7154 1918 8414 1946
rect 8442 1918 8447 1946
rect 9137 1918 9142 1946
rect 9170 1918 11690 1946
rect 14289 1918 14294 1946
rect 14322 1918 18382 1946
rect 18410 1918 18415 1946
rect 23081 1918 23086 1946
rect 23114 1918 24962 1946
rect 24934 1890 24962 1918
rect 3481 1862 3486 1890
rect 3514 1862 13678 1890
rect 13706 1862 13711 1890
rect 14681 1862 14686 1890
rect 14714 1862 16198 1890
rect 16226 1862 16231 1890
rect 18433 1862 18438 1890
rect 18466 1862 24822 1890
rect 24850 1862 24855 1890
rect 24934 1862 29638 1890
rect 29666 1862 29671 1890
rect 0 1834 56 1848
rect 32144 1834 32200 1848
rect 0 1806 770 1834
rect 3705 1806 3710 1834
rect 3738 1806 12614 1834
rect 12642 1806 12647 1834
rect 12726 1806 14294 1834
rect 14322 1806 14327 1834
rect 15913 1806 15918 1834
rect 15946 1806 24318 1834
rect 24346 1806 24351 1834
rect 27785 1806 27790 1834
rect 27818 1806 30142 1834
rect 30170 1806 30175 1834
rect 30641 1806 30646 1834
rect 30674 1806 32200 1834
rect 0 1792 56 1806
rect 742 1722 770 1806
rect 12726 1778 12754 1806
rect 32144 1792 32200 1806
rect 849 1750 854 1778
rect 882 1750 7126 1778
rect 7154 1750 7159 1778
rect 7905 1750 7910 1778
rect 7938 1750 11102 1778
rect 11130 1750 11135 1778
rect 11209 1750 11214 1778
rect 11242 1750 12754 1778
rect 12889 1750 12894 1778
rect 12922 1750 15526 1778
rect 15554 1750 15559 1778
rect 15946 1750 19166 1778
rect 19194 1750 19199 1778
rect 22297 1750 22302 1778
rect 22330 1750 24710 1778
rect 24738 1750 24743 1778
rect 28233 1750 28238 1778
rect 28266 1750 28574 1778
rect 28602 1750 28607 1778
rect 15946 1722 15974 1750
rect 742 1694 882 1722
rect 7121 1694 7126 1722
rect 7154 1694 10094 1722
rect 854 1666 882 1694
rect 10066 1666 10094 1694
rect 10878 1694 15190 1722
rect 15218 1694 15223 1722
rect 15302 1694 15974 1722
rect 18209 1694 18214 1722
rect 18242 1694 19726 1722
rect 19754 1694 19759 1722
rect 19889 1694 19894 1722
rect 19922 1694 20230 1722
rect 20258 1694 20263 1722
rect 21401 1694 21406 1722
rect 21434 1694 21798 1722
rect 21826 1694 21831 1722
rect 21910 1694 23254 1722
rect 23282 1694 23287 1722
rect 24313 1694 24318 1722
rect 24346 1694 25830 1722
rect 25858 1694 25863 1722
rect 30641 1694 30646 1722
rect 30674 1694 31318 1722
rect 31346 1694 31351 1722
rect 854 1638 6510 1666
rect 6538 1638 6543 1666
rect 10066 1638 10766 1666
rect 10794 1638 10799 1666
rect 0 1610 56 1624
rect 10878 1610 10906 1694
rect 15302 1666 15330 1694
rect 21910 1666 21938 1694
rect 10985 1638 10990 1666
rect 11018 1638 15330 1666
rect 15801 1638 15806 1666
rect 15834 1638 21938 1666
rect 25545 1638 25550 1666
rect 25578 1638 27230 1666
rect 27258 1638 27263 1666
rect 28065 1638 28070 1666
rect 28098 1638 30926 1666
rect 30954 1638 30959 1666
rect 32144 1610 32200 1624
rect 0 1582 1834 1610
rect 7177 1582 7182 1610
rect 7210 1582 10906 1610
rect 13169 1582 13174 1610
rect 13202 1582 13846 1610
rect 13874 1582 13879 1610
rect 14177 1582 14182 1610
rect 14210 1582 15638 1610
rect 15666 1582 15671 1610
rect 15745 1582 15750 1610
rect 15778 1582 16310 1610
rect 16338 1582 16343 1610
rect 16417 1582 16422 1610
rect 16450 1582 18774 1610
rect 18802 1582 18807 1610
rect 25769 1582 25774 1610
rect 25802 1582 27678 1610
rect 27706 1582 27711 1610
rect 31537 1582 31542 1610
rect 31570 1582 32200 1610
rect 0 1568 56 1582
rect 1806 1498 1834 1582
rect 1897 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2039 1582
rect 11897 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12039 1582
rect 21897 1554 21902 1582
rect 21930 1554 21954 1582
rect 21982 1554 22006 1582
rect 22034 1554 22039 1582
rect 32144 1568 32200 1582
rect 3257 1526 3262 1554
rect 3290 1526 4214 1554
rect 12161 1526 12166 1554
rect 12194 1526 12558 1554
rect 12586 1526 12591 1554
rect 15073 1526 15078 1554
rect 15106 1526 18438 1554
rect 18466 1526 18471 1554
rect 4186 1498 4214 1526
rect 1806 1470 2534 1498
rect 2562 1470 2567 1498
rect 4186 1470 13286 1498
rect 13314 1470 13319 1498
rect 13505 1470 13510 1498
rect 13538 1470 20342 1498
rect 20370 1470 20375 1498
rect 20505 1470 20510 1498
rect 20538 1470 25550 1498
rect 25578 1470 25583 1498
rect 6953 1414 6958 1442
rect 6986 1414 9086 1442
rect 9114 1414 9119 1442
rect 10761 1414 10766 1442
rect 10794 1414 13006 1442
rect 13034 1414 13039 1442
rect 14289 1414 14294 1442
rect 14322 1414 16814 1442
rect 16842 1414 16847 1442
rect 16926 1414 18494 1442
rect 18522 1414 18527 1442
rect 21233 1414 21238 1442
rect 21266 1414 26726 1442
rect 26754 1414 26759 1442
rect 0 1386 56 1400
rect 16926 1386 16954 1414
rect 32144 1386 32200 1400
rect 0 1358 350 1386
rect 378 1358 383 1386
rect 2529 1358 2534 1386
rect 2562 1358 7126 1386
rect 7154 1358 7159 1386
rect 7233 1358 7238 1386
rect 7266 1358 12838 1386
rect 12866 1358 12871 1386
rect 13897 1358 13902 1386
rect 13930 1358 15974 1386
rect 16002 1358 16007 1386
rect 16305 1358 16310 1386
rect 16338 1358 16954 1386
rect 18265 1358 18270 1386
rect 18298 1358 18942 1386
rect 18970 1358 18975 1386
rect 19217 1358 19222 1386
rect 19250 1358 25214 1386
rect 25242 1358 25247 1386
rect 25321 1358 25326 1386
rect 25354 1358 30254 1386
rect 30282 1358 30287 1386
rect 31313 1358 31318 1386
rect 31346 1358 32200 1386
rect 0 1344 56 1358
rect 32144 1344 32200 1358
rect 905 1302 910 1330
rect 938 1302 7070 1330
rect 7098 1302 7103 1330
rect 9193 1302 9198 1330
rect 9226 1302 15134 1330
rect 15162 1302 15167 1330
rect 15246 1302 21294 1330
rect 21322 1302 21327 1330
rect 21625 1302 21630 1330
rect 21658 1302 22302 1330
rect 22330 1302 22335 1330
rect 22465 1302 22470 1330
rect 22498 1302 26446 1330
rect 26474 1302 26479 1330
rect 30641 1302 30646 1330
rect 30674 1302 31374 1330
rect 31402 1302 31407 1330
rect 15246 1274 15274 1302
rect 1185 1246 1190 1274
rect 1218 1246 6790 1274
rect 6818 1246 6823 1274
rect 7345 1246 7350 1274
rect 7378 1246 13678 1274
rect 13706 1246 13711 1274
rect 13841 1246 13846 1274
rect 13874 1246 15274 1274
rect 15857 1246 15862 1274
rect 15890 1246 16198 1274
rect 16226 1246 16231 1274
rect 18769 1246 18774 1274
rect 18802 1246 19222 1274
rect 19250 1246 19255 1274
rect 20169 1246 20174 1274
rect 20202 1246 23646 1274
rect 23674 1246 23679 1274
rect 27001 1246 27006 1274
rect 27034 1246 28350 1274
rect 28378 1246 28383 1274
rect 4993 1190 4998 1218
rect 5026 1190 7462 1218
rect 7490 1190 7495 1218
rect 9977 1190 9982 1218
rect 10010 1190 12166 1218
rect 12194 1190 12199 1218
rect 13953 1190 13958 1218
rect 13986 1190 17150 1218
rect 17178 1190 17183 1218
rect 24761 1190 24766 1218
rect 24794 1190 29582 1218
rect 29610 1190 29615 1218
rect 0 1162 56 1176
rect 2227 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2369 1190
rect 12227 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12369 1190
rect 22227 1162 22232 1190
rect 22260 1162 22284 1190
rect 22312 1162 22336 1190
rect 22364 1162 22369 1190
rect 32144 1162 32200 1176
rect 0 1134 1638 1162
rect 1666 1134 1671 1162
rect 4377 1134 4382 1162
rect 4410 1134 10542 1162
rect 10570 1134 10575 1162
rect 10654 1134 12110 1162
rect 12138 1134 12143 1162
rect 13449 1134 13454 1162
rect 13482 1134 14686 1162
rect 14714 1134 14719 1162
rect 19049 1134 19054 1162
rect 19082 1134 21854 1162
rect 23473 1134 23478 1162
rect 23506 1134 25662 1162
rect 25690 1134 25695 1162
rect 26385 1134 26390 1162
rect 26418 1134 28126 1162
rect 28154 1134 28159 1162
rect 29185 1134 29190 1162
rect 29218 1134 30982 1162
rect 31010 1134 31015 1162
rect 31425 1134 31430 1162
rect 31458 1134 32200 1162
rect 0 1120 56 1134
rect 10654 1106 10682 1134
rect 21826 1106 21854 1134
rect 32144 1120 32200 1134
rect 2361 1078 2366 1106
rect 2394 1078 7070 1106
rect 7098 1078 7103 1106
rect 8297 1078 8302 1106
rect 8330 1078 10682 1106
rect 10710 1078 11158 1106
rect 11186 1078 11191 1106
rect 11601 1078 11606 1106
rect 11634 1078 14070 1106
rect 14098 1078 14103 1106
rect 17593 1078 17598 1106
rect 17626 1078 18466 1106
rect 19609 1078 19614 1106
rect 19642 1078 21182 1106
rect 21210 1078 21215 1106
rect 21826 1078 31094 1106
rect 31122 1078 31127 1106
rect 10710 1050 10738 1078
rect 18438 1050 18466 1078
rect 6673 1022 6678 1050
rect 6706 1022 10738 1050
rect 10817 1022 10822 1050
rect 10850 1022 14518 1050
rect 14546 1022 14551 1050
rect 15465 1022 15470 1050
rect 15498 1022 16366 1050
rect 16394 1022 16399 1050
rect 16753 1022 16758 1050
rect 16786 1022 17934 1050
rect 17962 1022 17967 1050
rect 18438 1022 20902 1050
rect 20930 1022 20935 1050
rect 22409 1022 22414 1050
rect 22442 1022 22694 1050
rect 22722 1022 22727 1050
rect 23081 1022 23086 1050
rect 23114 1022 23702 1050
rect 23730 1022 23735 1050
rect 28513 1022 28518 1050
rect 28546 1022 29918 1050
rect 29946 1022 29951 1050
rect 4186 966 8078 994
rect 8106 966 8111 994
rect 8185 966 8190 994
rect 8218 966 9142 994
rect 9170 966 9175 994
rect 10033 966 10038 994
rect 10066 966 13734 994
rect 13762 966 13767 994
rect 17369 966 17374 994
rect 17402 966 18214 994
rect 18242 966 18247 994
rect 19777 966 19782 994
rect 19810 966 20118 994
rect 20146 966 20151 994
rect 20225 966 20230 994
rect 20258 966 22582 994
rect 22610 966 22615 994
rect 23417 966 23422 994
rect 23450 966 24710 994
rect 24738 966 24743 994
rect 0 938 56 952
rect 4186 938 4214 966
rect 32144 938 32200 952
rect 0 910 854 938
rect 882 910 887 938
rect 961 910 966 938
rect 994 910 4214 938
rect 6393 910 6398 938
rect 6426 910 11214 938
rect 11242 910 11247 938
rect 12385 910 12390 938
rect 12418 910 24038 938
rect 24066 910 24071 938
rect 24313 910 24318 938
rect 24346 910 25886 938
rect 25914 910 25919 938
rect 31537 910 31542 938
rect 31570 910 32200 938
rect 0 896 56 910
rect 32144 896 32200 910
rect 798 854 1022 882
rect 1050 854 1055 882
rect 7513 854 7518 882
rect 7546 854 12782 882
rect 12810 854 12815 882
rect 13006 854 16198 882
rect 16226 854 16231 882
rect 16753 854 16758 882
rect 16786 854 17430 882
rect 17458 854 17463 882
rect 18041 854 18046 882
rect 18074 854 18998 882
rect 19026 854 19031 882
rect 19161 854 19166 882
rect 19194 854 20006 882
rect 20034 854 20039 882
rect 21826 854 21966 882
rect 21994 854 21999 882
rect 23641 854 23646 882
rect 23674 854 25214 882
rect 25242 854 25247 882
rect 25489 854 25494 882
rect 25522 854 27902 882
rect 27930 854 27935 882
rect 30641 854 30646 882
rect 30674 854 31346 882
rect 0 714 56 728
rect 798 714 826 854
rect 2585 798 2590 826
rect 2618 798 5838 826
rect 5866 798 5871 826
rect 5950 798 6846 826
rect 6874 798 6879 826
rect 7065 798 7070 826
rect 7098 798 8022 826
rect 8050 798 8055 826
rect 8409 798 8414 826
rect 8442 798 10094 826
rect 10122 798 10127 826
rect 1897 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2039 798
rect 5950 770 5978 798
rect 11897 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12039 798
rect 5049 742 5054 770
rect 5082 742 5978 770
rect 6281 742 6286 770
rect 6314 742 10878 770
rect 10906 742 10911 770
rect 13006 714 13034 854
rect 21826 826 21854 854
rect 18265 798 18270 826
rect 18298 798 18662 826
rect 18690 798 18695 826
rect 20505 798 20510 826
rect 20538 798 21854 826
rect 23193 798 23198 826
rect 23226 798 23590 826
rect 23618 798 23623 826
rect 24985 798 24990 826
rect 25018 798 25382 826
rect 25410 798 25415 826
rect 25545 798 25550 826
rect 25578 798 30142 826
rect 30170 798 30175 826
rect 21897 770 21902 798
rect 21930 770 21954 798
rect 21982 770 22006 798
rect 22034 770 22039 798
rect 14681 742 14686 770
rect 14714 742 21854 770
rect 22073 742 22078 770
rect 22106 742 22974 770
rect 23002 742 23007 770
rect 23865 742 23870 770
rect 23898 742 24374 770
rect 24402 742 24407 770
rect 24537 742 24542 770
rect 24570 742 25270 770
rect 25298 742 25303 770
rect 29521 742 29526 770
rect 29554 742 30590 770
rect 30618 742 30623 770
rect 21826 714 21854 742
rect 31318 714 31346 854
rect 32144 714 32200 728
rect 0 686 826 714
rect 6169 686 6174 714
rect 6202 686 7350 714
rect 7378 686 7383 714
rect 7961 686 7966 714
rect 7994 686 10094 714
rect 10122 686 10127 714
rect 10201 686 10206 714
rect 10234 686 13034 714
rect 14737 686 14742 714
rect 14770 686 17598 714
rect 17626 686 17631 714
rect 18377 686 18382 714
rect 18410 686 18690 714
rect 21826 686 22470 714
rect 22498 686 22503 714
rect 22577 686 22582 714
rect 22610 686 24766 714
rect 24794 686 24799 714
rect 25433 686 25438 714
rect 25466 686 29302 714
rect 29330 686 29335 714
rect 31318 686 32200 714
rect 0 672 56 686
rect 6785 630 6790 658
rect 6818 630 9310 658
rect 9338 630 9343 658
rect 9417 630 9422 658
rect 9450 630 10850 658
rect 11041 630 11046 658
rect 11074 630 11998 658
rect 12026 630 12031 658
rect 13561 630 13566 658
rect 13594 630 15806 658
rect 15834 630 15839 658
rect 17145 630 17150 658
rect 17178 630 17654 658
rect 17682 630 17687 658
rect 17817 630 17822 658
rect 17850 630 18550 658
rect 18578 630 18583 658
rect 10822 602 10850 630
rect 18662 602 18690 686
rect 32144 672 32200 686
rect 20057 630 20062 658
rect 20090 630 20790 658
rect 20818 630 20823 658
rect 20953 630 20958 658
rect 20986 630 22358 658
rect 22386 630 22391 658
rect 22969 630 22974 658
rect 23002 630 23926 658
rect 23954 630 23959 658
rect 2641 574 2646 602
rect 2674 574 10206 602
rect 10234 574 10239 602
rect 10822 574 11326 602
rect 11354 574 11359 602
rect 11657 574 11662 602
rect 11690 574 13034 602
rect 13113 574 13118 602
rect 13146 574 14854 602
rect 14882 574 14887 602
rect 17201 574 17206 602
rect 17234 574 18438 602
rect 18466 574 18471 602
rect 18662 574 24486 602
rect 24514 574 24519 602
rect 24761 574 24766 602
rect 24794 574 30702 602
rect 30730 574 30735 602
rect 13006 546 13034 574
rect 345 518 350 546
rect 378 518 6678 546
rect 6706 518 6711 546
rect 7289 518 7294 546
rect 7322 518 12894 546
rect 12922 518 12927 546
rect 13006 518 13258 546
rect 13337 518 13342 546
rect 13370 518 13790 546
rect 13818 518 13823 546
rect 13902 518 17654 546
rect 17682 518 17687 546
rect 18489 518 18494 546
rect 18522 518 19838 546
rect 19866 518 19871 546
rect 20281 518 20286 546
rect 20314 518 21854 546
rect 21882 518 21887 546
rect 22078 518 22694 546
rect 22722 518 22727 546
rect 24201 518 24206 546
rect 24234 518 26138 546
rect 26217 518 26222 546
rect 26250 518 31094 546
rect 31122 518 31127 546
rect 0 490 56 504
rect 13230 490 13258 518
rect 13902 490 13930 518
rect 22078 490 22106 518
rect 26110 490 26138 518
rect 32144 490 32200 504
rect 0 462 2086 490
rect 2114 462 2119 490
rect 6841 462 6846 490
rect 6874 462 7518 490
rect 7546 462 7551 490
rect 10369 462 10374 490
rect 10402 462 12446 490
rect 12474 462 12479 490
rect 13230 462 13930 490
rect 14009 462 14014 490
rect 14042 462 14406 490
rect 14434 462 14439 490
rect 15633 462 15638 490
rect 15666 462 16674 490
rect 16921 462 16926 490
rect 16954 462 17934 490
rect 17962 462 17967 490
rect 18713 462 18718 490
rect 18746 462 18751 490
rect 18937 462 18942 490
rect 18970 462 20622 490
rect 20650 462 20655 490
rect 21177 462 21182 490
rect 21210 462 22106 490
rect 22134 462 22442 490
rect 22633 462 22638 490
rect 22666 462 25438 490
rect 25466 462 25471 490
rect 26110 462 26782 490
rect 26810 462 26815 490
rect 29465 462 29470 490
rect 29498 462 29918 490
rect 29946 462 29951 490
rect 30585 462 30590 490
rect 30618 462 32200 490
rect 0 448 56 462
rect 5497 406 5502 434
rect 5530 406 7406 434
rect 7434 406 7439 434
rect 9081 406 9086 434
rect 9114 406 10430 434
rect 10458 406 10463 434
rect 12889 406 12894 434
rect 12922 406 15022 434
rect 15050 406 15055 434
rect 2227 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2369 406
rect 12227 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12369 406
rect 16646 378 16674 462
rect 18718 434 18746 462
rect 22134 434 22162 462
rect 17593 406 17598 434
rect 17626 406 18746 434
rect 19441 406 19446 434
rect 19474 406 22162 434
rect 22414 434 22442 462
rect 32144 448 32200 462
rect 22414 406 30086 434
rect 30114 406 30119 434
rect 22227 378 22232 406
rect 22260 378 22284 406
rect 22312 378 22336 406
rect 22364 378 22369 406
rect 4601 350 4606 378
rect 4634 350 6958 378
rect 6986 350 6991 378
rect 7289 350 7294 378
rect 7322 350 10822 378
rect 10850 350 10855 378
rect 13561 350 13566 378
rect 13594 350 16142 378
rect 16170 350 16175 378
rect 16646 350 19502 378
rect 19530 350 19535 378
rect 25209 350 25214 378
rect 25242 350 26670 378
rect 26698 350 26703 378
rect 2361 294 2366 322
rect 2394 294 2926 322
rect 2954 294 2959 322
rect 3033 294 3038 322
rect 3066 294 7182 322
rect 7210 294 7215 322
rect 7457 294 7462 322
rect 7490 294 9534 322
rect 9562 294 9567 322
rect 10089 294 10094 322
rect 10122 294 13846 322
rect 13874 294 13879 322
rect 13953 294 13958 322
rect 13986 294 18382 322
rect 18410 294 18415 322
rect 19385 294 19390 322
rect 19418 294 20398 322
rect 20426 294 20431 322
rect 22297 294 22302 322
rect 22330 294 22750 322
rect 22778 294 22783 322
rect 23982 294 27454 322
rect 27482 294 27487 322
rect 0 266 56 280
rect 23982 266 24010 294
rect 32144 266 32200 280
rect 0 238 2534 266
rect 2562 238 2567 266
rect 2809 238 2814 266
rect 2842 238 7014 266
rect 7042 238 7047 266
rect 12217 238 12222 266
rect 12250 238 15974 266
rect 16193 238 16198 266
rect 16226 238 20174 266
rect 20202 238 20207 266
rect 20342 238 24010 266
rect 24089 238 24094 266
rect 24122 238 25550 266
rect 25578 238 25583 266
rect 29801 238 29806 266
rect 29834 238 32200 266
rect 0 224 56 238
rect 15946 210 15974 238
rect 2137 182 2142 210
rect 2170 182 4606 210
rect 4634 182 4639 210
rect 4713 182 4718 210
rect 4746 182 8778 210
rect 10089 182 10094 210
rect 10122 182 13454 210
rect 13482 182 13487 210
rect 15946 182 20230 210
rect 20258 182 20263 210
rect 8750 154 8778 182
rect 20342 154 20370 238
rect 32144 224 32200 238
rect 21849 182 21854 210
rect 21882 182 23590 210
rect 23618 182 23623 210
rect 24761 182 24766 210
rect 24794 182 26446 210
rect 26474 182 26479 210
rect 1185 126 1190 154
rect 1218 126 8638 154
rect 8666 126 8671 154
rect 8750 126 10430 154
rect 10458 126 10463 154
rect 10705 126 10710 154
rect 10738 126 10743 154
rect 13337 126 13342 154
rect 13370 126 15974 154
rect 18321 126 18326 154
rect 18354 126 20370 154
rect 22521 126 22526 154
rect 22554 126 24374 154
rect 24402 126 24407 154
rect 10710 98 10738 126
rect 15946 98 15974 126
rect 10710 70 13958 98
rect 13986 70 13991 98
rect 15946 70 22414 98
rect 22442 70 22447 98
rect 22745 70 22750 98
rect 22778 70 24430 98
rect 24458 70 24463 98
rect 0 42 56 56
rect 32144 42 32200 56
rect 0 14 350 42
rect 378 14 383 42
rect 31369 14 31374 42
rect 31402 14 32200 42
rect 0 0 56 14
rect 32144 0 32200 14
<< via3 >>
rect 10486 6958 10514 6986
rect 15862 6902 15890 6930
rect 2086 6790 2114 6818
rect 9086 6790 9114 6818
rect 15862 6790 15890 6818
rect 2232 6650 2260 6678
rect 2284 6650 2312 6678
rect 2336 6650 2364 6678
rect 12232 6650 12260 6678
rect 12284 6650 12312 6678
rect 12336 6650 12364 6678
rect 22232 6650 22260 6678
rect 22284 6650 22312 6678
rect 22336 6650 22364 6678
rect 8918 6510 8946 6538
rect 10486 6342 10514 6370
rect 1902 6258 1930 6286
rect 1954 6258 1982 6286
rect 2006 6258 2034 6286
rect 11902 6258 11930 6286
rect 11954 6258 11982 6286
rect 12006 6258 12034 6286
rect 21902 6258 21930 6286
rect 21954 6258 21982 6286
rect 22006 6258 22034 6286
rect 12110 6230 12138 6258
rect 2086 6062 2114 6090
rect 8918 5950 8946 5978
rect 10094 5894 10122 5922
rect 12110 5894 12138 5922
rect 2232 5866 2260 5894
rect 2284 5866 2312 5894
rect 2336 5866 2364 5894
rect 12232 5866 12260 5894
rect 12284 5866 12312 5894
rect 12336 5866 12364 5894
rect 22232 5866 22260 5894
rect 22284 5866 22312 5894
rect 22336 5866 22364 5894
rect 2086 5838 2114 5866
rect 2086 5558 2114 5586
rect 22638 5558 22666 5586
rect 12110 5502 12138 5530
rect 1902 5474 1930 5502
rect 1954 5474 1982 5502
rect 2006 5474 2034 5502
rect 11902 5474 11930 5502
rect 11954 5474 11982 5502
rect 12006 5474 12034 5502
rect 21902 5474 21930 5502
rect 21954 5474 21982 5502
rect 22006 5474 22034 5502
rect 9142 5446 9170 5474
rect 22526 5278 22554 5306
rect 22638 5278 22666 5306
rect 7126 5222 7154 5250
rect 12110 5222 12138 5250
rect 22526 5166 22554 5194
rect 2232 5082 2260 5110
rect 2284 5082 2312 5110
rect 2336 5082 2364 5110
rect 10878 5054 10906 5082
rect 12232 5082 12260 5110
rect 12284 5082 12312 5110
rect 12336 5082 12364 5110
rect 22232 5082 22260 5110
rect 22284 5082 22312 5110
rect 22336 5082 22364 5110
rect 7574 4942 7602 4970
rect 14686 4998 14714 5026
rect 6790 4886 6818 4914
rect 9198 4886 9226 4914
rect 24094 4830 24122 4858
rect 2086 4774 2114 4802
rect 1902 4690 1930 4718
rect 1954 4690 1982 4718
rect 2006 4690 2034 4718
rect 11902 4690 11930 4718
rect 11954 4690 11982 4718
rect 12006 4690 12034 4718
rect 7574 4662 7602 4690
rect 21902 4690 21930 4718
rect 21954 4690 21982 4718
rect 22006 4690 22034 4718
rect 16758 4662 16786 4690
rect 6790 4550 6818 4578
rect 7518 4494 7546 4522
rect 10094 4438 10122 4466
rect 24094 4438 24122 4466
rect 9198 4382 9226 4410
rect 2232 4298 2260 4326
rect 2284 4298 2312 4326
rect 2336 4298 2364 4326
rect 12232 4298 12260 4326
rect 12284 4298 12312 4326
rect 12336 4298 12364 4326
rect 22232 4298 22260 4326
rect 22284 4298 22312 4326
rect 22336 4298 22364 4326
rect 2086 4270 2114 4298
rect 16758 4270 16786 4298
rect 11046 4214 11074 4242
rect 7518 4158 7546 4186
rect 15974 4158 16002 4186
rect 22918 4046 22946 4074
rect 5614 3990 5642 4018
rect 8414 3934 8442 3962
rect 1902 3906 1930 3934
rect 1954 3906 1982 3934
rect 2006 3906 2034 3934
rect 11902 3906 11930 3934
rect 11954 3906 11982 3934
rect 12006 3906 12034 3934
rect 21902 3906 21930 3934
rect 21954 3906 21982 3934
rect 22006 3906 22034 3934
rect 10430 3822 10458 3850
rect 15974 3822 16002 3850
rect 22918 3822 22946 3850
rect 5614 3766 5642 3794
rect 10430 3654 10458 3682
rect 8414 3598 8442 3626
rect 2232 3514 2260 3542
rect 2284 3514 2312 3542
rect 2336 3514 2364 3542
rect 12232 3514 12260 3542
rect 12284 3514 12312 3542
rect 12336 3514 12364 3542
rect 22232 3514 22260 3542
rect 22284 3514 22312 3542
rect 22336 3514 22364 3542
rect 12110 3374 12138 3402
rect 9254 3318 9282 3346
rect 13230 3262 13258 3290
rect 1902 3122 1930 3150
rect 1954 3122 1982 3150
rect 2006 3122 2034 3150
rect 11902 3122 11930 3150
rect 11954 3122 11982 3150
rect 12006 3122 12034 3150
rect 21902 3122 21930 3150
rect 21954 3122 21982 3150
rect 22006 3122 22034 3150
rect 9086 3094 9114 3122
rect 10038 3094 10066 3122
rect 24430 3094 24458 3122
rect 9254 2982 9282 3010
rect 12670 2926 12698 2954
rect 9142 2870 9170 2898
rect 2232 2730 2260 2758
rect 2284 2730 2312 2758
rect 2336 2730 2364 2758
rect 12232 2730 12260 2758
rect 12284 2730 12312 2758
rect 12336 2730 12364 2758
rect 22232 2730 22260 2758
rect 22284 2730 22312 2758
rect 22336 2730 22364 2758
rect 10094 2702 10122 2730
rect 13230 2702 13258 2730
rect 24430 2590 24458 2618
rect 12670 2534 12698 2562
rect 21798 2478 21826 2506
rect 1902 2338 1930 2366
rect 1954 2338 1982 2366
rect 2006 2338 2034 2366
rect 11902 2338 11930 2366
rect 11954 2338 11982 2366
rect 12006 2338 12034 2366
rect 21902 2338 21930 2366
rect 21954 2338 21982 2366
rect 22006 2338 22034 2366
rect 24990 2366 25018 2394
rect 7518 2310 7546 2338
rect 21798 2310 21826 2338
rect 7238 2198 7266 2226
rect 10822 2142 10850 2170
rect 7238 2086 7266 2114
rect 24318 2030 24346 2058
rect 2232 1946 2260 1974
rect 2284 1946 2312 1974
rect 2336 1946 2364 1974
rect 24990 1974 25018 2002
rect 12232 1946 12260 1974
rect 12284 1946 12312 1974
rect 12336 1946 12364 1974
rect 22232 1946 22260 1974
rect 22284 1946 22312 1974
rect 22336 1946 22364 1974
rect 7126 1918 7154 1946
rect 24318 1806 24346 1834
rect 7126 1750 7154 1778
rect 10990 1638 11018 1666
rect 16310 1582 16338 1610
rect 1902 1554 1930 1582
rect 1954 1554 1982 1582
rect 2006 1554 2034 1582
rect 11902 1554 11930 1582
rect 11954 1554 11982 1582
rect 12006 1554 12034 1582
rect 21902 1554 21930 1582
rect 21954 1554 21982 1582
rect 22006 1554 22034 1582
rect 16310 1358 16338 1386
rect 2232 1162 2260 1190
rect 2284 1162 2312 1190
rect 2336 1162 2364 1190
rect 12232 1162 12260 1190
rect 12284 1162 12312 1190
rect 12336 1162 12364 1190
rect 22232 1162 22260 1190
rect 22284 1162 22312 1190
rect 22336 1162 22364 1190
rect 12110 1134 12138 1162
rect 7070 1078 7098 1106
rect 10094 798 10122 826
rect 1902 770 1930 798
rect 1954 770 1982 798
rect 2006 770 2034 798
rect 11902 770 11930 798
rect 11954 770 11982 798
rect 12006 770 12034 798
rect 21902 770 21930 798
rect 21954 770 21982 798
rect 22006 770 22034 798
rect 14686 742 14714 770
rect 350 518 378 546
rect 7518 462 7546 490
rect 2232 378 2260 406
rect 2284 378 2312 406
rect 2336 378 2364 406
rect 12232 378 12260 406
rect 12284 378 12312 406
rect 12336 378 12364 406
rect 22232 378 22260 406
rect 22284 378 22312 406
rect 22336 378 22364 406
rect 4606 350 4634 378
rect 13958 294 13986 322
rect 4606 182 4634 210
rect 10094 182 10122 210
rect 13958 70 13986 98
rect 350 14 378 42
<< metal4 >>
rect 1888 6286 2048 7112
rect 1888 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2048 6286
rect 1888 5502 2048 6258
rect 2086 6818 2114 6823
rect 2086 6090 2114 6790
rect 2086 6057 2114 6062
rect 2218 6678 2378 7112
rect 10486 6986 10514 6991
rect 2218 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2378 6678
rect 2218 5894 2378 6650
rect 9086 6818 9114 6823
rect 8918 6538 8946 6543
rect 8918 5978 8946 6510
rect 8918 5945 8946 5950
rect 2086 5866 2114 5871
rect 2086 5586 2114 5838
rect 2086 5553 2114 5558
rect 2218 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2378 5894
rect 1888 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2048 5502
rect 1888 4718 2048 5474
rect 2218 5110 2378 5866
rect 2218 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2378 5110
rect 1888 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2048 4718
rect 1888 3934 2048 4690
rect 2086 4802 2114 4807
rect 2086 4298 2114 4774
rect 2086 4265 2114 4270
rect 2218 4326 2378 5082
rect 7126 5250 7154 5255
rect 6790 4914 6818 4919
rect 6790 4578 6818 4886
rect 6790 4545 6818 4550
rect 2218 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2378 4326
rect 1888 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2048 3934
rect 1888 3150 2048 3906
rect 1888 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2048 3150
rect 1888 2366 2048 3122
rect 1888 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2048 2366
rect 1888 1582 2048 2338
rect 1888 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2048 1582
rect 1888 798 2048 1554
rect 1888 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2048 798
rect 350 546 378 551
rect 350 42 378 518
rect 350 9 378 14
rect 1888 0 2048 770
rect 2218 3542 2378 4298
rect 5614 4018 5642 4023
rect 5614 3794 5642 3990
rect 5614 3761 5642 3766
rect 2218 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2378 3542
rect 2218 2758 2378 3514
rect 2218 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2378 2758
rect 2218 1974 2378 2730
rect 7126 2129 7154 5222
rect 7574 4970 7602 4975
rect 7574 4690 7602 4942
rect 7574 4657 7602 4662
rect 7518 4522 7546 4527
rect 7518 4186 7546 4494
rect 7518 4153 7546 4158
rect 8414 3962 8442 3967
rect 8414 3626 8442 3934
rect 8414 3593 8442 3598
rect 9086 3122 9114 6790
rect 10486 6370 10514 6958
rect 10486 6337 10514 6342
rect 11888 6286 12048 7112
rect 11888 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12048 6286
rect 12218 6678 12378 7112
rect 15862 6930 15890 6935
rect 15862 6818 15890 6902
rect 15862 6785 15890 6790
rect 12218 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12378 6678
rect 10094 5922 10122 5927
rect 9086 3089 9114 3094
rect 9142 5474 9170 5479
rect 9142 2898 9170 5446
rect 9198 4914 9226 4919
rect 9198 4410 9226 4886
rect 10094 4466 10122 5894
rect 11888 5502 12048 6258
rect 12110 6258 12138 6263
rect 12110 5922 12138 6230
rect 12110 5889 12138 5894
rect 12218 5894 12378 6650
rect 12218 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12378 5894
rect 11888 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12048 5502
rect 10094 4433 10122 4438
rect 10878 5082 10906 5087
rect 9198 4377 9226 4382
rect 10878 4289 10906 5054
rect 11888 4718 12048 5474
rect 12110 5530 12138 5535
rect 12110 5250 12138 5502
rect 12110 5217 12138 5222
rect 11888 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12048 4718
rect 10878 4261 11074 4289
rect 11046 4242 11074 4261
rect 11046 4209 11074 4214
rect 11888 3934 12048 4690
rect 11888 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12048 3934
rect 10430 3850 10458 3855
rect 10430 3682 10458 3822
rect 10430 3649 10458 3654
rect 9254 3346 9282 3351
rect 9254 3010 9282 3318
rect 11888 3150 12048 3906
rect 12218 5110 12378 5866
rect 12218 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12378 5110
rect 12218 4326 12378 5082
rect 21888 6286 22048 7112
rect 21888 6258 21902 6286
rect 21930 6258 21954 6286
rect 21982 6258 22006 6286
rect 22034 6258 22048 6286
rect 21888 5502 22048 6258
rect 21888 5474 21902 5502
rect 21930 5474 21954 5502
rect 21982 5474 22006 5502
rect 22034 5474 22048 5502
rect 12218 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12378 4326
rect 12218 3542 12378 4298
rect 12218 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12378 3542
rect 9254 2977 9282 2982
rect 10038 3122 10066 3127
rect 9142 2865 9170 2870
rect 10038 2759 10066 3094
rect 11888 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12048 3150
rect 10038 2731 10122 2759
rect 10094 2730 10122 2731
rect 10094 2697 10122 2702
rect 11888 2366 12048 3122
rect 7518 2338 7546 2343
rect 2218 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2378 1974
rect 2218 1190 2378 1946
rect 2218 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2378 1190
rect 2218 406 2378 1162
rect 7070 2101 7154 2129
rect 7238 2226 7266 2231
rect 7238 2114 7266 2198
rect 7070 1106 7098 2101
rect 7238 2081 7266 2086
rect 7126 1946 7154 1951
rect 7126 1778 7154 1918
rect 7126 1745 7154 1750
rect 7070 1073 7098 1078
rect 7518 490 7546 2310
rect 11888 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12048 2366
rect 10822 2170 10850 2175
rect 10822 2129 10850 2142
rect 10822 2101 10906 2129
rect 10878 1679 10906 2101
rect 10878 1666 11018 1679
rect 10878 1651 10990 1666
rect 10990 1633 11018 1638
rect 11888 1582 12048 2338
rect 11888 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12048 1582
rect 7518 457 7546 462
rect 10094 826 10122 831
rect 2218 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2378 406
rect 2218 0 2378 378
rect 4606 378 4634 383
rect 4606 210 4634 350
rect 4606 177 4634 182
rect 10094 210 10122 798
rect 10094 177 10122 182
rect 11888 798 12048 1554
rect 12110 3402 12138 3407
rect 12110 1162 12138 3374
rect 12110 1129 12138 1134
rect 12218 2758 12378 3514
rect 14686 5026 14714 5031
rect 13230 3290 13258 3295
rect 12218 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12378 2758
rect 12218 1974 12378 2730
rect 12670 2954 12698 2959
rect 12670 2562 12698 2926
rect 13230 2730 13258 3262
rect 13230 2697 13258 2702
rect 12670 2529 12698 2534
rect 12218 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12378 1974
rect 12218 1190 12378 1946
rect 12218 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12378 1190
rect 11888 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12048 798
rect 11888 0 12048 770
rect 12218 406 12378 1162
rect 14686 770 14714 4998
rect 21888 4718 22048 5474
rect 16758 4690 16786 4695
rect 16758 4298 16786 4662
rect 16758 4265 16786 4270
rect 21888 4690 21902 4718
rect 21930 4690 21954 4718
rect 21982 4690 22006 4718
rect 22034 4690 22048 4718
rect 15974 4186 16002 4191
rect 15974 3850 16002 4158
rect 15974 3817 16002 3822
rect 21888 3934 22048 4690
rect 21888 3906 21902 3934
rect 21930 3906 21954 3934
rect 21982 3906 22006 3934
rect 22034 3906 22048 3934
rect 21888 3150 22048 3906
rect 21888 3122 21902 3150
rect 21930 3122 21954 3150
rect 21982 3122 22006 3150
rect 22034 3122 22048 3150
rect 21798 2506 21826 2511
rect 21798 2338 21826 2478
rect 21798 2305 21826 2310
rect 21888 2366 22048 3122
rect 21888 2338 21902 2366
rect 21930 2338 21954 2366
rect 21982 2338 22006 2366
rect 22034 2338 22048 2366
rect 16310 1610 16338 1615
rect 16310 1386 16338 1582
rect 16310 1353 16338 1358
rect 21888 1582 22048 2338
rect 21888 1554 21902 1582
rect 21930 1554 21954 1582
rect 21982 1554 22006 1582
rect 22034 1554 22048 1582
rect 14686 737 14714 742
rect 21888 798 22048 1554
rect 21888 770 21902 798
rect 21930 770 21954 798
rect 21982 770 22006 798
rect 22034 770 22048 798
rect 12218 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12378 406
rect 12218 0 12378 378
rect 13958 322 13986 327
rect 13958 98 13986 294
rect 13958 65 13986 70
rect 21888 0 22048 770
rect 22218 6678 22378 7112
rect 22218 6650 22232 6678
rect 22260 6650 22284 6678
rect 22312 6650 22336 6678
rect 22364 6650 22378 6678
rect 22218 5894 22378 6650
rect 22218 5866 22232 5894
rect 22260 5866 22284 5894
rect 22312 5866 22336 5894
rect 22364 5866 22378 5894
rect 22218 5110 22378 5866
rect 22638 5586 22666 5591
rect 22526 5306 22554 5311
rect 22526 5194 22554 5278
rect 22638 5306 22666 5558
rect 22638 5273 22666 5278
rect 22526 5161 22554 5166
rect 22218 5082 22232 5110
rect 22260 5082 22284 5110
rect 22312 5082 22336 5110
rect 22364 5082 22378 5110
rect 22218 4326 22378 5082
rect 24094 4858 24122 4863
rect 24094 4466 24122 4830
rect 24094 4433 24122 4438
rect 22218 4298 22232 4326
rect 22260 4298 22284 4326
rect 22312 4298 22336 4326
rect 22364 4298 22378 4326
rect 22218 3542 22378 4298
rect 22918 4074 22946 4079
rect 22918 3850 22946 4046
rect 22918 3817 22946 3822
rect 22218 3514 22232 3542
rect 22260 3514 22284 3542
rect 22312 3514 22336 3542
rect 22364 3514 22378 3542
rect 22218 2758 22378 3514
rect 22218 2730 22232 2758
rect 22260 2730 22284 2758
rect 22312 2730 22336 2758
rect 22364 2730 22378 2758
rect 22218 1974 22378 2730
rect 24430 3122 24458 3127
rect 24430 2618 24458 3094
rect 24430 2585 24458 2590
rect 24990 2394 25018 2399
rect 22218 1946 22232 1974
rect 22260 1946 22284 1974
rect 22312 1946 22336 1974
rect 22364 1946 22378 1974
rect 22218 1190 22378 1946
rect 24318 2058 24346 2063
rect 24318 1834 24346 2030
rect 24990 2002 25018 2366
rect 24990 1969 25018 1974
rect 24318 1801 24346 1806
rect 22218 1162 22232 1190
rect 22260 1162 22284 1190
rect 22312 1162 22336 1190
rect 22364 1162 22378 1190
rect 22218 406 22378 1162
rect 22218 378 22232 406
rect 22260 378 22284 406
rect 22312 378 22336 406
rect 22364 378 22378 406
rect 22218 0 22378 378
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _000_
timestamp 1486834041
transform 1 0 13608 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _001_
timestamp 1486834041
transform 1 0 15568 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _002_
timestamp 1486834041
transform 1 0 19096 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _003_
timestamp 1486834041
transform 1 0 18760 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _004_
timestamp 1486834041
transform 1 0 16128 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _005_
timestamp 1486834041
transform 1 0 20496 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _006_
timestamp 1486834041
transform 1 0 20776 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _007_
timestamp 1486834041
transform 1 0 17248 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _008_
timestamp 1486834041
transform 1 0 18536 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _009_
timestamp 1486834041
transform 1 0 14616 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _010_
timestamp 1486834041
transform 1 0 16408 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _011_
timestamp 1486834041
transform 1 0 20328 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _012_
timestamp 1486834041
transform 1 0 19376 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _013_
timestamp 1486834041
transform 1 0 15568 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _014_
timestamp 1486834041
transform 1 0 11592 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _015_
timestamp 1486834041
transform 1 0 13608 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _016_
timestamp 1486834041
transform 1 0 14672 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _017_
timestamp 1486834041
transform 1 0 20328 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _018_
timestamp 1486834041
transform 1 0 13048 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _019_
timestamp 1486834041
transform 1 0 18816 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _020_
timestamp 1486834041
transform 1 0 19096 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _021_
timestamp 1486834041
transform 1 0 12712 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _022_
timestamp 1486834041
transform 1 0 15288 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _023_
timestamp 1486834041
transform 1 0 12432 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _024_
timestamp 1486834041
transform 1 0 19936 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _025_
timestamp 1486834041
transform 1 0 14168 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _026_
timestamp 1486834041
transform 1 0 16464 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _027_
timestamp 1486834041
transform 1 0 18368 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _028_
timestamp 1486834041
transform 1 0 18368 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _029_
timestamp 1486834041
transform 1 0 16912 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _030_
timestamp 1486834041
transform 1 0 12712 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _031_
timestamp 1486834041
transform 1 0 21672 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _032_
timestamp 1486834041
transform -1 0 23632 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _033_
timestamp 1486834041
transform -1 0 24472 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _034_
timestamp 1486834041
transform -1 0 25984 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _035_
timestamp 1486834041
transform -1 0 7224 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _036_
timestamp 1486834041
transform -1 0 8848 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _037_
timestamp 1486834041
transform -1 0 10304 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _038_
timestamp 1486834041
transform -1 0 11424 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _039_
timestamp 1486834041
transform -1 0 12656 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _040_
timestamp 1486834041
transform -1 0 16576 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _041_
timestamp 1486834041
transform -1 0 17864 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _042_
timestamp 1486834041
transform -1 0 25592 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _043_
timestamp 1486834041
transform -1 0 26488 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _044_
timestamp 1486834041
transform -1 0 27104 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _045_
timestamp 1486834041
transform -1 0 28336 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _046_
timestamp 1486834041
transform -1 0 28840 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _047_
timestamp 1486834041
transform -1 0 27944 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _048_
timestamp 1486834041
transform 1 0 29288 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _049_
timestamp 1486834041
transform 1 0 30520 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _050_
timestamp 1486834041
transform -1 0 29736 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _051_
timestamp 1486834041
transform -1 0 29568 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _052_
timestamp 1486834041
transform 1 0 6944 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _053_
timestamp 1486834041
transform 1 0 5768 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _054_
timestamp 1486834041
transform 1 0 9688 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _055_
timestamp 1486834041
transform 1 0 10248 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _056_
timestamp 1486834041
transform 1 0 11256 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _057_
timestamp 1486834041
transform 1 0 10472 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _058_
timestamp 1486834041
transform 1 0 8904 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _059_
timestamp 1486834041
transform 1 0 12768 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _060_
timestamp 1486834041
transform 1 0 12544 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _061_
timestamp 1486834041
transform 1 0 13608 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _062_
timestamp 1486834041
transform 1 0 13216 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _063_
timestamp 1486834041
transform 1 0 15120 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _064_
timestamp 1486834041
transform 1 0 16688 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _065_
timestamp 1486834041
transform 1 0 13608 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _066_
timestamp 1486834041
transform 1 0 11424 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _067_
timestamp 1486834041
transform 1 0 15904 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _068_
timestamp 1486834041
transform 1 0 16408 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _069_
timestamp 1486834041
transform 1 0 16912 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _070_
timestamp 1486834041
transform 1 0 17472 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _071_
timestamp 1486834041
transform 1 0 18144 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _072_
timestamp 1486834041
transform -1 0 2744 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _073_
timestamp 1486834041
transform -1 0 1344 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _074_
timestamp 1486834041
transform -1 0 1288 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _075_
timestamp 1486834041
transform -1 0 1288 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _076_
timestamp 1486834041
transform 1 0 17864 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _077_
timestamp 1486834041
transform 1 0 19432 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _078_
timestamp 1486834041
transform -1 0 1288 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _079_
timestamp 1486834041
transform 1 0 20720 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _080_
timestamp 1486834041
transform 1 0 20104 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _081_
timestamp 1486834041
transform 1 0 21224 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _082_
timestamp 1486834041
transform 1 0 21448 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _083_
timestamp 1486834041
transform 1 0 22120 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _084_
timestamp 1486834041
transform 1 0 22456 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _085_
timestamp 1486834041
transform 1 0 23352 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _086_
timestamp 1486834041
transform 1 0 24416 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _087_
timestamp 1486834041
transform 1 0 25368 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _088_
timestamp 1486834041
transform 1 0 26712 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _089_
timestamp 1486834041
transform 1 0 27328 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _090_
timestamp 1486834041
transform 1 0 29288 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _091_
timestamp 1486834041
transform 1 0 30408 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _092_
timestamp 1486834041
transform -1 0 12712 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _093_
timestamp 1486834041
transform -1 0 10472 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _094_
timestamp 1486834041
transform 1 0 29568 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _095_
timestamp 1486834041
transform -1 0 11144 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _096_
timestamp 1486834041
transform -1 0 10808 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _097_
timestamp 1486834041
transform -1 0 6832 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _098_
timestamp 1486834041
transform -1 0 4816 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _099_
timestamp 1486834041
transform -1 0 8008 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _100_
timestamp 1486834041
transform -1 0 6384 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _101_
timestamp 1486834041
transform -1 0 4256 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _102_
timestamp 1486834041
transform -1 0 4816 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _103_
timestamp 1486834041
transform -1 0 2744 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1486834041
transform -1 0 21896 0 -1 2744
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2
timestamp 1486834041
transform 1 0 448 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36
timestamp 1486834041
transform 1 0 2352 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70
timestamp 1486834041
transform 1 0 4256 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104
timestamp 1486834041
transform 1 0 6160 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 8064 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_172
timestamp 1486834041
transform 1 0 9968 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_206
timestamp 1486834041
transform 1 0 11872 0 1 392
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_222
timestamp 1486834041
transform 1 0 12768 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_240
timestamp 1486834041
transform 1 0 13776 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_274
timestamp 1486834041
transform 1 0 15680 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_303
timestamp 1486834041
transform 1 0 17304 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_305
timestamp 1486834041
transform 1 0 17416 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_336
timestamp 1486834041
transform 1 0 19152 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_370
timestamp 1486834041
transform 1 0 21056 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_404
timestamp 1486834041
transform 1 0 22960 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_438
timestamp 1486834041
transform 1 0 24864 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_472
timestamp 1486834041
transform 1 0 26768 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_478
timestamp 1486834041
transform 1 0 27104 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_512
timestamp 1486834041
transform 1 0 29008 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_546
timestamp 1486834041
transform 1 0 30912 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_2
timestamp 1486834041
transform 1 0 448 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_6
timestamp 1486834041
transform 1 0 672 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_8
timestamp 1486834041
transform 1 0 784 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_17
timestamp 1486834041
transform 1 0 1288 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_33
timestamp 1486834041
transform 1 0 2184 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_43
timestamp 1486834041
transform 1 0 2744 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_59
timestamp 1486834041
transform 1 0 3640 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_67
timestamp 1486834041
transform 1 0 4088 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_69
timestamp 1486834041
transform 1 0 4200 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_72
timestamp 1486834041
transform 1 0 4368 0 -1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_136
timestamp 1486834041
transform 1 0 7952 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_142
timestamp 1486834041
transform 1 0 8288 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_158
timestamp 1486834041
transform 1 0 9184 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_166
timestamp 1486834041
transform 1 0 9632 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_170
timestamp 1486834041
transform 1 0 9856 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_172
timestamp 1486834041
transform 1 0 9968 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_189
timestamp 1486834041
transform 1 0 10920 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_205
timestamp 1486834041
transform 1 0 11816 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_209
timestamp 1486834041
transform 1 0 12040 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1486834041
transform 1 0 12208 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_221
timestamp 1486834041
transform 1 0 12712 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_282
timestamp 1486834041
transform 1 0 16128 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_284
timestamp 1486834041
transform 1 0 16240 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_349
timestamp 1486834041
transform 1 0 19880 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_416
timestamp 1486834041
transform 1 0 23632 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_478
timestamp 1486834041
transform 1 0 27104 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_486
timestamp 1486834041
transform 1 0 27552 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_492
timestamp 1486834041
transform 1 0 27888 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_508
timestamp 1486834041
transform 1 0 28784 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_512
timestamp 1486834041
transform 1 0 29008 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_530
timestamp 1486834041
transform 1 0 30016 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_2
timestamp 1486834041
transform 1 0 448 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_6
timestamp 1486834041
transform 1 0 672 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_8
timestamp 1486834041
transform 1 0 784 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_17
timestamp 1486834041
transform 1 0 1288 0 1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_33
timestamp 1486834041
transform 1 0 2184 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1486834041
transform 1 0 2408 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1486834041
transform 1 0 5992 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_107
timestamp 1486834041
transform 1 0 6328 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 9912 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_177
timestamp 1486834041
transform 1 0 10248 0 1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_209
timestamp 1486834041
transform 1 0 12040 0 1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_225
timestamp 1486834041
transform 1 0 12936 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_233
timestamp 1486834041
transform 1 0 13384 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_247
timestamp 1486834041
transform 1 0 14168 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_291
timestamp 1486834041
transform 1 0 16632 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_300
timestamp 1486834041
transform 1 0 17136 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_381
timestamp 1486834041
transform 1 0 21672 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_451
timestamp 1486834041
transform 1 0 25592 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_457
timestamp 1486834041
transform 1 0 25928 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_467
timestamp 1486834041
transform 1 0 26488 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_469
timestamp 1486834041
transform 1 0 26600 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_478
timestamp 1486834041
transform 1 0 27104 0 1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_510
timestamp 1486834041
transform 1 0 28896 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_514
timestamp 1486834041
transform 1 0 29120 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_516
timestamp 1486834041
transform 1 0 29232 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_527
timestamp 1486834041
transform 1 0 29848 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_531
timestamp 1486834041
transform 1 0 30072 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1486834041
transform 1 0 448 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1486834041
transform 1 0 4032 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_72
timestamp 1486834041
transform 1 0 4368 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_88
timestamp 1486834041
transform 1 0 5264 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_96
timestamp 1486834041
transform 1 0 5712 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_108
timestamp 1486834041
transform 1 0 6384 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_116
timestamp 1486834041
transform 1 0 6832 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_126
timestamp 1486834041
transform 1 0 7392 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_134
timestamp 1486834041
transform 1 0 7840 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_138
timestamp 1486834041
transform 1 0 8064 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_142
timestamp 1486834041
transform 1 0 8288 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_206
timestamp 1486834041
transform 1 0 11872 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_212
timestamp 1486834041
transform 1 0 12208 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_228
timestamp 1486834041
transform 1 0 13104 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_236
timestamp 1486834041
transform 1 0 13552 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_259
timestamp 1486834041
transform 1 0 14840 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_263
timestamp 1486834041
transform 1 0 15064 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_290
timestamp 1486834041
transform 1 0 16576 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_306
timestamp 1486834041
transform 1 0 17472 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_310
timestamp 1486834041
transform 1 0 17696 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_312
timestamp 1486834041
transform 1 0 17808 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_343
timestamp 1486834041
transform 1 0 19544 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_347
timestamp 1486834041
transform 1 0 19768 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_349
timestamp 1486834041
transform 1 0 19880 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_408
timestamp 1486834041
transform 1 0 23184 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_416
timestamp 1486834041
transform 1 0 23632 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_458
timestamp 1486834041
transform 1 0 25984 0 -1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_500
timestamp 1486834041
transform 1 0 28336 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_509
timestamp 1486834041
transform 1 0 28840 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_525
timestamp 1486834041
transform 1 0 29736 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_529
timestamp 1486834041
transform 1 0 29960 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1486834041
transform 1 0 448 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 2240 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1486834041
transform 1 0 2408 0 1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1486834041
transform 1 0 5992 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_107
timestamp 1486834041
transform 1 0 6328 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_123
timestamp 1486834041
transform 1 0 7224 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_127
timestamp 1486834041
transform 1 0 7448 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_137
timestamp 1486834041
transform 1 0 8008 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_161
timestamp 1486834041
transform 1 0 9352 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_169
timestamp 1486834041
transform 1 0 9800 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_173
timestamp 1486834041
transform 1 0 10024 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_177
timestamp 1486834041
transform 1 0 10248 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_193
timestamp 1486834041
transform 1 0 11144 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_197
timestamp 1486834041
transform 1 0 11368 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_206
timestamp 1486834041
transform 1 0 11872 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_214
timestamp 1486834041
transform 1 0 12320 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_226
timestamp 1486834041
transform 1 0 12992 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_234
timestamp 1486834041
transform 1 0 13440 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_236
timestamp 1486834041
transform 1 0 13552 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_247
timestamp 1486834041
transform 1 0 14168 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_263
timestamp 1486834041
transform 1 0 15064 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_271
timestamp 1486834041
transform 1 0 15512 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_275
timestamp 1486834041
transform 1 0 15736 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_277
timestamp 1486834041
transform 1 0 15848 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_286
timestamp 1486834041
transform 1 0 16352 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_295
timestamp 1486834041
transform 1 0 16856 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_311
timestamp 1486834041
transform 1 0 17752 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_317
timestamp 1486834041
transform 1 0 18088 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_325
timestamp 1486834041
transform 1 0 18536 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_337
timestamp 1486834041
transform 1 0 19208 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_361
timestamp 1486834041
transform 1 0 20552 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_363
timestamp 1486834041
transform 1 0 20664 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_372
timestamp 1486834041
transform 1 0 21168 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_376
timestamp 1486834041
transform 1 0 21392 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_387
timestamp 1486834041
transform 1 0 22008 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_403
timestamp 1486834041
transform 1 0 22904 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_407
timestamp 1486834041
transform 1 0 23128 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_431
timestamp 1486834041
transform 1 0 24472 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_439
timestamp 1486834041
transform 1 0 24920 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_457
timestamp 1486834041
transform 1 0 25928 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_489
timestamp 1486834041
transform 1 0 27720 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_505
timestamp 1486834041
transform 1 0 28616 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_513
timestamp 1486834041
transform 1 0 29064 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_527
timestamp 1486834041
transform 1 0 29848 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_531
timestamp 1486834041
transform 1 0 30072 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_2
timestamp 1486834041
transform 1 0 448 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_6
timestamp 1486834041
transform 1 0 672 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_8
timestamp 1486834041
transform 1 0 784 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_17
timestamp 1486834041
transform 1 0 1288 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_49
timestamp 1486834041
transform 1 0 3080 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_65
timestamp 1486834041
transform 1 0 3976 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_69
timestamp 1486834041
transform 1 0 4200 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_80
timestamp 1486834041
transform 1 0 4816 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_112
timestamp 1486834041
transform 1 0 6608 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_128
timestamp 1486834041
transform 1 0 7504 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_136
timestamp 1486834041
transform 1 0 7952 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_142
timestamp 1486834041
transform 1 0 8288 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_174
timestamp 1486834041
transform 1 0 10080 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_176
timestamp 1486834041
transform 1 0 10192 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_193
timestamp 1486834041
transform 1 0 11144 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_203
timestamp 1486834041
transform 1 0 11704 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_207
timestamp 1486834041
transform 1 0 11928 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_209
timestamp 1486834041
transform 1 0 12040 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_212
timestamp 1486834041
transform 1 0 12208 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_220
timestamp 1486834041
transform 1 0 12656 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_224
timestamp 1486834041
transform 1 0 12880 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_226
timestamp 1486834041
transform 1 0 12992 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_235
timestamp 1486834041
transform 1 0 13496 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_267
timestamp 1486834041
transform 1 0 15288 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_275
timestamp 1486834041
transform 1 0 15736 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_279
timestamp 1486834041
transform 1 0 15960 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_282
timestamp 1486834041
transform 1 0 16128 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_290
timestamp 1486834041
transform 1 0 16576 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_294
timestamp 1486834041
transform 1 0 16800 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_304
timestamp 1486834041
transform 1 0 17360 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_320
timestamp 1486834041
transform 1 0 18256 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_328
timestamp 1486834041
transform 1 0 18704 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_332
timestamp 1486834041
transform 1 0 18928 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_334
timestamp 1486834041
transform 1 0 19040 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_343
timestamp 1486834041
transform 1 0 19544 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_347
timestamp 1486834041
transform 1 0 19768 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_349
timestamp 1486834041
transform 1 0 19880 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_352
timestamp 1486834041
transform 1 0 20048 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_368
timestamp 1486834041
transform 1 0 20944 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_376
timestamp 1486834041
transform 1 0 21392 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_378
timestamp 1486834041
transform 1 0 21504 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_385
timestamp 1486834041
transform 1 0 21896 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_397
timestamp 1486834041
transform 1 0 22568 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_413
timestamp 1486834041
transform 1 0 23464 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_417
timestamp 1486834041
transform 1 0 23688 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_419
timestamp 1486834041
transform 1 0 23800 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_422
timestamp 1486834041
transform 1 0 23968 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_454
timestamp 1486834041
transform 1 0 25760 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_470
timestamp 1486834041
transform 1 0 26656 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_478
timestamp 1486834041
transform 1 0 27104 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_492
timestamp 1486834041
transform 1 0 27888 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_524
timestamp 1486834041
transform 1 0 29680 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_528
timestamp 1486834041
transform 1 0 29904 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_530
timestamp 1486834041
transform 1 0 30016 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1486834041
transform 1 0 448 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 2240 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1486834041
transform 1 0 2408 0 1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1486834041
transform 1 0 5992 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_107
timestamp 1486834041
transform 1 0 6328 0 1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_171
timestamp 1486834041
transform 1 0 9912 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_177
timestamp 1486834041
transform 1 0 10248 0 1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_241
timestamp 1486834041
transform 1 0 13832 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_247
timestamp 1486834041
transform 1 0 14168 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_279
timestamp 1486834041
transform 1 0 15960 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_295
timestamp 1486834041
transform 1 0 16856 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_303
timestamp 1486834041
transform 1 0 17304 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_305
timestamp 1486834041
transform 1 0 17416 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_314
timestamp 1486834041
transform 1 0 17920 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_317
timestamp 1486834041
transform 1 0 18088 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_349
timestamp 1486834041
transform 1 0 19880 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_365
timestamp 1486834041
transform 1 0 20776 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_381
timestamp 1486834041
transform 1 0 21672 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_387
timestamp 1486834041
transform 1 0 22008 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_403
timestamp 1486834041
transform 1 0 22904 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_419
timestamp 1486834041
transform 1 0 23800 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_435
timestamp 1486834041
transform 1 0 24696 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_443
timestamp 1486834041
transform 1 0 25144 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_457
timestamp 1486834041
transform 1 0 25928 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_465
timestamp 1486834041
transform 1 0 26376 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_469
timestamp 1486834041
transform 1 0 26600 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_479
timestamp 1486834041
transform 1 0 27160 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_511
timestamp 1486834041
transform 1 0 28952 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_519
timestamp 1486834041
transform 1 0 29400 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_523
timestamp 1486834041
transform 1 0 29624 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_527
timestamp 1486834041
transform 1 0 29848 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_535
timestamp 1486834041
transform 1 0 30296 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_2
timestamp 1486834041
transform 1 0 448 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_34
timestamp 1486834041
transform 1 0 2240 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_43
timestamp 1486834041
transform 1 0 2744 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_59
timestamp 1486834041
transform 1 0 3640 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_67
timestamp 1486834041
transform 1 0 4088 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_69
timestamp 1486834041
transform 1 0 4200 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_72
timestamp 1486834041
transform 1 0 4368 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_104
timestamp 1486834041
transform 1 0 6160 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_116
timestamp 1486834041
transform 1 0 6832 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_132
timestamp 1486834041
transform 1 0 7728 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_142
timestamp 1486834041
transform 1 0 8288 0 -1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_206
timestamp 1486834041
transform 1 0 11872 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_212
timestamp 1486834041
transform 1 0 12208 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_244
timestamp 1486834041
transform 1 0 14000 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_260
timestamp 1486834041
transform 1 0 14896 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_264
timestamp 1486834041
transform 1 0 15120 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_266
timestamp 1486834041
transform 1 0 15232 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_275
timestamp 1486834041
transform 1 0 15736 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_279
timestamp 1486834041
transform 1 0 15960 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_282
timestamp 1486834041
transform 1 0 16128 0 -1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_346
timestamp 1486834041
transform 1 0 19712 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_352
timestamp 1486834041
transform 1 0 20048 0 -1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_416
timestamp 1486834041
transform 1 0 23632 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_422
timestamp 1486834041
transform 1 0 23968 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_438
timestamp 1486834041
transform 1 0 24864 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_470
timestamp 1486834041
transform 1 0 26656 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_486
timestamp 1486834041
transform 1 0 27552 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_492
timestamp 1486834041
transform 1 0 27888 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_524
timestamp 1486834041
transform 1 0 29680 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_528
timestamp 1486834041
transform 1 0 29904 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_530
timestamp 1486834041
transform 1 0 30016 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1486834041
transform 1 0 448 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 2240 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_37
timestamp 1486834041
transform 1 0 2408 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_69
timestamp 1486834041
transform 1 0 4200 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_71
timestamp 1486834041
transform 1 0 4312 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_80
timestamp 1486834041
transform 1 0 4816 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_96
timestamp 1486834041
transform 1 0 5712 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_107
timestamp 1486834041
transform 1 0 6328 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_139
timestamp 1486834041
transform 1 0 8120 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_155
timestamp 1486834041
transform 1 0 9016 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_163
timestamp 1486834041
transform 1 0 9464 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_177
timestamp 1486834041
transform 1 0 10248 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_187
timestamp 1486834041
transform 1 0 10808 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_219
timestamp 1486834041
transform 1 0 12600 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_229
timestamp 1486834041
transform 1 0 13160 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_247
timestamp 1486834041
transform 1 0 14168 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_255
timestamp 1486834041
transform 1 0 14616 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_264
timestamp 1486834041
transform 1 0 15120 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_296
timestamp 1486834041
transform 1 0 16912 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_304
timestamp 1486834041
transform 1 0 17360 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_313
timestamp 1486834041
transform 1 0 17864 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_317
timestamp 1486834041
transform 1 0 18088 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_326
timestamp 1486834041
transform 1 0 18592 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_358
timestamp 1486834041
transform 1 0 20384 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_368
timestamp 1486834041
transform 1 0 20944 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_384
timestamp 1486834041
transform 1 0 21840 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_387
timestamp 1486834041
transform 1 0 22008 0 1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_451
timestamp 1486834041
transform 1 0 25592 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_457
timestamp 1486834041
transform 1 0 25928 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_489
timestamp 1486834041
transform 1 0 27720 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_505
timestamp 1486834041
transform 1 0 28616 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_513
timestamp 1486834041
transform 1 0 29064 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_527
timestamp 1486834041
transform 1 0 29848 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_531
timestamp 1486834041
transform 1 0 30072 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1486834041
transform 1 0 448 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1486834041
transform 1 0 4032 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_72
timestamp 1486834041
transform 1 0 4368 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_136
timestamp 1486834041
transform 1 0 7952 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_142
timestamp 1486834041
transform 1 0 8288 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_206
timestamp 1486834041
transform 1 0 11872 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_212
timestamp 1486834041
transform 1 0 12208 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_276
timestamp 1486834041
transform 1 0 15792 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_282
timestamp 1486834041
transform 1 0 16128 0 -1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_314
timestamp 1486834041
transform 1 0 17920 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_338
timestamp 1486834041
transform 1 0 19264 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_346
timestamp 1486834041
transform 1 0 19712 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_352
timestamp 1486834041
transform 1 0 20048 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_416
timestamp 1486834041
transform 1 0 23632 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_422
timestamp 1486834041
transform 1 0 23968 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_486
timestamp 1486834041
transform 1 0 27552 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_492
timestamp 1486834041
transform 1 0 27888 0 -1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_524
timestamp 1486834041
transform 1 0 29680 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_532
timestamp 1486834041
transform 1 0 30128 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_536
timestamp 1486834041
transform 1 0 30352 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_2
timestamp 1486834041
transform 1 0 448 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_18
timestamp 1486834041
transform 1 0 1344 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1486834041
transform 1 0 2240 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1486834041
transform 1 0 2408 0 1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1486834041
transform 1 0 5992 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_107
timestamp 1486834041
transform 1 0 6328 0 1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_171
timestamp 1486834041
transform 1 0 9912 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_177
timestamp 1486834041
transform 1 0 10248 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_193
timestamp 1486834041
transform 1 0 11144 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_209
timestamp 1486834041
transform 1 0 12040 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_241
timestamp 1486834041
transform 1 0 13832 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_255
timestamp 1486834041
transform 1 0 14616 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_287
timestamp 1486834041
transform 1 0 16408 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_295
timestamp 1486834041
transform 1 0 16856 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_304
timestamp 1486834041
transform 1 0 17360 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_312
timestamp 1486834041
transform 1 0 17808 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_314
timestamp 1486834041
transform 1 0 17920 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_317
timestamp 1486834041
transform 1 0 18088 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_349
timestamp 1486834041
transform 1 0 19880 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_358
timestamp 1486834041
transform 1 0 20384 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_374
timestamp 1486834041
transform 1 0 21280 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_382
timestamp 1486834041
transform 1 0 21728 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_384
timestamp 1486834041
transform 1 0 21840 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_387
timestamp 1486834041
transform 1 0 22008 0 1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_451
timestamp 1486834041
transform 1 0 25592 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_457
timestamp 1486834041
transform 1 0 25928 0 1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_521
timestamp 1486834041
transform 1 0 29512 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_527
timestamp 1486834041
transform 1 0 29848 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_531
timestamp 1486834041
transform 1 0 30072 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_2
timestamp 1486834041
transform 1 0 448 0 -1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_34
timestamp 1486834041
transform 1 0 2240 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_50
timestamp 1486834041
transform 1 0 3136 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_58
timestamp 1486834041
transform 1 0 3584 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_72
timestamp 1486834041
transform 1 0 4368 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_136
timestamp 1486834041
transform 1 0 7952 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_142
timestamp 1486834041
transform 1 0 8288 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_206
timestamp 1486834041
transform 1 0 11872 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_212
timestamp 1486834041
transform 1 0 12208 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_224
timestamp 1486834041
transform 1 0 12880 0 -1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_256
timestamp 1486834041
transform 1 0 14672 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_272
timestamp 1486834041
transform 1 0 15568 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_282
timestamp 1486834041
transform 1 0 16128 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_286
timestamp 1486834041
transform 1 0 16352 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_296
timestamp 1486834041
transform 1 0 16912 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_312
timestamp 1486834041
transform 1 0 17808 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_320
timestamp 1486834041
transform 1 0 18256 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_330
timestamp 1486834041
transform 1 0 18816 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_346
timestamp 1486834041
transform 1 0 19712 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_352
timestamp 1486834041
transform 1 0 20048 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_416
timestamp 1486834041
transform 1 0 23632 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_422
timestamp 1486834041
transform 1 0 23968 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_486
timestamp 1486834041
transform 1 0 27552 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_492
timestamp 1486834041
transform 1 0 27888 0 -1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_524
timestamp 1486834041
transform 1 0 29680 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_528
timestamp 1486834041
transform 1 0 29904 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_530
timestamp 1486834041
transform 1 0 30016 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1486834041
transform 1 0 448 0 1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1486834041
transform 1 0 2240 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1486834041
transform 1 0 2408 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1486834041
transform 1 0 5992 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_107
timestamp 1486834041
transform 1 0 6328 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_171
timestamp 1486834041
transform 1 0 9912 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_177
timestamp 1486834041
transform 1 0 10248 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_241
timestamp 1486834041
transform 1 0 13832 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_247
timestamp 1486834041
transform 1 0 14168 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_263
timestamp 1486834041
transform 1 0 15064 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_271
timestamp 1486834041
transform 1 0 15512 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_280
timestamp 1486834041
transform 1 0 16016 0 1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_312
timestamp 1486834041
transform 1 0 17808 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_314
timestamp 1486834041
transform 1 0 17920 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_317
timestamp 1486834041
transform 1 0 18088 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_321
timestamp 1486834041
transform 1 0 18312 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_330
timestamp 1486834041
transform 1 0 18816 0 1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_362
timestamp 1486834041
transform 1 0 20608 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_378
timestamp 1486834041
transform 1 0 21504 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_382
timestamp 1486834041
transform 1 0 21728 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_384
timestamp 1486834041
transform 1 0 21840 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_387
timestamp 1486834041
transform 1 0 22008 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_451
timestamp 1486834041
transform 1 0 25592 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_457
timestamp 1486834041
transform 1 0 25928 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_521
timestamp 1486834041
transform 1 0 29512 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_527
timestamp 1486834041
transform 1 0 29848 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_531
timestamp 1486834041
transform 1 0 30072 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1486834041
transform 1 0 448 0 -1 5880
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1486834041
transform 1 0 4032 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_72
timestamp 1486834041
transform 1 0 4368 0 -1 5880
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_136
timestamp 1486834041
transform 1 0 7952 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_142
timestamp 1486834041
transform 1 0 8288 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_158
timestamp 1486834041
transform 1 0 9184 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_166
timestamp 1486834041
transform 1 0 9632 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_178
timestamp 1486834041
transform 1 0 10304 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_186
timestamp 1486834041
transform 1 0 10752 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_198
timestamp 1486834041
transform 1 0 11424 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_206
timestamp 1486834041
transform 1 0 11872 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_220
timestamp 1486834041
transform 1 0 12656 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_229
timestamp 1486834041
transform 1 0 13160 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_245
timestamp 1486834041
transform 1 0 14056 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_253
timestamp 1486834041
transform 1 0 14504 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_263
timestamp 1486834041
transform 1 0 15064 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_279
timestamp 1486834041
transform 1 0 15960 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_290
timestamp 1486834041
transform 1 0 16576 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_322
timestamp 1486834041
transform 1 0 18368 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_338
timestamp 1486834041
transform 1 0 19264 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_348
timestamp 1486834041
transform 1 0 19824 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_352
timestamp 1486834041
transform 1 0 20048 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_368
timestamp 1486834041
transform 1 0 20944 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_376
timestamp 1486834041
transform 1 0 21392 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_380
timestamp 1486834041
transform 1 0 21616 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_389
timestamp 1486834041
transform 1 0 22120 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_405
timestamp 1486834041
transform 1 0 23016 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_413
timestamp 1486834041
transform 1 0 23464 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_417
timestamp 1486834041
transform 1 0 23688 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_419
timestamp 1486834041
transform 1 0 23800 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_422
timestamp 1486834041
transform 1 0 23968 0 -1 5880
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_486
timestamp 1486834041
transform 1 0 27552 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_492
timestamp 1486834041
transform 1 0 27888 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_508
timestamp 1486834041
transform 1 0 28784 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_516
timestamp 1486834041
transform 1 0 29232 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1486834041
transform 1 0 448 0 1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1486834041
transform 1 0 2240 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1486834041
transform 1 0 2408 0 1 5880
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1486834041
transform 1 0 5992 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_107
timestamp 1486834041
transform 1 0 6328 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_123
timestamp 1486834041
transform 1 0 7224 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_139
timestamp 1486834041
transform 1 0 8120 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_143
timestamp 1486834041
transform 1 0 8344 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_152
timestamp 1486834041
transform 1 0 8848 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_168
timestamp 1486834041
transform 1 0 9744 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_172
timestamp 1486834041
transform 1 0 9968 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_174
timestamp 1486834041
transform 1 0 10080 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_177
timestamp 1486834041
transform 1 0 10248 0 1 5880
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_241
timestamp 1486834041
transform 1 0 13832 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_247
timestamp 1486834041
transform 1 0 14168 0 1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_279
timestamp 1486834041
transform 1 0 15960 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_295
timestamp 1486834041
transform 1 0 16856 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_299
timestamp 1486834041
transform 1 0 17080 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_301
timestamp 1486834041
transform 1 0 17192 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_310
timestamp 1486834041
transform 1 0 17696 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_314
timestamp 1486834041
transform 1 0 17920 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_317
timestamp 1486834041
transform 1 0 18088 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_347
timestamp 1486834041
transform 1 0 19768 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_355
timestamp 1486834041
transform 1 0 20216 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_373
timestamp 1486834041
transform 1 0 21224 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_381
timestamp 1486834041
transform 1 0 21672 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_387
timestamp 1486834041
transform 1 0 22008 0 1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_419
timestamp 1486834041
transform 1 0 23800 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_435
timestamp 1486834041
transform 1 0 24696 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_451
timestamp 1486834041
transform 1 0 25592 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_457
timestamp 1486834041
transform 1 0 25928 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_473
timestamp 1486834041
transform 1 0 26824 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_481
timestamp 1486834041
transform 1 0 27272 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_493
timestamp 1486834041
transform 1 0 27944 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_509
timestamp 1486834041
transform 1 0 28840 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_527
timestamp 1486834041
transform 1 0 29848 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_531
timestamp 1486834041
transform 1 0 30072 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_2
timestamp 1486834041
transform 1 0 448 0 -1 6664
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_18
timestamp 1486834041
transform 1 0 1344 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_20
timestamp 1486834041
transform 1 0 1456 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_27
timestamp 1486834041
transform 1 0 1848 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_31
timestamp 1486834041
transform 1 0 2072 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_33
timestamp 1486834041
transform 1 0 2184 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_36
timestamp 1486834041
transform 1 0 2352 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_44
timestamp 1486834041
transform 1 0 2800 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_46
timestamp 1486834041
transform 1 0 2912 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_61
timestamp 1486834041
transform 1 0 3752 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_65
timestamp 1486834041
transform 1 0 3976 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_67
timestamp 1486834041
transform 1 0 4088 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_70
timestamp 1486834041
transform 1 0 4256 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_72
timestamp 1486834041
transform 1 0 4368 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_87
timestamp 1486834041
transform 1 0 5208 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_95
timestamp 1486834041
transform 1 0 5656 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_99
timestamp 1486834041
transform 1 0 5880 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_101
timestamp 1486834041
transform 1 0 5992 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_118
timestamp 1486834041
transform 1 0 6944 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_138
timestamp 1486834041
transform 1 0 8064 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_146
timestamp 1486834041
transform 1 0 8512 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_150
timestamp 1486834041
transform 1 0 8736 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_165
timestamp 1486834041
transform 1 0 9576 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_169
timestamp 1486834041
transform 1 0 9800 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_172
timestamp 1486834041
transform 1 0 9968 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_176
timestamp 1486834041
transform 1 0 10192 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_191
timestamp 1486834041
transform 1 0 11032 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_199
timestamp 1486834041
transform 1 0 11480 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_203
timestamp 1486834041
transform 1 0 11704 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_220
timestamp 1486834041
transform 1 0 12656 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_240
timestamp 1486834041
transform 1 0 13776 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_248
timestamp 1486834041
transform 1 0 14224 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_252
timestamp 1486834041
transform 1 0 14448 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_254
timestamp 1486834041
transform 1 0 14560 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_269
timestamp 1486834041
transform 1 0 15400 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_271
timestamp 1486834041
transform 1 0 15512 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_274
timestamp 1486834041
transform 1 0 15680 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_278
timestamp 1486834041
transform 1 0 15904 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_280
timestamp 1486834041
transform 1 0 16016 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_295
timestamp 1486834041
transform 1 0 16856 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_303
timestamp 1486834041
transform 1 0 17304 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_305
timestamp 1486834041
transform 1 0 17416 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_322
timestamp 1486834041
transform 1 0 18368 0 -1 6664
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_338
timestamp 1486834041
transform 1 0 19264 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_342
timestamp 1486834041
transform 1 0 19488 0 -1 6664
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_358
timestamp 1486834041
transform 1 0 20384 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_373
timestamp 1486834041
transform 1 0 21224 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_376
timestamp 1486834041
transform 1 0 21392 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_384
timestamp 1486834041
transform 1 0 21840 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_399
timestamp 1486834041
transform 1 0 22680 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_407
timestamp 1486834041
transform 1 0 23128 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_410
timestamp 1486834041
transform 1 0 23296 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_425
timestamp 1486834041
transform 1 0 24136 0 -1 6664
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_441
timestamp 1486834041
transform 1 0 25032 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_444
timestamp 1486834041
transform 1 0 25200 0 -1 6664
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_460
timestamp 1486834041
transform 1 0 26096 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_478
timestamp 1486834041
transform 1 0 27104 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_486
timestamp 1486834041
transform 1 0 27552 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_488
timestamp 1486834041
transform 1 0 27664 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_503
timestamp 1486834041
transform 1 0 28504 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_507
timestamp 1486834041
transform 1 0 28728 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_509
timestamp 1486834041
transform 1 0 28840 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_512
timestamp 1486834041
transform 1 0 29008 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_514
timestamp 1486834041
transform 1 0 29120 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_529
timestamp 1486834041
transform 1 0 29960 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_560
timestamp 1486834041
transform 1 0 31696 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform 1 0 30184 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform 1 0 30072 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform 1 0 30968 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform 1 0 30856 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform 1 0 30072 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform 1 0 30968 0 1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform 1 0 30184 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform 1 0 30856 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform 1 0 30856 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform 1 0 30968 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform 1 0 30968 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform 1 0 29232 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform 1 0 30856 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform 1 0 30968 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 30856 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 30184 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform 1 0 30968 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 30072 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform 1 0 30184 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform 1 0 30016 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform 1 0 28952 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform 1 0 29288 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 30016 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform 1 0 30072 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform 1 0 30184 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 30072 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 30968 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 30856 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 30072 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 30968 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform 1 0 30184 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 30856 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform -1 0 3752 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform -1 0 18368 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform -1 0 19768 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform -1 0 21224 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform -1 0 22680 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform -1 0 24136 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform -1 0 25592 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform -1 0 26992 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform -1 0 28504 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform -1 0 29960 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform 1 0 30912 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform -1 0 5208 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform -1 0 6944 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform 1 0 7168 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform 1 0 8792 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform 1 0 10248 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform 1 0 11872 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform 1 0 12880 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform -1 0 15400 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform -1 0 16856 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform 1 0 12880 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform 1 0 14056 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform 1 0 13664 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform 1 0 14280 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform 1 0 14000 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform 1 0 14448 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform 1 0 15064 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform 1 0 14784 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform 1 0 15232 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform 1 0 15848 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform 1 0 15736 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform 1 0 16296 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform -1 0 17304 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform 1 0 17080 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform 1 0 17584 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform 1 0 17192 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform 1 0 17864 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform 1 0 18368 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform 1 0 18088 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform 1 0 18648 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform 1 0 18312 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform 1 0 21616 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform -1 0 21616 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform -1 0 22960 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform -1 0 23184 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform -1 0 22400 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform -1 0 22792 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform 1 0 19488 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform 1 0 18872 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform 1 0 20272 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform 1 0 19656 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform 1 0 20048 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform 1 0 20832 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform -1 0 20832 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform 1 0 20440 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform 1 0 21392 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform -1 0 24080 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform 1 0 25200 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform 1 0 25536 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform 1 0 24752 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform 1 0 25984 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform 1 0 25032 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform 1 0 26320 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform -1 0 23576 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform -1 0 23184 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform -1 0 24864 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform 1 0 23968 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform 1 0 23576 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform -1 0 24024 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform 1 0 24360 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform 1 0 24752 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform 1 0 23968 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output105
timestamp 1486834041
transform -1 0 1848 0 -1 6664
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_16
timestamp 1486834041
transform 1 0 336 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 31864 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_17
timestamp 1486834041
transform 1 0 336 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 31864 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_18
timestamp 1486834041
transform 1 0 336 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 31864 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_19
timestamp 1486834041
transform 1 0 336 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 31864 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_20
timestamp 1486834041
transform 1 0 336 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 31864 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_21
timestamp 1486834041
transform 1 0 336 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 31864 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_22
timestamp 1486834041
transform 1 0 336 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 31864 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_23
timestamp 1486834041
transform 1 0 336 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 31864 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_24
timestamp 1486834041
transform 1 0 336 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 31864 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_25
timestamp 1486834041
transform 1 0 336 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 31864 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_26
timestamp 1486834041
transform 1 0 336 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 31864 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_27
timestamp 1486834041
transform 1 0 336 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 31864 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_28
timestamp 1486834041
transform 1 0 336 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 31864 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_29
timestamp 1486834041
transform 1 0 336 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 31864 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_30
timestamp 1486834041
transform 1 0 336 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 31864 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_31
timestamp 1486834041
transform 1 0 336 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 31864 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_32
timestamp 1486834041
transform 1 0 2240 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_33
timestamp 1486834041
transform 1 0 4144 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34
timestamp 1486834041
transform 1 0 6048 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1486834041
transform 1 0 7952 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1486834041
transform 1 0 9856 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1486834041
transform 1 0 11760 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1486834041
transform 1 0 13664 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_39
timestamp 1486834041
transform 1 0 15568 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_40
timestamp 1486834041
transform 1 0 17472 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_41
timestamp 1486834041
transform 1 0 19376 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_42
timestamp 1486834041
transform 1 0 21280 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_43
timestamp 1486834041
transform 1 0 23184 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_44
timestamp 1486834041
transform 1 0 25088 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_45
timestamp 1486834041
transform 1 0 26992 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_46
timestamp 1486834041
transform 1 0 28896 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_47
timestamp 1486834041
transform 1 0 30800 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_48
timestamp 1486834041
transform 1 0 4256 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_49
timestamp 1486834041
transform 1 0 8176 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_50
timestamp 1486834041
transform 1 0 12096 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_51
timestamp 1486834041
transform 1 0 16016 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_52
timestamp 1486834041
transform 1 0 19936 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_53
timestamp 1486834041
transform 1 0 23856 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_54
timestamp 1486834041
transform 1 0 27776 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_55
timestamp 1486834041
transform 1 0 31640 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_56
timestamp 1486834041
transform 1 0 2296 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_57
timestamp 1486834041
transform 1 0 6216 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_58
timestamp 1486834041
transform 1 0 10136 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_59
timestamp 1486834041
transform 1 0 14056 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_60
timestamp 1486834041
transform 1 0 17976 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_61
timestamp 1486834041
transform 1 0 21896 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_62
timestamp 1486834041
transform 1 0 25816 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_63
timestamp 1486834041
transform 1 0 29736 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_64
timestamp 1486834041
transform 1 0 4256 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_65
timestamp 1486834041
transform 1 0 8176 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_66
timestamp 1486834041
transform 1 0 12096 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_67
timestamp 1486834041
transform 1 0 16016 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_68
timestamp 1486834041
transform 1 0 19936 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_69
timestamp 1486834041
transform 1 0 23856 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_70
timestamp 1486834041
transform 1 0 27776 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_71
timestamp 1486834041
transform 1 0 31640 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_72
timestamp 1486834041
transform 1 0 2296 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_73
timestamp 1486834041
transform 1 0 6216 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_74
timestamp 1486834041
transform 1 0 10136 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_75
timestamp 1486834041
transform 1 0 14056 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_76
timestamp 1486834041
transform 1 0 17976 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_77
timestamp 1486834041
transform 1 0 21896 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_78
timestamp 1486834041
transform 1 0 25816 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_79
timestamp 1486834041
transform 1 0 29736 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_80
timestamp 1486834041
transform 1 0 4256 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_81
timestamp 1486834041
transform 1 0 8176 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_82
timestamp 1486834041
transform 1 0 12096 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_83
timestamp 1486834041
transform 1 0 16016 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_84
timestamp 1486834041
transform 1 0 19936 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_85
timestamp 1486834041
transform 1 0 23856 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_86
timestamp 1486834041
transform 1 0 27776 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_87
timestamp 1486834041
transform 1 0 31640 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_88
timestamp 1486834041
transform 1 0 2296 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_89
timestamp 1486834041
transform 1 0 6216 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_90
timestamp 1486834041
transform 1 0 10136 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_91
timestamp 1486834041
transform 1 0 14056 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_92
timestamp 1486834041
transform 1 0 17976 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_93
timestamp 1486834041
transform 1 0 21896 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_94
timestamp 1486834041
transform 1 0 25816 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_95
timestamp 1486834041
transform 1 0 29736 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_96
timestamp 1486834041
transform 1 0 4256 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_97
timestamp 1486834041
transform 1 0 8176 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_98
timestamp 1486834041
transform 1 0 12096 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_99
timestamp 1486834041
transform 1 0 16016 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_100
timestamp 1486834041
transform 1 0 19936 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_101
timestamp 1486834041
transform 1 0 23856 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_102
timestamp 1486834041
transform 1 0 27776 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_103
timestamp 1486834041
transform 1 0 31640 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_104
timestamp 1486834041
transform 1 0 2296 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_105
timestamp 1486834041
transform 1 0 6216 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_106
timestamp 1486834041
transform 1 0 10136 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_107
timestamp 1486834041
transform 1 0 14056 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_108
timestamp 1486834041
transform 1 0 17976 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_109
timestamp 1486834041
transform 1 0 21896 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_110
timestamp 1486834041
transform 1 0 25816 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_111
timestamp 1486834041
transform 1 0 29736 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_112
timestamp 1486834041
transform 1 0 4256 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_113
timestamp 1486834041
transform 1 0 8176 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_114
timestamp 1486834041
transform 1 0 12096 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_115
timestamp 1486834041
transform 1 0 16016 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_116
timestamp 1486834041
transform 1 0 19936 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_117
timestamp 1486834041
transform 1 0 23856 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_118
timestamp 1486834041
transform 1 0 27776 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_119
timestamp 1486834041
transform 1 0 31640 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_120
timestamp 1486834041
transform 1 0 2296 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_121
timestamp 1486834041
transform 1 0 6216 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_122
timestamp 1486834041
transform 1 0 10136 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_123
timestamp 1486834041
transform 1 0 14056 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_124
timestamp 1486834041
transform 1 0 17976 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_125
timestamp 1486834041
transform 1 0 21896 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_126
timestamp 1486834041
transform 1 0 25816 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_127
timestamp 1486834041
transform 1 0 29736 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_128
timestamp 1486834041
transform 1 0 4256 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_129
timestamp 1486834041
transform 1 0 8176 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_130
timestamp 1486834041
transform 1 0 12096 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_131
timestamp 1486834041
transform 1 0 16016 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_132
timestamp 1486834041
transform 1 0 19936 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_133
timestamp 1486834041
transform 1 0 23856 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_134
timestamp 1486834041
transform 1 0 27776 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_135
timestamp 1486834041
transform 1 0 31640 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_136
timestamp 1486834041
transform 1 0 2296 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_137
timestamp 1486834041
transform 1 0 6216 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_138
timestamp 1486834041
transform 1 0 10136 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_139
timestamp 1486834041
transform 1 0 14056 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_140
timestamp 1486834041
transform 1 0 17976 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_141
timestamp 1486834041
transform 1 0 21896 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_142
timestamp 1486834041
transform 1 0 25816 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_143
timestamp 1486834041
transform 1 0 29736 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_144
timestamp 1486834041
transform 1 0 4256 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_145
timestamp 1486834041
transform 1 0 8176 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_146
timestamp 1486834041
transform 1 0 12096 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_147
timestamp 1486834041
transform 1 0 16016 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_148
timestamp 1486834041
transform 1 0 19936 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_149
timestamp 1486834041
transform 1 0 23856 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_150
timestamp 1486834041
transform 1 0 27776 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_151
timestamp 1486834041
transform 1 0 31640 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_152
timestamp 1486834041
transform 1 0 2296 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_153
timestamp 1486834041
transform 1 0 6216 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_154
timestamp 1486834041
transform 1 0 10136 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_155
timestamp 1486834041
transform 1 0 14056 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_156
timestamp 1486834041
transform 1 0 17976 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_157
timestamp 1486834041
transform 1 0 21896 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1486834041
transform 1 0 25816 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1486834041
transform 1 0 29736 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_160
timestamp 1486834041
transform 1 0 2240 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_161
timestamp 1486834041
transform 1 0 4144 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_162
timestamp 1486834041
transform 1 0 6048 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1486834041
transform 1 0 7952 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1486834041
transform 1 0 9856 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1486834041
transform 1 0 11760 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1486834041
transform 1 0 13664 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_167
timestamp 1486834041
transform 1 0 15568 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_168
timestamp 1486834041
transform 1 0 17472 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_169
timestamp 1486834041
transform 1 0 19376 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_170
timestamp 1486834041
transform 1 0 21280 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_171
timestamp 1486834041
transform 1 0 23184 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_172
timestamp 1486834041
transform 1 0 25088 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_173
timestamp 1486834041
transform 1 0 26992 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_174
timestamp 1486834041
transform 1 0 28896 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_175
timestamp 1486834041
transform 1 0 30800 0 -1 6664
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 0 56 56 0 FreeSans 224 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 2240 56 2296 0 FreeSans 224 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 2464 56 2520 0 FreeSans 224 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 2688 56 2744 0 FreeSans 224 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 2912 56 2968 0 FreeSans 224 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 3136 56 3192 0 FreeSans 224 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 3360 56 3416 0 FreeSans 224 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 3584 56 3640 0 FreeSans 224 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 3808 56 3864 0 FreeSans 224 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 4032 56 4088 0 FreeSans 224 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 4256 56 4312 0 FreeSans 224 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 224 56 280 0 FreeSans 224 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 4480 56 4536 0 FreeSans 224 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 4704 56 4760 0 FreeSans 224 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 4928 56 4984 0 FreeSans 224 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 5152 56 5208 0 FreeSans 224 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 5376 56 5432 0 FreeSans 224 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 5600 56 5656 0 FreeSans 224 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 5824 56 5880 0 FreeSans 224 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 6048 56 6104 0 FreeSans 224 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 6272 56 6328 0 FreeSans 224 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 6496 56 6552 0 FreeSans 224 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 448 56 504 0 FreeSans 224 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 6720 56 6776 0 FreeSans 224 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 6944 56 7000 0 FreeSans 224 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 672 56 728 0 FreeSans 224 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 896 56 952 0 FreeSans 224 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 1120 56 1176 0 FreeSans 224 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 1344 56 1400 0 FreeSans 224 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 1568 56 1624 0 FreeSans 224 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 1792 56 1848 0 FreeSans 224 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 2016 56 2072 0 FreeSans 224 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 32144 0 32200 56 0 FreeSans 224 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 32144 2240 32200 2296 0 FreeSans 224 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 32144 2464 32200 2520 0 FreeSans 224 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 32144 2688 32200 2744 0 FreeSans 224 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 32144 2912 32200 2968 0 FreeSans 224 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 32144 3136 32200 3192 0 FreeSans 224 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 32144 3360 32200 3416 0 FreeSans 224 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 32144 3584 32200 3640 0 FreeSans 224 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 32144 3808 32200 3864 0 FreeSans 224 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 32144 4032 32200 4088 0 FreeSans 224 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 32144 4256 32200 4312 0 FreeSans 224 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 32144 224 32200 280 0 FreeSans 224 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 32144 4480 32200 4536 0 FreeSans 224 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 32144 4704 32200 4760 0 FreeSans 224 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 32144 4928 32200 4984 0 FreeSans 224 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 32144 5152 32200 5208 0 FreeSans 224 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 32144 5376 32200 5432 0 FreeSans 224 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 32144 5600 32200 5656 0 FreeSans 224 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 32144 5824 32200 5880 0 FreeSans 224 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 32144 6048 32200 6104 0 FreeSans 224 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 32144 6272 32200 6328 0 FreeSans 224 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 32144 6496 32200 6552 0 FreeSans 224 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 32144 448 32200 504 0 FreeSans 224 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 32144 6720 32200 6776 0 FreeSans 224 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 32144 6944 32200 7000 0 FreeSans 224 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 32144 672 32200 728 0 FreeSans 224 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 32144 896 32200 952 0 FreeSans 224 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 32144 1120 32200 1176 0 FreeSans 224 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 32144 1344 32200 1400 0 FreeSans 224 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 32144 1568 32200 1624 0 FreeSans 224 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 32144 1792 32200 1848 0 FreeSans 224 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 32144 2016 32200 2072 0 FreeSans 224 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 25648 0 25704 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 27888 0 27944 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 28112 0 28168 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 28336 0 28392 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 28560 0 28616 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 28784 0 28840 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 29008 0 29064 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 29232 0 29288 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 29456 0 29512 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 29680 0 29736 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 29904 0 29960 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 25872 0 25928 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 26096 0 26152 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 26320 0 26376 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 26544 0 26600 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 26768 0 26824 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 26992 0 27048 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 27216 0 27272 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 27440 0 27496 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 27664 0 27720 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 2912 7056 2968 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 17472 7056 17528 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 18928 7056 18984 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 20384 7056 20440 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 21840 7056 21896 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 23296 7056 23352 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 24752 7056 24808 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 26208 7056 26264 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 27664 7056 27720 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 29120 7056 29176 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 30576 7056 30632 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 4368 7056 4424 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 5824 7056 5880 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 7280 7056 7336 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 8736 7056 8792 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 10192 7056 10248 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 11648 7056 11704 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 13104 7056 13160 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 14560 7056 14616 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 16016 7056 16072 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 2128 0 2184 56 0 FreeSans 224 0 0 0 N1END[0]
port 104 nsew signal input
flabel metal2 s 2352 0 2408 56 0 FreeSans 224 0 0 0 N1END[1]
port 105 nsew signal input
flabel metal2 s 2576 0 2632 56 0 FreeSans 224 0 0 0 N1END[2]
port 106 nsew signal input
flabel metal2 s 2800 0 2856 56 0 FreeSans 224 0 0 0 N1END[3]
port 107 nsew signal input
flabel metal2 s 4816 0 4872 56 0 FreeSans 224 0 0 0 N2END[0]
port 108 nsew signal input
flabel metal2 s 5040 0 5096 56 0 FreeSans 224 0 0 0 N2END[1]
port 109 nsew signal input
flabel metal2 s 5264 0 5320 56 0 FreeSans 224 0 0 0 N2END[2]
port 110 nsew signal input
flabel metal2 s 5488 0 5544 56 0 FreeSans 224 0 0 0 N2END[3]
port 111 nsew signal input
flabel metal2 s 5712 0 5768 56 0 FreeSans 224 0 0 0 N2END[4]
port 112 nsew signal input
flabel metal2 s 5936 0 5992 56 0 FreeSans 224 0 0 0 N2END[5]
port 113 nsew signal input
flabel metal2 s 6160 0 6216 56 0 FreeSans 224 0 0 0 N2END[6]
port 114 nsew signal input
flabel metal2 s 6384 0 6440 56 0 FreeSans 224 0 0 0 N2END[7]
port 115 nsew signal input
flabel metal2 s 3024 0 3080 56 0 FreeSans 224 0 0 0 N2MID[0]
port 116 nsew signal input
flabel metal2 s 3248 0 3304 56 0 FreeSans 224 0 0 0 N2MID[1]
port 117 nsew signal input
flabel metal2 s 3472 0 3528 56 0 FreeSans 224 0 0 0 N2MID[2]
port 118 nsew signal input
flabel metal2 s 3696 0 3752 56 0 FreeSans 224 0 0 0 N2MID[3]
port 119 nsew signal input
flabel metal2 s 3920 0 3976 56 0 FreeSans 224 0 0 0 N2MID[4]
port 120 nsew signal input
flabel metal2 s 4144 0 4200 56 0 FreeSans 224 0 0 0 N2MID[5]
port 121 nsew signal input
flabel metal2 s 4368 0 4424 56 0 FreeSans 224 0 0 0 N2MID[6]
port 122 nsew signal input
flabel metal2 s 4592 0 4648 56 0 FreeSans 224 0 0 0 N2MID[7]
port 123 nsew signal input
flabel metal2 s 6608 0 6664 56 0 FreeSans 224 0 0 0 N4END[0]
port 124 nsew signal input
flabel metal2 s 8848 0 8904 56 0 FreeSans 224 0 0 0 N4END[10]
port 125 nsew signal input
flabel metal2 s 9072 0 9128 56 0 FreeSans 224 0 0 0 N4END[11]
port 126 nsew signal input
flabel metal2 s 9296 0 9352 56 0 FreeSans 224 0 0 0 N4END[12]
port 127 nsew signal input
flabel metal2 s 9520 0 9576 56 0 FreeSans 224 0 0 0 N4END[13]
port 128 nsew signal input
flabel metal2 s 9744 0 9800 56 0 FreeSans 224 0 0 0 N4END[14]
port 129 nsew signal input
flabel metal2 s 9968 0 10024 56 0 FreeSans 224 0 0 0 N4END[15]
port 130 nsew signal input
flabel metal2 s 6832 0 6888 56 0 FreeSans 224 0 0 0 N4END[1]
port 131 nsew signal input
flabel metal2 s 7056 0 7112 56 0 FreeSans 224 0 0 0 N4END[2]
port 132 nsew signal input
flabel metal2 s 7280 0 7336 56 0 FreeSans 224 0 0 0 N4END[3]
port 133 nsew signal input
flabel metal2 s 7504 0 7560 56 0 FreeSans 224 0 0 0 N4END[4]
port 134 nsew signal input
flabel metal2 s 7728 0 7784 56 0 FreeSans 224 0 0 0 N4END[5]
port 135 nsew signal input
flabel metal2 s 7952 0 8008 56 0 FreeSans 224 0 0 0 N4END[6]
port 136 nsew signal input
flabel metal2 s 8176 0 8232 56 0 FreeSans 224 0 0 0 N4END[7]
port 137 nsew signal input
flabel metal2 s 8400 0 8456 56 0 FreeSans 224 0 0 0 N4END[8]
port 138 nsew signal input
flabel metal2 s 8624 0 8680 56 0 FreeSans 224 0 0 0 N4END[9]
port 139 nsew signal input
flabel metal2 s 10192 0 10248 56 0 FreeSans 224 0 0 0 NN4END[0]
port 140 nsew signal input
flabel metal2 s 12432 0 12488 56 0 FreeSans 224 0 0 0 NN4END[10]
port 141 nsew signal input
flabel metal2 s 12656 0 12712 56 0 FreeSans 224 0 0 0 NN4END[11]
port 142 nsew signal input
flabel metal2 s 12880 0 12936 56 0 FreeSans 224 0 0 0 NN4END[12]
port 143 nsew signal input
flabel metal2 s 13104 0 13160 56 0 FreeSans 224 0 0 0 NN4END[13]
port 144 nsew signal input
flabel metal2 s 13328 0 13384 56 0 FreeSans 224 0 0 0 NN4END[14]
port 145 nsew signal input
flabel metal2 s 13552 0 13608 56 0 FreeSans 224 0 0 0 NN4END[15]
port 146 nsew signal input
flabel metal2 s 10416 0 10472 56 0 FreeSans 224 0 0 0 NN4END[1]
port 147 nsew signal input
flabel metal2 s 10640 0 10696 56 0 FreeSans 224 0 0 0 NN4END[2]
port 148 nsew signal input
flabel metal2 s 10864 0 10920 56 0 FreeSans 224 0 0 0 NN4END[3]
port 149 nsew signal input
flabel metal2 s 11088 0 11144 56 0 FreeSans 224 0 0 0 NN4END[4]
port 150 nsew signal input
flabel metal2 s 11312 0 11368 56 0 FreeSans 224 0 0 0 NN4END[5]
port 151 nsew signal input
flabel metal2 s 11536 0 11592 56 0 FreeSans 224 0 0 0 NN4END[6]
port 152 nsew signal input
flabel metal2 s 11760 0 11816 56 0 FreeSans 224 0 0 0 NN4END[7]
port 153 nsew signal input
flabel metal2 s 11984 0 12040 56 0 FreeSans 224 0 0 0 NN4END[8]
port 154 nsew signal input
flabel metal2 s 12208 0 12264 56 0 FreeSans 224 0 0 0 NN4END[9]
port 155 nsew signal input
flabel metal2 s 13776 0 13832 56 0 FreeSans 224 0 0 0 S1BEG[0]
port 156 nsew signal output
flabel metal2 s 14000 0 14056 56 0 FreeSans 224 0 0 0 S1BEG[1]
port 157 nsew signal output
flabel metal2 s 14224 0 14280 56 0 FreeSans 224 0 0 0 S1BEG[2]
port 158 nsew signal output
flabel metal2 s 14448 0 14504 56 0 FreeSans 224 0 0 0 S1BEG[3]
port 159 nsew signal output
flabel metal2 s 14672 0 14728 56 0 FreeSans 224 0 0 0 S2BEG[0]
port 160 nsew signal output
flabel metal2 s 14896 0 14952 56 0 FreeSans 224 0 0 0 S2BEG[1]
port 161 nsew signal output
flabel metal2 s 15120 0 15176 56 0 FreeSans 224 0 0 0 S2BEG[2]
port 162 nsew signal output
flabel metal2 s 15344 0 15400 56 0 FreeSans 224 0 0 0 S2BEG[3]
port 163 nsew signal output
flabel metal2 s 15568 0 15624 56 0 FreeSans 224 0 0 0 S2BEG[4]
port 164 nsew signal output
flabel metal2 s 15792 0 15848 56 0 FreeSans 224 0 0 0 S2BEG[5]
port 165 nsew signal output
flabel metal2 s 16016 0 16072 56 0 FreeSans 224 0 0 0 S2BEG[6]
port 166 nsew signal output
flabel metal2 s 16240 0 16296 56 0 FreeSans 224 0 0 0 S2BEG[7]
port 167 nsew signal output
flabel metal2 s 16464 0 16520 56 0 FreeSans 224 0 0 0 S2BEGb[0]
port 168 nsew signal output
flabel metal2 s 16688 0 16744 56 0 FreeSans 224 0 0 0 S2BEGb[1]
port 169 nsew signal output
flabel metal2 s 16912 0 16968 56 0 FreeSans 224 0 0 0 S2BEGb[2]
port 170 nsew signal output
flabel metal2 s 17136 0 17192 56 0 FreeSans 224 0 0 0 S2BEGb[3]
port 171 nsew signal output
flabel metal2 s 17360 0 17416 56 0 FreeSans 224 0 0 0 S2BEGb[4]
port 172 nsew signal output
flabel metal2 s 17584 0 17640 56 0 FreeSans 224 0 0 0 S2BEGb[5]
port 173 nsew signal output
flabel metal2 s 17808 0 17864 56 0 FreeSans 224 0 0 0 S2BEGb[6]
port 174 nsew signal output
flabel metal2 s 18032 0 18088 56 0 FreeSans 224 0 0 0 S2BEGb[7]
port 175 nsew signal output
flabel metal2 s 18256 0 18312 56 0 FreeSans 224 0 0 0 S4BEG[0]
port 176 nsew signal output
flabel metal2 s 20496 0 20552 56 0 FreeSans 224 0 0 0 S4BEG[10]
port 177 nsew signal output
flabel metal2 s 20720 0 20776 56 0 FreeSans 224 0 0 0 S4BEG[11]
port 178 nsew signal output
flabel metal2 s 20944 0 21000 56 0 FreeSans 224 0 0 0 S4BEG[12]
port 179 nsew signal output
flabel metal2 s 21168 0 21224 56 0 FreeSans 224 0 0 0 S4BEG[13]
port 180 nsew signal output
flabel metal2 s 21392 0 21448 56 0 FreeSans 224 0 0 0 S4BEG[14]
port 181 nsew signal output
flabel metal2 s 21616 0 21672 56 0 FreeSans 224 0 0 0 S4BEG[15]
port 182 nsew signal output
flabel metal2 s 18480 0 18536 56 0 FreeSans 224 0 0 0 S4BEG[1]
port 183 nsew signal output
flabel metal2 s 18704 0 18760 56 0 FreeSans 224 0 0 0 S4BEG[2]
port 184 nsew signal output
flabel metal2 s 18928 0 18984 56 0 FreeSans 224 0 0 0 S4BEG[3]
port 185 nsew signal output
flabel metal2 s 19152 0 19208 56 0 FreeSans 224 0 0 0 S4BEG[4]
port 186 nsew signal output
flabel metal2 s 19376 0 19432 56 0 FreeSans 224 0 0 0 S4BEG[5]
port 187 nsew signal output
flabel metal2 s 19600 0 19656 56 0 FreeSans 224 0 0 0 S4BEG[6]
port 188 nsew signal output
flabel metal2 s 19824 0 19880 56 0 FreeSans 224 0 0 0 S4BEG[7]
port 189 nsew signal output
flabel metal2 s 20048 0 20104 56 0 FreeSans 224 0 0 0 S4BEG[8]
port 190 nsew signal output
flabel metal2 s 20272 0 20328 56 0 FreeSans 224 0 0 0 S4BEG[9]
port 191 nsew signal output
flabel metal2 s 21840 0 21896 56 0 FreeSans 224 0 0 0 SS4BEG[0]
port 192 nsew signal output
flabel metal2 s 24080 0 24136 56 0 FreeSans 224 0 0 0 SS4BEG[10]
port 193 nsew signal output
flabel metal2 s 24304 0 24360 56 0 FreeSans 224 0 0 0 SS4BEG[11]
port 194 nsew signal output
flabel metal2 s 24528 0 24584 56 0 FreeSans 224 0 0 0 SS4BEG[12]
port 195 nsew signal output
flabel metal2 s 24752 0 24808 56 0 FreeSans 224 0 0 0 SS4BEG[13]
port 196 nsew signal output
flabel metal2 s 24976 0 25032 56 0 FreeSans 224 0 0 0 SS4BEG[14]
port 197 nsew signal output
flabel metal2 s 25200 0 25256 56 0 FreeSans 224 0 0 0 SS4BEG[15]
port 198 nsew signal output
flabel metal2 s 22064 0 22120 56 0 FreeSans 224 0 0 0 SS4BEG[1]
port 199 nsew signal output
flabel metal2 s 22288 0 22344 56 0 FreeSans 224 0 0 0 SS4BEG[2]
port 200 nsew signal output
flabel metal2 s 22512 0 22568 56 0 FreeSans 224 0 0 0 SS4BEG[3]
port 201 nsew signal output
flabel metal2 s 22736 0 22792 56 0 FreeSans 224 0 0 0 SS4BEG[4]
port 202 nsew signal output
flabel metal2 s 22960 0 23016 56 0 FreeSans 224 0 0 0 SS4BEG[5]
port 203 nsew signal output
flabel metal2 s 23184 0 23240 56 0 FreeSans 224 0 0 0 SS4BEG[6]
port 204 nsew signal output
flabel metal2 s 23408 0 23464 56 0 FreeSans 224 0 0 0 SS4BEG[7]
port 205 nsew signal output
flabel metal2 s 23632 0 23688 56 0 FreeSans 224 0 0 0 SS4BEG[8]
port 206 nsew signal output
flabel metal2 s 23856 0 23912 56 0 FreeSans 224 0 0 0 SS4BEG[9]
port 207 nsew signal output
flabel metal2 s 25424 0 25480 56 0 FreeSans 224 0 0 0 UserCLK
port 208 nsew signal input
flabel metal2 s 1456 7056 1512 7112 0 FreeSans 224 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal4 s 1888 0 2048 7112 0 FreeSans 736 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 1888 0 2048 28 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 1888 7084 2048 7112 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 11888 0 12048 7112 0 FreeSans 736 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 11888 0 12048 28 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 11888 7084 12048 7112 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 21888 0 22048 7112 0 FreeSans 736 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 21888 0 22048 28 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 21888 7084 22048 7112 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 2218 0 2378 7112 0 FreeSans 736 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 2218 0 2378 28 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 2218 7084 2378 7112 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 12218 0 12378 7112 0 FreeSans 736 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 12218 0 12378 28 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 12218 7084 12378 7112 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 22218 0 22378 7112 0 FreeSans 736 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 22218 0 22378 28 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 22218 7084 22378 7112 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
rlabel metal1 16100 6272 16100 6272 0 VDD
rlabel metal1 16100 6664 16100 6664 0 VSS
rlabel metal3 203 28 203 28 0 FrameData[0]
rlabel metal2 14252 5824 14252 5824 0 FrameData[10]
rlabel metal3 15092 2520 15092 2520 0 FrameData[11]
rlabel metal3 791 2716 791 2716 0 FrameData[12]
rlabel metal2 12180 1372 12180 1372 0 FrameData[13]
rlabel metal3 931 3164 931 3164 0 FrameData[14]
rlabel metal2 13692 3920 13692 3920 0 FrameData[15]
rlabel metal2 14756 3962 14756 3962 0 FrameData[16]
rlabel metal3 3647 3836 3647 3836 0 FrameData[17]
rlabel metal2 10612 4172 10612 4172 0 FrameData[18]
rlabel metal3 1071 4284 1071 4284 0 FrameData[19]
rlabel metal3 1295 252 1295 252 0 FrameData[1]
rlabel metal2 14084 3556 14084 3556 0 FrameData[20]
rlabel metal3 931 4732 931 4732 0 FrameData[21]
rlabel metal3 13468 3360 13468 3360 0 FrameData[22]
rlabel metal2 10052 4704 10052 4704 0 FrameData[23]
rlabel metal2 15764 4200 15764 4200 0 FrameData[24]
rlabel metal2 14308 5432 14308 5432 0 FrameData[25]
rlabel metal3 1071 5852 1071 5852 0 FrameData[26]
rlabel metal3 1071 6076 1071 6076 0 FrameData[27]
rlabel metal3 931 6300 931 6300 0 FrameData[28]
rlabel metal3 2121 6524 2121 6524 0 FrameData[29]
rlabel metal3 1071 476 1071 476 0 FrameData[2]
rlabel metal3 427 6748 427 6748 0 FrameData[30]
rlabel metal3 483 6972 483 6972 0 FrameData[31]
rlabel metal3 427 700 427 700 0 FrameData[3]
rlabel metal3 455 924 455 924 0 FrameData[4]
rlabel metal3 847 1148 847 1148 0 FrameData[5]
rlabel metal3 203 1372 203 1372 0 FrameData[6]
rlabel metal3 931 1596 931 1596 0 FrameData[7]
rlabel metal3 399 1820 399 1820 0 FrameData[8]
rlabel metal3 1435 2044 1435 2044 0 FrameData[9]
rlabel metal3 31773 28 31773 28 0 FrameData_O[0]
rlabel metal3 31717 2268 31717 2268 0 FrameData_O[10]
rlabel metal2 31556 2380 31556 2380 0 FrameData_O[11]
rlabel metal2 31332 2660 31332 2660 0 FrameData_O[12]
rlabel metal2 30660 3080 30660 3080 0 FrameData_O[13]
rlabel metal2 31556 3108 31556 3108 0 FrameData_O[14]
rlabel metal2 30772 3584 30772 3584 0 FrameData_O[15]
rlabel metal2 31444 3444 31444 3444 0 FrameData_O[16]
rlabel metal3 31801 3836 31801 3836 0 FrameData_O[17]
rlabel metal2 31556 3948 31556 3948 0 FrameData_O[18]
rlabel metal3 31801 4284 31801 4284 0 FrameData_O[19]
rlabel metal3 30989 252 30989 252 0 FrameData_O[1]
rlabel metal3 31773 4508 31773 4508 0 FrameData_O[20]
rlabel metal3 31801 4732 31801 4732 0 FrameData_O[21]
rlabel metal3 31773 4956 31773 4956 0 FrameData_O[22]
rlabel metal2 30660 5208 30660 5208 0 FrameData_O[23]
rlabel metal3 31857 5404 31857 5404 0 FrameData_O[24]
rlabel metal3 31409 5628 31409 5628 0 FrameData_O[25]
rlabel metal3 31773 5852 31773 5852 0 FrameData_O[26]
rlabel metal2 30604 6216 30604 6216 0 FrameData_O[27]
rlabel metal2 29540 6244 29540 6244 0 FrameData_O[28]
rlabel metal2 31108 6132 31108 6132 0 FrameData_O[29]
rlabel metal3 31381 476 31381 476 0 FrameData_O[2]
rlabel metal2 31164 5852 31164 5852 0 FrameData_O[30]
rlabel metal2 31332 5796 31332 5796 0 FrameData_O[31]
rlabel metal3 31745 700 31745 700 0 FrameData_O[3]
rlabel metal2 31556 812 31556 812 0 FrameData_O[4]
rlabel metal2 31444 1036 31444 1036 0 FrameData_O[5]
rlabel metal3 31745 1372 31745 1372 0 FrameData_O[6]
rlabel metal2 31556 1540 31556 1540 0 FrameData_O[7]
rlabel metal2 30660 1960 30660 1960 0 FrameData_O[8]
rlabel metal2 31444 1876 31444 1876 0 FrameData_O[9]
rlabel metal2 25676 595 25676 595 0 FrameStrobe[0]
rlabel metal2 25508 1064 25508 1064 0 FrameStrobe[10]
rlabel metal2 26404 1204 26404 1204 0 FrameStrobe[11]
rlabel metal2 28364 651 28364 651 0 FrameStrobe[12]
rlabel metal3 28420 1764 28420 1764 0 FrameStrobe[13]
rlabel metal2 28812 861 28812 861 0 FrameStrobe[14]
rlabel metal3 28448 5068 28448 5068 0 FrameStrobe[15]
rlabel metal2 29260 427 29260 427 0 FrameStrobe[16]
rlabel metal2 29484 203 29484 203 0 FrameStrobe[17]
rlabel metal2 29708 651 29708 651 0 FrameStrobe[18]
rlabel metal2 29932 259 29932 259 0 FrameStrobe[19]
rlabel metal2 25900 399 25900 399 0 FrameStrobe[1]
rlabel metal2 26124 343 26124 343 0 FrameStrobe[2]
rlabel metal2 26348 203 26348 203 0 FrameStrobe[3]
rlabel metal2 8764 6132 8764 6132 0 FrameStrobe[4]
rlabel metal2 26796 259 26796 259 0 FrameStrobe[5]
rlabel metal2 27020 595 27020 595 0 FrameStrobe[6]
rlabel metal2 27244 847 27244 847 0 FrameStrobe[7]
rlabel metal2 27468 175 27468 175 0 FrameStrobe[8]
rlabel metal2 27692 819 27692 819 0 FrameStrobe[9]
rlabel metal2 2940 7049 2940 7049 0 FrameStrobe_O[0]
rlabel metal2 17500 7049 17500 7049 0 FrameStrobe_O[10]
rlabel metal2 19180 6356 19180 6356 0 FrameStrobe_O[11]
rlabel metal2 20412 7049 20412 7049 0 FrameStrobe_O[12]
rlabel metal2 21868 7049 21868 7049 0 FrameStrobe_O[13]
rlabel metal2 23324 7049 23324 7049 0 FrameStrobe_O[14]
rlabel metal2 24892 6188 24892 6188 0 FrameStrobe_O[15]
rlabel metal2 26236 7049 26236 7049 0 FrameStrobe_O[16]
rlabel metal2 27692 7049 27692 7049 0 FrameStrobe_O[17]
rlabel metal2 29148 7049 29148 7049 0 FrameStrobe_O[18]
rlabel metal2 30604 6825 30604 6825 0 FrameStrobe_O[19]
rlabel metal2 4396 7049 4396 7049 0 FrameStrobe_O[1]
rlabel metal2 5852 6797 5852 6797 0 FrameStrobe_O[2]
rlabel metal2 7308 7049 7308 7049 0 FrameStrobe_O[3]
rlabel metal2 8764 7049 8764 7049 0 FrameStrobe_O[4]
rlabel metal2 10220 7049 10220 7049 0 FrameStrobe_O[5]
rlabel metal2 11676 6797 11676 6797 0 FrameStrobe_O[6]
rlabel metal2 13132 6825 13132 6825 0 FrameStrobe_O[7]
rlabel metal2 14588 7049 14588 7049 0 FrameStrobe_O[8]
rlabel metal2 16044 7049 16044 7049 0 FrameStrobe_O[9]
rlabel metal2 2156 119 2156 119 0 N1END[0]
rlabel metal2 2380 175 2380 175 0 N1END[1]
rlabel metal2 2604 427 2604 427 0 N1END[2]
rlabel metal2 2828 147 2828 147 0 N1END[3]
rlabel metal2 4844 1715 4844 1715 0 N2END[0]
rlabel metal2 5068 399 5068 399 0 N2END[1]
rlabel metal2 5292 1351 5292 1351 0 N2END[2]
rlabel metal2 5516 231 5516 231 0 N2END[3]
rlabel metal2 5740 1015 5740 1015 0 N2END[4]
rlabel metal2 5964 1127 5964 1127 0 N2END[5]
rlabel metal2 6188 371 6188 371 0 N2END[6]
rlabel metal2 14308 1624 14308 1624 0 N2END[7]
rlabel metal2 3052 175 3052 175 0 N2MID[0]
rlabel metal2 3276 791 3276 791 0 N2MID[1]
rlabel metal2 3500 959 3500 959 0 N2MID[2]
rlabel metal2 3724 931 3724 931 0 N2MID[3]
rlabel metal2 3948 1687 3948 1687 0 N2MID[4]
rlabel metal2 4172 1043 4172 1043 0 N2MID[5]
rlabel metal2 10556 1120 10556 1120 0 N2MID[6]
rlabel metal2 4620 1575 4620 1575 0 N2MID[7]
rlabel metal4 15876 6860 15876 6860 0 N4END[0]
rlabel metal2 14196 2324 14196 2324 0 N4END[10]
rlabel metal3 14420 3528 14420 3528 0 N4END[11]
rlabel metal2 9324 343 9324 343 0 N4END[12]
rlabel metal2 9548 175 9548 175 0 N4END[13]
rlabel metal3 2730 4396 2730 4396 0 N4END[14]
rlabel metal2 2660 3108 2660 3108 0 N4END[15]
rlabel metal2 6860 259 6860 259 0 N4END[1]
rlabel metal2 14028 3948 14028 3948 0 N4END[2]
rlabel metal2 10836 616 10836 616 0 N4END[3]
rlabel metal2 7532 455 7532 455 0 N4END[4]
rlabel metal3 15960 6496 15960 6496 0 N4END[5]
rlabel metal2 10108 504 10108 504 0 N4END[6]
rlabel metal2 8204 511 8204 511 0 N4END[7]
rlabel metal2 13468 2296 13468 2296 0 N4END[8]
rlabel metal2 1204 560 1204 560 0 N4END[9]
rlabel metal2 2660 784 2660 784 0 NN4END[0]
rlabel metal2 12460 259 12460 259 0 NN4END[10]
rlabel metal2 12684 511 12684 511 0 NN4END[11]
rlabel metal2 12908 231 12908 231 0 NN4END[12]
rlabel metal2 13132 259 13132 259 0 NN4END[13]
rlabel metal2 13356 91 13356 91 0 NN4END[14]
rlabel metal2 13580 203 13580 203 0 NN4END[15]
rlabel metal2 10444 91 10444 91 0 NN4END[1]
rlabel metal2 10668 707 10668 707 0 NN4END[2]
rlabel metal2 10892 399 10892 399 0 NN4END[3]
rlabel metal3 9520 1764 9520 1764 0 NN4END[4]
rlabel metal2 11340 315 11340 315 0 NN4END[5]
rlabel metal2 6692 3304 6692 3304 0 NN4END[6]
rlabel metal3 11256 3388 11256 3388 0 NN4END[7]
rlabel metal2 12012 343 12012 343 0 NN4END[8]
rlabel metal2 12236 147 12236 147 0 NN4END[9]
rlabel metal2 13804 287 13804 287 0 S1BEG[0]
rlabel metal2 14028 259 14028 259 0 S1BEG[1]
rlabel metal2 14252 455 14252 455 0 S1BEG[2]
rlabel metal2 14476 651 14476 651 0 S1BEG[3]
rlabel metal2 14700 343 14700 343 0 S2BEG[0]
rlabel metal2 14924 483 14924 483 0 S2BEG[1]
rlabel metal2 15148 343 15148 343 0 S2BEG[2]
rlabel metal2 15372 343 15372 343 0 S2BEG[3]
rlabel metal2 15596 455 15596 455 0 S2BEG[4]
rlabel metal2 15820 259 15820 259 0 S2BEG[5]
rlabel metal2 16044 259 16044 259 0 S2BEG[6]
rlabel metal2 16268 455 16268 455 0 S2BEG[7]
rlabel metal2 16492 343 16492 343 0 S2BEGb[0]
rlabel metal2 16716 231 16716 231 0 S2BEGb[1]
rlabel metal2 16940 259 16940 259 0 S2BEGb[2]
rlabel metal2 17164 343 17164 343 0 S2BEGb[3]
rlabel metal2 17388 511 17388 511 0 S2BEGb[4]
rlabel metal2 17612 231 17612 231 0 S2BEGb[5]
rlabel metal2 17836 343 17836 343 0 S2BEGb[6]
rlabel metal2 18060 455 18060 455 0 S2BEGb[7]
rlabel metal2 18284 427 18284 427 0 S4BEG[0]
rlabel metal3 21910 868 21910 868 0 S4BEG[10]
rlabel metal2 20748 861 20748 861 0 S4BEG[11]
rlabel metal2 20972 343 20972 343 0 S4BEG[12]
rlabel metal3 22092 504 22092 504 0 S4BEG[13]
rlabel metal3 21616 1708 21616 1708 0 S4BEG[14]
rlabel metal2 21644 679 21644 679 0 S4BEG[15]
rlabel metal2 18508 287 18508 287 0 S4BEG[1]
rlabel metal2 18732 203 18732 203 0 S4BEG[2]
rlabel metal2 18956 259 18956 259 0 S4BEG[3]
rlabel metal2 19180 455 19180 455 0 S4BEG[4]
rlabel metal2 19404 175 19404 175 0 S4BEG[5]
rlabel metal2 19628 567 19628 567 0 S4BEG[6]
rlabel metal2 19852 203 19852 203 0 S4BEG[7]
rlabel metal2 20076 343 20076 343 0 S4BEG[8]
rlabel metal2 20300 287 20300 287 0 S4BEG[9]
rlabel metal2 21868 119 21868 119 0 SS4BEG[0]
rlabel metal2 24108 147 24108 147 0 SS4BEG[10]
rlabel metal2 24332 483 24332 483 0 SS4BEG[11]
rlabel metal2 24556 399 24556 399 0 SS4BEG[12]
rlabel metal2 24780 119 24780 119 0 SS4BEG[13]
rlabel metal2 25004 427 25004 427 0 SS4BEG[14]
rlabel metal2 25228 203 25228 203 0 SS4BEG[15]
rlabel metal2 22092 399 22092 399 0 SS4BEG[1]
rlabel metal2 22316 175 22316 175 0 SS4BEG[2]
rlabel metal2 22540 91 22540 91 0 SS4BEG[3]
rlabel metal2 22764 63 22764 63 0 SS4BEG[4]
rlabel metal2 22988 343 22988 343 0 SS4BEG[5]
rlabel metal2 23212 427 23212 427 0 SS4BEG[6]
rlabel metal2 23436 511 23436 511 0 SS4BEG[7]
rlabel metal2 23660 455 23660 455 0 SS4BEG[8]
rlabel metal2 23884 399 23884 399 0 SS4BEG[9]
rlabel metal2 25452 259 25452 259 0 UserCLK
rlabel metal2 1596 6692 1596 6692 0 UserCLKo
rlabel metal2 14028 2044 14028 2044 0 net1
rlabel metal2 31108 3836 31108 3836 0 net10
rlabel metal3 13020 784 13020 784 0 net100
rlabel metal3 29232 1036 29232 1036 0 net101
rlabel metal4 13972 196 13972 196 0 net102
rlabel metal2 10444 3640 10444 3640 0 net103
rlabel metal2 14140 4676 14140 4676 0 net104
rlabel metal3 15092 4200 15092 4200 0 net105
rlabel metal2 19180 4284 19180 4284 0 net11
rlabel metal2 29316 644 29316 644 0 net12
rlabel metal4 24108 4648 24108 4648 0 net13
rlabel metal2 14980 4508 14980 4508 0 net14
rlabel metal2 15652 3794 15652 3794 0 net15
rlabel metal2 16772 5124 16772 5124 0 net16
rlabel metal2 31108 4900 31108 4900 0 net17
rlabel metal3 22092 4620 22092 4620 0 net18
rlabel metal2 16828 6132 16828 6132 0 net19
rlabel metal3 16996 6020 16996 6020 0 net2
rlabel metal2 18732 4984 18732 4984 0 net20
rlabel metal2 18732 5460 18732 5460 0 net21
rlabel metal2 29372 5096 29372 5096 0 net22
rlabel metal3 22148 448 22148 448 0 net23
rlabel metal2 13076 5264 13076 5264 0 net24
rlabel metal3 23604 4816 23604 4816 0 net25
rlabel metal2 25564 1148 25564 1148 0 net26
rlabel metal2 16604 2128 16604 2128 0 net27
rlabel metal3 29512 1652 29512 1652 0 net28
rlabel metal2 26852 4648 26852 4648 0 net29
rlabel metal2 31108 2296 31108 2296 0 net3
rlabel metal3 20454 1148 20454 1148 0 net30
rlabel metal3 22050 6020 22050 6020 0 net31
rlabel metal2 14980 5768 14980 5768 0 net32
rlabel metal2 3668 6412 3668 6412 0 net33
rlabel metal3 22232 1372 22232 1372 0 net34
rlabel metal2 22428 3696 22428 3696 0 net35
rlabel metal3 23996 1428 23996 1428 0 net36
rlabel metal4 25004 2184 25004 2184 0 net37
rlabel metal2 24052 6300 24052 6300 0 net38
rlabel metal3 26544 6020 26544 6020 0 net39
rlabel metal2 23548 4592 23548 4592 0 net4
rlabel metal2 29596 3668 29596 3668 0 net40
rlabel metal2 30828 4732 30828 4732 0 net41
rlabel metal2 29456 1316 29456 1316 0 net42
rlabel metal2 29204 1092 29204 1092 0 net43
rlabel metal2 5124 6692 5124 6692 0 net44
rlabel metal2 6860 6440 6860 6440 0 net45
rlabel metal2 6916 6328 6916 6328 0 net46
rlabel metal2 8540 6300 8540 6300 0 net47
rlabel metal2 9940 6104 9940 6104 0 net48
rlabel metal2 11060 6104 11060 6104 0 net49
rlabel metal2 15932 5180 15932 5180 0 net5
rlabel metal3 12628 5740 12628 5740 0 net50
rlabel metal2 15316 6104 15316 6104 0 net51
rlabel metal3 17136 6468 17136 6468 0 net52
rlabel metal2 12908 560 12908 560 0 net53
rlabel metal2 14140 2772 14140 2772 0 net54
rlabel metal3 11900 980 11900 980 0 net55
rlabel metal2 14364 2100 14364 2100 0 net56
rlabel metal2 14084 840 14084 840 0 net57
rlabel metal3 12684 1036 12684 1036 0 net58
rlabel metal3 12180 1316 12180 1316 0 net59
rlabel metal3 15960 2912 15960 2912 0 net6
rlabel metal3 14000 588 14000 588 0 net60
rlabel metal2 15428 952 15428 952 0 net61
rlabel metal2 13916 1792 13916 1792 0 net62
rlabel metal2 15820 616 15820 616 0 net63
rlabel metal2 15484 1372 15484 1372 0 net64
rlabel metal2 17080 588 17080 588 0 net65
rlabel metal2 13972 1260 13972 1260 0 net66
rlabel metal3 13916 504 13916 504 0 net67
rlabel metal2 17276 1736 17276 1736 0 net68
rlabel metal3 17360 1036 17360 1036 0 net69
rlabel metal3 22120 3668 22120 3668 0 net7
rlabel metal3 17836 588 17836 588 0 net70
rlabel metal2 18172 2128 18172 2128 0 net71
rlabel metal2 18732 2352 18732 2352 0 net72
rlabel metal2 2436 3052 2436 3052 0 net73
rlabel metal2 21756 1596 21756 1596 0 net74
rlabel metal3 21980 2548 21980 2548 0 net75
rlabel metal2 22820 1736 22820 1736 0 net76
rlabel metal3 23408 1036 23408 1036 0 net77
rlabel metal2 24724 2520 24724 2520 0 net78
rlabel metal3 23520 3108 23520 3108 0 net79
rlabel metal2 27692 3528 27692 3528 0 net8
rlabel metal3 7028 4424 7028 4424 0 net80
rlabel metal3 2562 2604 2562 2604 0 net81
rlabel metal2 13524 1848 13524 1848 0 net82
rlabel metal3 18984 1708 18984 1708 0 net83
rlabel metal3 19964 980 19964 980 0 net84
rlabel metal2 14756 1540 14756 1540 0 net85
rlabel metal3 20916 2100 20916 2100 0 net86
rlabel metal2 20496 1372 20496 1372 0 net87
rlabel metal2 21588 952 21588 952 0 net88
rlabel metal2 23996 1680 23996 1680 0 net89
rlabel metal2 20692 3416 20692 3416 0 net9
rlabel metal2 25508 588 25508 588 0 net90
rlabel metal2 16772 2744 16772 2744 0 net91
rlabel metal2 15092 2212 15092 2212 0 net92
rlabel metal3 10668 1120 10668 1120 0 net93
rlabel metal2 14812 4480 14812 4480 0 net94
rlabel metal2 2380 1064 2380 1064 0 net95
rlabel metal2 23492 1960 23492 1960 0 net96
rlabel metal3 24948 1904 24948 1904 0 net97
rlabel metal3 27748 588 27748 588 0 net98
rlabel metal2 24052 952 24052 952 0 net99
<< properties >>
string FIXED_BBOX 0 0 32200 7112
<< end >>
