module GF_SRAM (A_SRAM0,
    A_SRAM1,
    A_SRAM2,
    A_SRAM3,
    A_SRAM4,
    A_SRAM5,
    A_SRAM6,
    A_SRAM7,
    A_SRAM8,
    CEN_SRAM,
    CLK_SRAM,
    CONFIGURED_top,
    D_SRAM0,
    D_SRAM1,
    D_SRAM2,
    D_SRAM3,
    D_SRAM4,
    D_SRAM5,
    D_SRAM6,
    D_SRAM7,
    GWEN_SRAM,
    Q_SRAM0,
    Q_SRAM1,
    Q_SRAM2,
    Q_SRAM3,
    Q_SRAM4,
    Q_SRAM5,
    Q_SRAM6,
    Q_SRAM7,
    Tile_X0Y0_UserCLKo,
    Tile_X0Y1_UserCLK,
    WEN_SRAM0,
    WEN_SRAM1,
    WEN_SRAM2,
    WEN_SRAM3,
    WEN_SRAM4,
    WEN_SRAM5,
    WEN_SRAM6,
    WEN_SRAM7,
    VDD,
    VSS,
    Tile_X0Y0_E1END,
    Tile_X0Y0_E2END,
    Tile_X0Y0_E2MID,
    Tile_X0Y0_E6END,
    Tile_X0Y0_EE4END,
    Tile_X0Y0_FrameData,
    Tile_X0Y0_FrameData_O,
    Tile_X0Y0_FrameStrobe_O,
    Tile_X0Y0_N1BEG,
    Tile_X0Y0_N2BEG,
    Tile_X0Y0_N2BEGb,
    Tile_X0Y0_N4BEG,
    Tile_X0Y0_S1END,
    Tile_X0Y0_S2END,
    Tile_X0Y0_S2MID,
    Tile_X0Y0_S4END,
    Tile_X0Y0_W1BEG,
    Tile_X0Y0_W2BEG,
    Tile_X0Y0_W2BEGb,
    Tile_X0Y0_W6BEG,
    Tile_X0Y0_WW4BEG,
    Tile_X0Y1_E1END,
    Tile_X0Y1_E2END,
    Tile_X0Y1_E2MID,
    Tile_X0Y1_E6END,
    Tile_X0Y1_EE4END,
    Tile_X0Y1_FrameData,
    Tile_X0Y1_FrameData_O,
    Tile_X0Y1_FrameStrobe,
    Tile_X0Y1_N1END,
    Tile_X0Y1_N2END,
    Tile_X0Y1_N2MID,
    Tile_X0Y1_N4END,
    Tile_X0Y1_S1BEG,
    Tile_X0Y1_S2BEG,
    Tile_X0Y1_S2BEGb,
    Tile_X0Y1_S4BEG,
    Tile_X0Y1_W1BEG,
    Tile_X0Y1_W2BEG,
    Tile_X0Y1_W2BEGb,
    Tile_X0Y1_W6BEG,
    Tile_X0Y1_WW4BEG);
 output A_SRAM0;
 output A_SRAM1;
 output A_SRAM2;
 output A_SRAM3;
 output A_SRAM4;
 output A_SRAM5;
 output A_SRAM6;
 output A_SRAM7;
 output A_SRAM8;
 output CEN_SRAM;
 output CLK_SRAM;
 input CONFIGURED_top;
 output D_SRAM0;
 output D_SRAM1;
 output D_SRAM2;
 output D_SRAM3;
 output D_SRAM4;
 output D_SRAM5;
 output D_SRAM6;
 output D_SRAM7;
 output GWEN_SRAM;
 input Q_SRAM0;
 input Q_SRAM1;
 input Q_SRAM2;
 input Q_SRAM3;
 input Q_SRAM4;
 input Q_SRAM5;
 input Q_SRAM6;
 input Q_SRAM7;
 output Tile_X0Y0_UserCLKo;
 input Tile_X0Y1_UserCLK;
 output WEN_SRAM0;
 output WEN_SRAM1;
 output WEN_SRAM2;
 output WEN_SRAM3;
 output WEN_SRAM4;
 output WEN_SRAM5;
 output WEN_SRAM6;
 output WEN_SRAM7;
 inout VDD;
 inout VSS;
 input [3:0] Tile_X0Y0_E1END;
 input [7:0] Tile_X0Y0_E2END;
 input [7:0] Tile_X0Y0_E2MID;
 input [11:0] Tile_X0Y0_E6END;
 input [15:0] Tile_X0Y0_EE4END;
 input [31:0] Tile_X0Y0_FrameData;
 output [31:0] Tile_X0Y0_FrameData_O;
 output [19:0] Tile_X0Y0_FrameStrobe_O;
 output [3:0] Tile_X0Y0_N1BEG;
 output [7:0] Tile_X0Y0_N2BEG;
 output [7:0] Tile_X0Y0_N2BEGb;
 output [15:0] Tile_X0Y0_N4BEG;
 input [3:0] Tile_X0Y0_S1END;
 input [7:0] Tile_X0Y0_S2END;
 input [7:0] Tile_X0Y0_S2MID;
 input [15:0] Tile_X0Y0_S4END;
 output [3:0] Tile_X0Y0_W1BEG;
 output [7:0] Tile_X0Y0_W2BEG;
 output [7:0] Tile_X0Y0_W2BEGb;
 output [11:0] Tile_X0Y0_W6BEG;
 output [15:0] Tile_X0Y0_WW4BEG;
 input [3:0] Tile_X0Y1_E1END;
 input [7:0] Tile_X0Y1_E2END;
 input [7:0] Tile_X0Y1_E2MID;
 input [11:0] Tile_X0Y1_E6END;
 input [15:0] Tile_X0Y1_EE4END;
 input [31:0] Tile_X0Y1_FrameData;
 output [31:0] Tile_X0Y1_FrameData_O;
 input [19:0] Tile_X0Y1_FrameStrobe;
 input [3:0] Tile_X0Y1_N1END;
 input [7:0] Tile_X0Y1_N2END;
 input [7:0] Tile_X0Y1_N2MID;
 input [15:0] Tile_X0Y1_N4END;
 output [3:0] Tile_X0Y1_S1BEG;
 output [7:0] Tile_X0Y1_S2BEG;
 output [7:0] Tile_X0Y1_S2BEGb;
 output [15:0] Tile_X0Y1_S4BEG;
 output [3:0] Tile_X0Y1_W1BEG;
 output [7:0] Tile_X0Y1_W2BEG;
 output [7:0] Tile_X0Y1_W2BEGb;
 output [11:0] Tile_X0Y1_W6BEG;
 output [15:0] Tile_X0Y1_WW4BEG;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG0 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG1 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG2 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG3 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG0 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG1 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG2 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG3 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG4 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG5 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG6 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG7 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb0 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb1 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb2 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb3 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb4 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb5 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb6 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb7 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG0 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG1 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG2 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG3 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG0 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG1 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG2 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG3 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG4 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG5 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG6 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG7 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG0 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG1 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG2 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG3 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG4 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG5 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG6 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG7 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb0 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb1 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb2 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb3 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb4 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb5 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb6 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb7 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG10 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG11 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG2 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG3 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG4 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG5 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG6 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG7 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG8 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG9 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG10 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG11 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG12 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG13 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG14 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG15 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG4 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG5 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG6 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG7 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG8 ;
 wire \Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG9 ;
 wire \Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_10.A ;
 wire \Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_11.A ;
 wire \Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_8.A ;
 wire \Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_9.A ;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG0 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG1 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG2 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG3 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG0 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG1 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG2 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG3 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG4 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG5 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG6 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG7 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG0 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG1 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG2 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG3 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG4 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG5 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG6 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG7 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb0 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb1 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb2 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb3 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb4 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb5 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb6 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb7 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG10 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG11 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG2 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG3 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG4 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG5 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG6 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG7 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG8 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG9 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG10 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG11 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG12 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG13 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG14 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG15 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG4 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG5 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG6 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG7 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG8 ;
 wire \Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG9 ;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire clknet_0_Tile_X0Y1_UserCLK;
 wire clknet_1_0__leaf_Tile_X0Y1_UserCLK;
 wire clknet_1_1__leaf_Tile_X0Y1_UserCLK;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0210_ (.I(Tile_X0Y1_N2MID[6]),
    .ZN(_0139_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0211_ (.I(Tile_X0Y1_N2END[3]),
    .ZN(_0140_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0212_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .ZN(_0141_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0213_ (.I(Tile_X0Y0_S2MID[2]),
    .ZN(_0142_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0214_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q ),
    .ZN(_0143_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0215_ (.I(CONFIGURED_top),
    .ZN(_0144_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0216_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ),
    .ZN(_0145_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0217_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ),
    .ZN(_0146_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0218_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_0147_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0219_ (.I(Tile_X0Y0_E2END[4]),
    .ZN(_0148_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0220_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ),
    .ZN(_0149_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0221_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ),
    .ZN(_0150_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0222_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ),
    .ZN(_0151_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0223_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ),
    .ZN(_0152_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0224_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ),
    .ZN(_0153_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0225_ (.I(Tile_X0Y1_E6END[4]),
    .ZN(_0154_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0226_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ),
    .ZN(_0155_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0227_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .ZN(_0156_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0228_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .ZN(_0157_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0229_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ),
    .ZN(_0158_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0230_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_0159_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0231_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .ZN(_0160_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0232_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .ZN(_0161_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0233_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .ZN(_0162_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0234_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .ZN(_0163_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0235_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .ZN(_0164_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0236_ (.I0(Tile_X0Y0_E2MID[7]),
    .I1(Tile_X0Y0_E2END[7]),
    .I2(Tile_X0Y0_E6END[8]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit10.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit11.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0237_ (.I0(Tile_X0Y1_N2MID[0]),
    .I1(Tile_X0Y1_N2END[0]),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG0 ),
    .I3(Tile_X0Y0_S2MID[0]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q ),
    .Z(_0165_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0238_ (.I0(Tile_X0Y1_E2MID[7]),
    .I1(Tile_X0Y1_E2END[7]),
    .I2(Tile_X0Y1_E6END[7]),
    .I3(_0165_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0239_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb0 ),
    .I1(Tile_X0Y0_S2MID[0]),
    .I2(Tile_X0Y1_N2MID[0]),
    .I3(Tile_X0Y0_S2END[0]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit9.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit8.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0240_ (.I0(Tile_X0Y1_E2MID[3]),
    .I1(Tile_X0Y1_E2MID[6]),
    .I2(Tile_X0Y1_E2END[1]),
    .I3(Tile_X0Y1_E2END[2]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .Z(_0166_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0241_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .A2(Tile_X0Y1_E2MID[0]),
    .ZN(_0167_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0242_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .A2(_0141_),
    .ZN(_0168_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0243_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .A2(_0140_),
    .B(_0167_),
    .ZN(_0169_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0244_ (.A1(Tile_X0Y1_N2END[2]),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .B(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .C(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .ZN(_0170_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0245_ (.A1(_0139_),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .B(_0170_),
    .ZN(_0171_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _0246_ (.A1(_0141_),
    .A2(_0166_),
    .B1(_0168_),
    .B2(_0169_),
    .C(_0171_),
    .ZN(_0172_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0247_ (.I0(Tile_X0Y1_E2END[4]),
    .I1(Tile_X0Y0_S2MID[3]),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .Z(_0173_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _0248_ (.A1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG0 ),
    .A2(_0168_),
    .B1(_0173_),
    .B2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .C(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .ZN(_0174_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0249_ (.A1(_0141_),
    .A2(Tile_X0Y1_E2END[5]),
    .ZN(_0175_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0250_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(_0142_),
    .ZN(_0176_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0251_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .A3(Tile_X0Y1_E2END[3]),
    .ZN(_0177_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0252_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .A2(_0175_),
    .B(_0177_),
    .C(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .ZN(_0178_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0253_ (.A1(_0176_),
    .A2(_0178_),
    .B(_0143_),
    .ZN(_0179_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0254_ (.A1(_0143_),
    .A2(_0172_),
    .B1(_0174_),
    .B2(_0179_),
    .C(_0144_),
    .ZN(net10),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0255_ (.A1(Tile_X0Y0_E6END[1]),
    .A2(_0145_),
    .ZN(_0180_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0256_ (.A1(_0145_),
    .A2(Tile_X0Y0_S1END[1]),
    .ZN(_0181_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0257_ (.A1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ),
    .A3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1 ),
    .ZN(_0182_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0258_ (.A1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_0181_),
    .B(_0182_),
    .C(_0180_),
    .ZN(_0183_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0259_ (.I0(Tile_X0Y0_E1END[1]),
    .I1(Tile_X0Y0_E6END[9]),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .I3(_0183_),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit4.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit5.Q ),
    .Z(_0184_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0260_ (.I0(Tile_X0Y1_N1END[1]),
    .I1(Tile_X0Y1_N4END[1]),
    .I2(_0184_),
    .I3(Tile_X0Y0_S4END[5]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q ),
    .Z(_0185_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0261_ (.A1(Tile_X0Y1_E6END[1]),
    .A2(_0157_),
    .ZN(_0186_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0262_ (.A1(_0157_),
    .A2(_0184_),
    .ZN(_0187_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0263_ (.A1(Tile_X0Y1_N1END[1]),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .A3(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .ZN(_0188_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0264_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_0187_),
    .B(_0188_),
    .C(_0186_),
    .ZN(_0189_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0265_ (.I0(Tile_X0Y1_E1END[1]),
    .I1(_0185_),
    .I2(Tile_X0Y1_E6END[5]),
    .I3(_0189_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0266_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1 ),
    .I1(Tile_X0Y1_N4END[5]),
    .I2(Tile_X0Y0_S1END[1]),
    .I3(Tile_X0Y0_S4END[1]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit2.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit3.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0267_ (.I0(Tile_X0Y0_E1END[1]),
    .I1(Tile_X0Y0_E6END[5]),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .I3(_0183_),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit0.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit1.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0268_ (.A1(Tile_X0Y0_E6END[2]),
    .A2(_0146_),
    .ZN(_0190_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0269_ (.A1(_0146_),
    .A2(Tile_X0Y0_S1END[2]),
    .ZN(_0191_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0270_ (.A1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ),
    .A2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ),
    .A3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2 ),
    .ZN(_0192_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0271_ (.A1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0191_),
    .B(_0192_),
    .C(_0190_),
    .ZN(_0193_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0272_ (.I0(Tile_X0Y0_E1END[2]),
    .I1(Tile_X0Y0_E6END[10]),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .I3(_0193_),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit6.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit7.Q ),
    .Z(_0194_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0273_ (.I0(Tile_X0Y1_N1END[2]),
    .I1(Tile_X0Y1_N4END[2]),
    .I2(_0194_),
    .I3(Tile_X0Y0_S4END[6]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q ),
    .Z(_0195_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0274_ (.A1(Tile_X0Y1_E6END[2]),
    .A2(_0158_),
    .ZN(_0196_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0275_ (.A1(Tile_X0Y1_N1END[2]),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ),
    .A3(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .ZN(_0197_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0276_ (.A1(_0158_),
    .A2(_0194_),
    .ZN(_0198_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0277_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0198_),
    .B(_0197_),
    .C(_0196_),
    .ZN(_0199_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0278_ (.I0(Tile_X0Y1_E1END[2]),
    .I1(_0195_),
    .I2(Tile_X0Y1_E6END[6]),
    .I3(_0199_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0279_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2 ),
    .I1(Tile_X0Y1_N4END[6]),
    .I2(Tile_X0Y0_S1END[2]),
    .I3(Tile_X0Y0_S4END[2]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit4.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit5.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0280_ (.I0(Tile_X0Y0_E1END[2]),
    .I1(Tile_X0Y0_E6END[6]),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .I3(_0193_),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit2.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit3.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0281_ (.A1(Tile_X0Y0_E6END[3]),
    .A2(_0147_),
    .ZN(_0200_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0282_ (.A1(_0147_),
    .A2(Tile_X0Y0_S1END[3]),
    .ZN(_0201_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0283_ (.A1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ),
    .A2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ),
    .A3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3 ),
    .ZN(_0202_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0284_ (.A1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_0201_),
    .B(_0202_),
    .C(_0200_),
    .ZN(_0203_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0285_ (.I0(Tile_X0Y0_E1END[3]),
    .I1(Tile_X0Y0_E6END[11]),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .I3(_0203_),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit8.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit9.Q ),
    .Z(_0204_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0286_ (.I0(Tile_X0Y1_N1END[3]),
    .I1(Tile_X0Y1_N4END[3]),
    .I2(_0204_),
    .I3(Tile_X0Y0_S4END[7]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q ),
    .Z(_0205_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0287_ (.A1(Tile_X0Y1_E6END[3]),
    .A2(_0159_),
    .ZN(_0206_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0288_ (.A1(_0159_),
    .A2(_0204_),
    .ZN(_0207_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0289_ (.A1(Tile_X0Y1_N1END[3]),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .A3(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .ZN(_0208_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0290_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_0207_),
    .B(_0208_),
    .C(_0206_),
    .ZN(_0209_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0291_ (.I0(Tile_X0Y1_E1END[3]),
    .I1(_0205_),
    .I2(Tile_X0Y1_E6END[7]),
    .I3(_0209_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0292_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3 ),
    .I1(Tile_X0Y1_N4END[7]),
    .I2(Tile_X0Y0_S1END[3]),
    .I3(Tile_X0Y0_S4END[3]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit6.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit7.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0293_ (.I0(Tile_X0Y0_E1END[3]),
    .I1(Tile_X0Y0_E6END[7]),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .I3(_0203_),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit4.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit5.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0294_ (.I0(Tile_X0Y0_E2MID[7]),
    .I1(Tile_X0Y0_E2END[7]),
    .I2(Tile_X0Y0_E6END[7]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit6.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit7.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0295_ (.I0(Tile_X0Y0_E2MID[6]),
    .I1(Tile_X0Y0_E2END[6]),
    .I2(Tile_X0Y0_E6END[9]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit12.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit13.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0296_ (.I0(Tile_X0Y1_N2MID[1]),
    .I1(Tile_X0Y1_N2END[1]),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG1 ),
    .I3(Tile_X0Y0_S2MID[1]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q ),
    .Z(_0000_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0297_ (.I0(Tile_X0Y1_E2MID[6]),
    .I1(Tile_X0Y1_E2END[6]),
    .I2(Tile_X0Y1_E6END[6]),
    .I3(_0000_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0298_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb1 ),
    .I1(Tile_X0Y0_S2MID[1]),
    .I2(Tile_X0Y1_N2MID[1]),
    .I3(Tile_X0Y0_S2END[1]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit11.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit10.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0299_ (.I0(Tile_X0Y0_E2MID[6]),
    .I1(Tile_X0Y0_E2END[6]),
    .I2(Tile_X0Y0_E6END[6]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit8.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit9.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0300_ (.I0(Tile_X0Y0_E2MID[5]),
    .I1(Tile_X0Y0_E2END[5]),
    .I2(Tile_X0Y0_E6END[10]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit14.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit15.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0301_ (.I0(Tile_X0Y1_N2MID[2]),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG2 ),
    .I2(Tile_X0Y1_N2END[2]),
    .I3(Tile_X0Y0_S2MID[2]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q ),
    .Z(_0001_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0302_ (.I0(Tile_X0Y1_E2MID[5]),
    .I1(Tile_X0Y1_E6END[5]),
    .I2(Tile_X0Y1_E2END[5]),
    .I3(_0001_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0303_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb2 ),
    .I1(Tile_X0Y1_N2MID[2]),
    .I2(Tile_X0Y0_S2MID[2]),
    .I3(Tile_X0Y0_S2END[2]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit12.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit13.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0304_ (.I0(Tile_X0Y0_E2MID[5]),
    .I1(Tile_X0Y0_E2END[5]),
    .I2(Tile_X0Y0_E6END[5]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit10.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit11.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0305_ (.I0(Tile_X0Y0_E2MID[4]),
    .I1(Tile_X0Y0_E2END[4]),
    .I2(Tile_X0Y0_E6END[11]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit16.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit17.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0306_ (.I0(Tile_X0Y1_N2MID[3]),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG3 ),
    .I2(Tile_X0Y1_N2END[3]),
    .I3(Tile_X0Y0_S2MID[3]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .Z(_0002_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0307_ (.I0(Tile_X0Y1_E2MID[4]),
    .I1(Tile_X0Y1_E6END[4]),
    .I2(Tile_X0Y1_E2END[4]),
    .I3(_0002_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0308_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb3 ),
    .I1(Tile_X0Y1_N2MID[3]),
    .I2(Tile_X0Y0_S2MID[3]),
    .I3(Tile_X0Y0_S2END[3]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit14.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit15.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0309_ (.I0(Tile_X0Y0_E2MID[4]),
    .I1(Tile_X0Y0_E2END[4]),
    .I2(Tile_X0Y0_E6END[4]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit12.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit13.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0310_ (.I0(Tile_X0Y0_E1END[0]),
    .I1(Tile_X0Y0_E2END[3]),
    .I2(Tile_X0Y0_E2MID[3]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit19.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit18.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0311_ (.I0(Tile_X0Y1_N2MID[4]),
    .I1(Tile_X0Y1_N2END[4]),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG4 ),
    .I3(Tile_X0Y0_S2MID[4]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q ),
    .Z(_0003_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0312_ (.I0(Tile_X0Y1_E2MID[3]),
    .I1(Tile_X0Y1_E2END[3]),
    .I2(Tile_X0Y1_E6END[3]),
    .I3(_0003_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0313_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb4 ),
    .I1(Tile_X0Y0_S2MID[4]),
    .I2(Tile_X0Y1_N2MID[4]),
    .I3(Tile_X0Y0_S2END[4]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit17.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit16.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0314_ (.I0(Tile_X0Y0_E2MID[3]),
    .I1(Tile_X0Y0_E2END[3]),
    .I2(Tile_X0Y0_E6END[3]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit14.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit15.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0315_ (.I0(Tile_X0Y0_E1END[1]),
    .I1(Tile_X0Y0_E2MID[2]),
    .I2(Tile_X0Y0_E2END[2]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit20.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit21.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0316_ (.I0(Tile_X0Y1_N2MID[5]),
    .I1(Tile_X0Y1_N2END[5]),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG5 ),
    .I3(Tile_X0Y0_S2MID[5]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q ),
    .Z(_0004_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0317_ (.I0(Tile_X0Y1_E2MID[2]),
    .I1(Tile_X0Y1_E6END[2]),
    .I2(Tile_X0Y1_E2END[2]),
    .I3(_0004_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0318_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb5 ),
    .I1(Tile_X0Y0_S2MID[5]),
    .I2(Tile_X0Y1_N2MID[5]),
    .I3(Tile_X0Y0_S2END[5]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit19.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit18.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0319_ (.I0(Tile_X0Y0_E2MID[2]),
    .I1(Tile_X0Y0_E2END[2]),
    .I2(Tile_X0Y0_E6END[2]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit16.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit17.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0320_ (.I0(Tile_X0Y0_E1END[2]),
    .I1(Tile_X0Y0_E2MID[1]),
    .I2(Tile_X0Y0_E2END[1]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit22.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit23.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0321_ (.I0(Tile_X0Y1_N2MID[6]),
    .I1(Tile_X0Y1_N2END[6]),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG6 ),
    .I3(Tile_X0Y0_S2MID[6]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q ),
    .Z(_0005_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0322_ (.I0(Tile_X0Y1_E2MID[1]),
    .I1(Tile_X0Y1_E6END[1]),
    .I2(Tile_X0Y1_E2END[1]),
    .I3(_0005_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0323_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb6 ),
    .I1(Tile_X0Y0_S2MID[6]),
    .I2(Tile_X0Y1_N2MID[6]),
    .I3(Tile_X0Y0_S2END[6]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit21.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit20.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0324_ (.I0(Tile_X0Y0_E2MID[1]),
    .I1(Tile_X0Y0_E2END[1]),
    .I2(Tile_X0Y0_E6END[1]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0325_ (.I0(Tile_X0Y0_E1END[3]),
    .I1(Tile_X0Y0_E2MID[0]),
    .I2(Tile_X0Y0_E2END[0]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit24.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit25.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0326_ (.I0(Tile_X0Y1_N2MID[7]),
    .I1(Tile_X0Y1_N2END[7]),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG7 ),
    .I3(Tile_X0Y0_S2MID[7]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q ),
    .Z(_0006_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0327_ (.I0(Tile_X0Y1_E2MID[0]),
    .I1(Tile_X0Y1_E2END[0]),
    .I2(Tile_X0Y1_E6END[0]),
    .I3(_0006_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0328_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb7 ),
    .I1(Tile_X0Y0_S2MID[7]),
    .I2(Tile_X0Y1_N2MID[7]),
    .I3(Tile_X0Y0_S2END[7]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit23.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit22.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0329_ (.I0(Tile_X0Y0_E2MID[0]),
    .I1(Tile_X0Y0_E2END[0]),
    .I2(Tile_X0Y0_E6END[0]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit20.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0330_ (.A1(Tile_X0Y0_E6END[0]),
    .A2(_0155_),
    .ZN(_0007_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0331_ (.A1(Tile_X0Y0_S1END[0]),
    .A2(_0155_),
    .ZN(_0008_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0332_ (.A1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ),
    .A2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ),
    .A3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0 ),
    .ZN(_0009_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0333_ (.A1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(_0008_),
    .B(_0009_),
    .C(_0007_),
    .ZN(_0010_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0334_ (.I0(Tile_X0Y0_E1END[0]),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .I2(Tile_X0Y0_E6END[8]),
    .I3(_0010_),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit3.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit2.Q ),
    .Z(_0011_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0335_ (.I0(Tile_X0Y1_N1END[0]),
    .I1(Tile_X0Y1_N4END[0]),
    .I2(_0011_),
    .I3(Tile_X0Y0_S4END[4]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q ),
    .Z(_0012_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0336_ (.A1(_0156_),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .A3(_0011_),
    .ZN(_0013_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0337_ (.A1(Tile_X0Y1_N1END[0]),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .ZN(_0014_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0338_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(_0014_),
    .ZN(_0015_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0339_ (.A1(Tile_X0Y1_E6END[0]),
    .A2(_0156_),
    .B(_0015_),
    .ZN(_0016_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0340_ (.A1(_0013_),
    .A2(_0016_),
    .ZN(_0017_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0341_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(_0013_),
    .A3(_0016_),
    .Z(_0018_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0342_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(_0012_),
    .B(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .ZN(_0019_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0343_ (.A1(_0154_),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .ZN(_0020_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0344_ (.A1(Tile_X0Y1_E1END[0]),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .B(_0020_),
    .ZN(_0021_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0345_ (.A1(_0018_),
    .A2(_0019_),
    .B1(_0021_),
    .B2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .ZN(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0346_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0 ),
    .I1(Q_SRAM4),
    .I2(Tile_X0Y0_S1END[0]),
    .I3(Q_SRAM6),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit7.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit6.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0347_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1 ),
    .I1(Q_SRAM5),
    .I2(Tile_X0Y0_S1END[1]),
    .I3(Q_SRAM7),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit9.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit8.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0348_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2 ),
    .I1(Q_SRAM4),
    .I2(Tile_X0Y0_S1END[2]),
    .I3(Q_SRAM6),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit11.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit10.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0349_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3 ),
    .I1(Q_SRAM5),
    .I2(Tile_X0Y0_S1END[3]),
    .I3(Q_SRAM7),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit13.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit12.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0350_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit14.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit15.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0351_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .I2(Q_SRAM6),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit17.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit16.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0352_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .I2(Q_SRAM6),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit19.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit18.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0353_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit20.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit21.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0354_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit22.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit23.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0355_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .I2(Q_SRAM6),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit25.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit24.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0356_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .I2(Q_SRAM6),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit27.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit26.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0357_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit28.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit29.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0358_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit30.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit31.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0359_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .I2(Q_SRAM6),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit1.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit0.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0360_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .I2(Q_SRAM6),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit3.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit2.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0361_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit5.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0362_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit6.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit7.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0363_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .I2(Q_SRAM6),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit9.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit8.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0364_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .I2(Q_SRAM6),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit11.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit10.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0365_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit13.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0366_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit14.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit15.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0367_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .I2(Q_SRAM6),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit17.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit16.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0368_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .I2(Q_SRAM6),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit19.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit18.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0369_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0 ),
    .I1(Tile_X0Y1_N4END[4]),
    .I2(Tile_X0Y0_S1END[0]),
    .I3(Tile_X0Y0_S4END[0]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit0.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit1.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0370_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit21.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0371_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3 ),
    .I1(Tile_X0Y1_N4END[7]),
    .I2(Tile_X0Y0_S1END[3]),
    .I3(Tile_X0Y0_S4END[3]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit30.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit31.Q ),
    .Z(_0022_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0372_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(_0022_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit22.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit23.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0373_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2 ),
    .I1(Tile_X0Y1_N4END[6]),
    .I2(Tile_X0Y0_S1END[2]),
    .I3(Tile_X0Y0_S4END[2]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit29.Q ),
    .Z(_0023_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0374_ (.I0(Q_SRAM4),
    .I1(Q_SRAM6),
    .I2(_0023_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit25.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0375_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1 ),
    .I1(Tile_X0Y1_N4END[5]),
    .I2(Tile_X0Y0_S1END[1]),
    .I3(Tile_X0Y0_S4END[1]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit26.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit27.Q ),
    .Z(_0024_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0376_ (.I0(Q_SRAM5),
    .I1(_0024_),
    .I2(Q_SRAM6),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit27.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit26.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0377_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0 ),
    .I1(Tile_X0Y1_N4END[4]),
    .I2(Tile_X0Y0_S1END[0]),
    .I3(Tile_X0Y0_S4END[0]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit25.Q ),
    .Z(_0025_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0378_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(_0025_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit29.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0379_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3 ),
    .I1(Tile_X0Y1_N4END[7]),
    .I2(Tile_X0Y0_S1END[3]),
    .I3(Tile_X0Y0_S4END[3]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit23.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0380_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit31.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG8 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0381_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2 ),
    .I1(Tile_X0Y1_N4END[6]),
    .I2(Tile_X0Y0_S1END[2]),
    .I3(Tile_X0Y0_S4END[2]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit21.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0382_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .I2(Q_SRAM6),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit1.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit0.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG9 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0383_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1 ),
    .I1(Tile_X0Y1_N4END[5]),
    .I2(Tile_X0Y0_S1END[1]),
    .I3(Tile_X0Y0_S4END[1]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit19.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0384_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .I2(Q_SRAM6),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit3.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit2.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG10 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0385_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0 ),
    .I1(Tile_X0Y1_N4END[4]),
    .I2(Tile_X0Y0_S1END[0]),
    .I3(Tile_X0Y0_S4END[0]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit17.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0386_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit5.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG11 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0387_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3 ),
    .I1(Tile_X0Y1_N4END[7]),
    .I2(Tile_X0Y0_S1END[3]),
    .I3(Tile_X0Y0_S4END[3]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit15.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0388_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit7.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG12 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0389_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2 ),
    .I1(Tile_X0Y1_N4END[6]),
    .I2(Tile_X0Y0_S1END[2]),
    .I3(Tile_X0Y0_S4END[2]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit13.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0390_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .I2(Q_SRAM6),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit9.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit8.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG13 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0391_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1 ),
    .I1(Tile_X0Y1_N4END[5]),
    .I2(Tile_X0Y0_S1END[1]),
    .I3(Tile_X0Y0_S4END[1]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit11.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0392_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .I2(Q_SRAM6),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit11.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit10.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG14 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0393_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0 ),
    .I1(Tile_X0Y1_N4END[4]),
    .I2(Tile_X0Y0_S1END[0]),
    .I3(Tile_X0Y0_S4END[0]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit9.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0394_ (.I0(Q_SRAM4),
    .I1(Q_SRAM7),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit13.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG15 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0395_ (.I0(Tile_X0Y1_N4END[4]),
    .I1(Tile_X0Y0_S4END[0]),
    .I2(_0022_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit15.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0396_ (.I0(Tile_X0Y1_N4END[5]),
    .I1(Tile_X0Y0_S4END[1]),
    .I2(_0023_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit17.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0397_ (.I0(Tile_X0Y1_N4END[6]),
    .I1(Tile_X0Y0_S4END[2]),
    .I2(_0024_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit19.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0398_ (.I0(Tile_X0Y1_N4END[7]),
    .I1(Tile_X0Y0_S4END[3]),
    .I2(_0025_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit21.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0399_ (.I0(Q_SRAM7),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .I2(_0022_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit23.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0400_ (.I0(Q_SRAM6),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .I2(_0023_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit25.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0401_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .I2(_0024_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit26.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit27.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0402_ (.I0(Q_SRAM4),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .I2(_0025_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit29.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0403_ (.I0(Q_SRAM4),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit31.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit30.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG8 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0404_ (.I0(Q_SRAM5),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit1.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit0.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG9 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0405_ (.I0(Q_SRAM6),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit3.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit2.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG10 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0406_ (.I0(Q_SRAM7),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .I2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit5.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit4.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG11 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0407_ (.A1(_0149_),
    .A2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .ZN(_0026_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0408_ (.A1(Tile_X0Y0_E2MID[0]),
    .A2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ),
    .A3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ),
    .ZN(_0027_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0409_ (.A1(Tile_X0Y0_E2END[0]),
    .A2(_0149_),
    .ZN(_0028_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0410_ (.A1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ),
    .A2(_0028_),
    .B(_0027_),
    .C(_0026_),
    .ZN(net5),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0411_ (.A1(_0150_),
    .A2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .ZN(_0029_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0412_ (.A1(Tile_X0Y0_E2MID[1]),
    .A2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ),
    .A3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ),
    .ZN(_0030_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0413_ (.A1(Tile_X0Y0_E2END[1]),
    .A2(_0150_),
    .ZN(_0031_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0414_ (.A1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ),
    .A2(_0031_),
    .B(_0030_),
    .C(_0029_),
    .ZN(net6),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0415_ (.A1(_0151_),
    .A2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .ZN(_0032_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0416_ (.A1(Tile_X0Y0_E2MID[2]),
    .A2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ),
    .A3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ),
    .ZN(_0033_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0417_ (.A1(Tile_X0Y0_E2END[2]),
    .A2(_0151_),
    .ZN(_0034_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0418_ (.A1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ),
    .A2(_0034_),
    .B(_0033_),
    .C(_0032_),
    .ZN(net7),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0419_ (.A1(_0152_),
    .A2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .ZN(_0035_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0420_ (.A1(Tile_X0Y0_E2MID[3]),
    .A2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ),
    .A3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ),
    .ZN(_0036_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0421_ (.A1(Tile_X0Y0_E2END[3]),
    .A2(_0152_),
    .ZN(_0037_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0422_ (.A1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ),
    .A2(_0037_),
    .B(_0036_),
    .C(_0035_),
    .ZN(net8),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0423_ (.A1(_0153_),
    .A2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .ZN(_0038_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0424_ (.A1(Tile_X0Y0_E2MID[4]),
    .A2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ),
    .A3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ),
    .ZN(_0039_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0425_ (.A1(_0148_),
    .A2(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ),
    .B1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ),
    .B2(_0038_),
    .C(_0039_),
    .ZN(net9),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0426_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .I2(_0025_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ),
    .Z(_0040_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0427_ (.I0(Tile_X0Y0_E1END[0]),
    .I1(Tile_X0Y0_EE4END[0]),
    .I2(Tile_X0Y0_E6END[8]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ),
    .Z(_0041_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0428_ (.I0(_0041_),
    .I1(_0040_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0429_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .I2(_0024_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ),
    .Z(_0042_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0430_ (.I0(Tile_X0Y0_E1END[1]),
    .I1(Tile_X0Y0_E6END[9]),
    .I2(Tile_X0Y0_EE4END[1]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ),
    .Z(_0043_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0431_ (.I0(_0043_),
    .I1(_0042_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0432_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .I2(_0023_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ),
    .Z(_0044_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0433_ (.I0(Tile_X0Y0_E1END[2]),
    .I1(Tile_X0Y0_E6END[10]),
    .I2(Tile_X0Y0_EE4END[2]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ),
    .Z(_0045_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0434_ (.I0(_0045_),
    .I1(_0044_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit30.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0435_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .I2(_0022_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit0.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit31.Q ),
    .Z(_0046_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0436_ (.I0(Tile_X0Y0_E1END[3]),
    .I1(Tile_X0Y0_E6END[11]),
    .I2(Tile_X0Y0_EE4END[3]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit0.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit31.Q ),
    .Z(_0047_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0437_ (.I0(_0047_),
    .I1(_0046_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit1.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0438_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .I2(_0025_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit27.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit26.Q ),
    .Z(_0048_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0439_ (.I0(Tile_X0Y0_E1END[0]),
    .I1(Tile_X0Y0_EE4END[12]),
    .I2(Tile_X0Y0_E6END[4]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit26.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit27.Q ),
    .Z(_0049_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0440_ (.I0(_0049_),
    .I1(_0048_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit28.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0441_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .I2(_0024_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit30.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit29.Q ),
    .Z(_0050_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0442_ (.I0(Tile_X0Y0_E1END[1]),
    .I1(Tile_X0Y0_E6END[5]),
    .I2(Tile_X0Y0_EE4END[13]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit30.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit29.Q ),
    .Z(_0051_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0443_ (.I0(_0051_),
    .I1(_0050_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit31.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0444_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .I2(_0023_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit1.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit0.Q ),
    .Z(_0052_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0445_ (.I0(Tile_X0Y0_E1END[2]),
    .I1(Tile_X0Y0_E6END[6]),
    .I2(Tile_X0Y0_EE4END[14]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit1.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit0.Q ),
    .Z(_0053_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0446_ (.I0(_0053_),
    .I1(_0052_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit2.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0447_ (.I0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .I2(_0022_),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit4.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit3.Q ),
    .Z(_0054_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0448_ (.I0(Tile_X0Y0_E1END[3]),
    .I1(Tile_X0Y0_E6END[7]),
    .I2(Tile_X0Y0_EE4END[15]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit4.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit3.Q ),
    .Z(_0055_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0449_ (.I0(_0055_),
    .I1(_0054_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit5.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0450_ (.I0(Tile_X0Y0_E6END[0]),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .I2(Tile_X0Y0_E6END[4]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit7.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit6.Q ),
    .Z(_0056_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0451_ (.I0(Tile_X0Y0_EE4END[0]),
    .I1(Tile_X0Y0_EE4END[4]),
    .I2(Tile_X0Y0_EE4END[8]),
    .I3(Tile_X0Y0_EE4END[12]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit7.Q ),
    .Z(_0057_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0452_ (.I0(_0057_),
    .I1(_0056_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit8.Q ),
    .Z(net16),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0453_ (.I0(Tile_X0Y0_E6END[1]),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .I2(Tile_X0Y0_E6END[5]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit9.Q ),
    .Z(_0058_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0454_ (.I0(Tile_X0Y0_EE4END[1]),
    .I1(Tile_X0Y0_EE4END[5]),
    .I2(Tile_X0Y0_EE4END[9]),
    .I3(Tile_X0Y0_EE4END[13]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit9.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit10.Q ),
    .Z(_0059_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0455_ (.I0(_0059_),
    .I1(_0058_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit11.Q ),
    .Z(net17),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0456_ (.I0(Tile_X0Y0_E6END[2]),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .I2(Tile_X0Y0_E6END[6]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit13.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit12.Q ),
    .Z(_0060_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0457_ (.I0(Tile_X0Y0_EE4END[2]),
    .I1(Tile_X0Y0_EE4END[6]),
    .I2(Tile_X0Y0_EE4END[10]),
    .I3(Tile_X0Y0_EE4END[14]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit13.Q ),
    .Z(_0061_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0458_ (.I0(_0061_),
    .I1(_0060_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit14.Q ),
    .Z(net18),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0459_ (.I0(Tile_X0Y0_E6END[3]),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .I2(Tile_X0Y0_E6END[7]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit15.Q ),
    .Z(_0062_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0460_ (.I0(Tile_X0Y0_EE4END[3]),
    .I1(Tile_X0Y0_EE4END[7]),
    .I2(Tile_X0Y0_EE4END[11]),
    .I3(Tile_X0Y0_EE4END[15]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit15.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit16.Q ),
    .Z(_0063_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0461_ (.I0(_0063_),
    .I1(_0062_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit17.Q ),
    .Z(net19),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0462_ (.I0(Tile_X0Y0_E6END[0]),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .I2(Tile_X0Y0_E6END[4]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit19.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit18.Q ),
    .Z(_0064_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0463_ (.I0(Tile_X0Y0_EE4END[0]),
    .I1(Tile_X0Y0_EE4END[4]),
    .I2(Tile_X0Y0_EE4END[8]),
    .I3(Tile_X0Y0_EE4END[12]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit18.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit19.Q ),
    .Z(_0065_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0464_ (.I0(_0065_),
    .I1(_0064_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit20.Q ),
    .Z(net278),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0465_ (.I0(Tile_X0Y0_E6END[1]),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .I2(Tile_X0Y0_E6END[5]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit22.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit21.Q ),
    .Z(_0066_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0466_ (.I0(Tile_X0Y0_EE4END[1]),
    .I1(Tile_X0Y0_EE4END[5]),
    .I2(Tile_X0Y0_EE4END[9]),
    .I3(Tile_X0Y0_EE4END[13]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit21.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit22.Q ),
    .Z(_0067_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0467_ (.I0(_0067_),
    .I1(_0066_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit23.Q ),
    .Z(net279),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0468_ (.I0(Tile_X0Y0_E6END[2]),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .I2(Tile_X0Y0_E6END[6]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit25.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit24.Q ),
    .Z(_0068_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0469_ (.I0(Tile_X0Y0_EE4END[2]),
    .I1(Tile_X0Y0_EE4END[6]),
    .I2(Tile_X0Y0_EE4END[10]),
    .I3(Tile_X0Y0_EE4END[14]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit25.Q ),
    .Z(_0069_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0470_ (.I0(_0069_),
    .I1(_0068_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit26.Q ),
    .Z(net280),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0471_ (.I0(Tile_X0Y0_E6END[3]),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .I2(Tile_X0Y0_E6END[7]),
    .I3(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit27.Q ),
    .Z(_0070_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0472_ (.I0(Tile_X0Y0_EE4END[3]),
    .I1(Tile_X0Y0_EE4END[7]),
    .I2(Tile_X0Y0_EE4END[11]),
    .I3(Tile_X0Y0_EE4END[15]),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit28.Q ),
    .Z(_0071_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0473_ (.I0(_0071_),
    .I1(_0070_),
    .S(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit29.Q ),
    .Z(net281),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0474_ (.I0(Tile_X0Y0_E1END[0]),
    .I1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .I2(Tile_X0Y0_E6END[4]),
    .I3(_0010_),
    .S0(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame8_bit31.Q ),
    .S1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame8_bit30.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0475_ (.I0(Tile_X0Y1_E1END[0]),
    .I1(Tile_X0Y1_E6END[8]),
    .I2(_0012_),
    .I3(_0017_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0476_ (.I0(Tile_X0Y1_E1END[1]),
    .I1(Tile_X0Y1_E6END[9]),
    .I2(_0185_),
    .I3(_0189_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0477_ (.I0(Tile_X0Y1_E1END[2]),
    .I1(Tile_X0Y1_E6END[10]),
    .I2(_0195_),
    .I3(_0199_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0478_ (.I0(Tile_X0Y1_E1END[3]),
    .I1(Tile_X0Y1_E6END[11]),
    .I2(_0205_),
    .I3(_0209_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0479_ (.I0(Tile_X0Y1_E2MID[7]),
    .I1(Tile_X0Y1_E2END[7]),
    .I2(Tile_X0Y1_E6END[8]),
    .I3(_0165_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0480_ (.I0(Tile_X0Y1_E2MID[6]),
    .I1(Tile_X0Y1_E2END[6]),
    .I2(Tile_X0Y1_E6END[9]),
    .I3(_0000_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0481_ (.I0(Tile_X0Y1_E2MID[5]),
    .I1(Tile_X0Y1_E6END[10]),
    .I2(Tile_X0Y1_E2END[5]),
    .I3(_0001_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0482_ (.I0(Tile_X0Y1_E2MID[4]),
    .I1(Tile_X0Y1_E6END[11]),
    .I2(Tile_X0Y1_E2END[4]),
    .I3(_0002_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0483_ (.I0(Tile_X0Y1_E1END[0]),
    .I1(Tile_X0Y1_E2END[3]),
    .I2(Tile_X0Y1_E2MID[3]),
    .I3(_0003_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0484_ (.I0(Tile_X0Y1_E1END[1]),
    .I1(Tile_X0Y1_E2MID[2]),
    .I2(Tile_X0Y1_E2END[2]),
    .I3(_0004_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0485_ (.I0(Tile_X0Y1_E1END[2]),
    .I1(Tile_X0Y1_E2MID[1]),
    .I2(Tile_X0Y1_E2END[1]),
    .I3(_0005_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0486_ (.I0(Tile_X0Y1_E1END[3]),
    .I1(Tile_X0Y1_E2END[0]),
    .I2(Tile_X0Y1_E2MID[0]),
    .I3(_0006_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0487_ (.I0(Tile_X0Y1_N1END[0]),
    .I1(Q_SRAM0),
    .I2(_0011_),
    .I3(Q_SRAM2),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0488_ (.I0(Tile_X0Y1_N1END[1]),
    .I1(Q_SRAM1),
    .I2(_0184_),
    .I3(Q_SRAM3),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0489_ (.I0(Tile_X0Y1_N1END[2]),
    .I1(Q_SRAM0),
    .I2(_0194_),
    .I3(Q_SRAM2),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0490_ (.I0(Tile_X0Y1_N1END[3]),
    .I1(Q_SRAM1),
    .I2(_0204_),
    .I3(Q_SRAM3),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0491_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(_0165_),
    .I3(_0006_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0492_ (.I0(Q_SRAM1),
    .I1(_0000_),
    .I2(Q_SRAM2),
    .I3(_0005_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0493_ (.I0(Q_SRAM1),
    .I1(_0001_),
    .I2(Q_SRAM2),
    .I3(_0004_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0494_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(_0002_),
    .I3(_0003_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0495_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(_0002_),
    .I3(_0003_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0496_ (.I0(Q_SRAM1),
    .I1(_0001_),
    .I2(Q_SRAM2),
    .I3(_0004_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0497_ (.I0(Q_SRAM1),
    .I1(_0000_),
    .I2(Q_SRAM2),
    .I3(_0005_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0498_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(_0165_),
    .I3(_0006_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0499_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(_0165_),
    .I3(_0006_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0500_ (.I0(Q_SRAM1),
    .I1(_0000_),
    .I2(Q_SRAM2),
    .I3(_0005_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0501_ (.I0(Q_SRAM1),
    .I1(_0001_),
    .I2(Q_SRAM2),
    .I3(_0004_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0502_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(_0002_),
    .I3(_0003_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0503_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(_0002_),
    .I3(_0003_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0504_ (.I0(Q_SRAM1),
    .I1(_0001_),
    .I2(Q_SRAM2),
    .I3(_0004_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0505_ (.I0(Q_SRAM1),
    .I1(_0000_),
    .I2(Q_SRAM2),
    .I3(_0005_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0506_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(_0165_),
    .I3(_0006_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0507_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(_0205_),
    .I3(_0006_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0508_ (.I0(Q_SRAM1),
    .I1(_0195_),
    .I2(Q_SRAM2),
    .I3(_0005_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0509_ (.I0(Q_SRAM1),
    .I1(_0185_),
    .I2(Q_SRAM2),
    .I3(_0004_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0510_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(_0012_),
    .I3(_0003_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0511_ (.I0(Tile_X0Y1_N1END[3]),
    .I1(Tile_X0Y1_N4END[3]),
    .I2(_0204_),
    .I3(Tile_X0Y0_S4END[7]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q ),
    .Z(_0072_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0512_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(_0072_),
    .I3(_0002_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0513_ (.I0(Tile_X0Y1_N1END[2]),
    .I1(Tile_X0Y1_N4END[2]),
    .I2(_0194_),
    .I3(Tile_X0Y0_S4END[6]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .Z(_0073_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0514_ (.I0(Q_SRAM1),
    .I1(_0073_),
    .I2(Q_SRAM2),
    .I3(_0001_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0515_ (.I0(Tile_X0Y1_N1END[1]),
    .I1(Tile_X0Y1_N4END[1]),
    .I2(_0184_),
    .I3(Tile_X0Y0_S4END[5]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q ),
    .Z(_0074_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0516_ (.I0(Q_SRAM1),
    .I1(_0074_),
    .I2(Q_SRAM2),
    .I3(_0000_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0517_ (.I0(Tile_X0Y1_N1END[0]),
    .I1(Tile_X0Y1_N4END[0]),
    .I2(_0011_),
    .I3(Tile_X0Y0_S4END[4]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .Z(_0075_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0518_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(_0075_),
    .I3(_0165_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0519_ (.I0(Tile_X0Y1_N1END[3]),
    .I1(Tile_X0Y1_N4END[3]),
    .I2(_0204_),
    .I3(Tile_X0Y0_S4END[7]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0520_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .I3(_0006_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG8 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0521_ (.I0(Tile_X0Y1_N1END[2]),
    .I1(Tile_X0Y1_N4END[2]),
    .I2(_0194_),
    .I3(Tile_X0Y0_S4END[6]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0522_ (.I0(Q_SRAM1),
    .I1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .I2(Q_SRAM2),
    .I3(_0005_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG9 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0523_ (.I0(Tile_X0Y1_N1END[1]),
    .I1(Tile_X0Y1_N4END[1]),
    .I2(_0184_),
    .I3(Tile_X0Y0_S4END[5]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0524_ (.I0(Q_SRAM1),
    .I1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .I2(Q_SRAM2),
    .I3(_0004_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG10 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0525_ (.I0(Tile_X0Y1_N1END[0]),
    .I1(Tile_X0Y1_N4END[0]),
    .I2(_0011_),
    .I3(Tile_X0Y0_S4END[4]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0526_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .I3(_0003_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG11 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0527_ (.I0(Tile_X0Y1_N1END[3]),
    .I1(Tile_X0Y1_N4END[3]),
    .I2(_0204_),
    .I3(Tile_X0Y0_S4END[7]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q ),
    .Z(_0076_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0528_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(_0076_),
    .I3(_0002_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG12 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0529_ (.I0(Tile_X0Y1_N1END[2]),
    .I1(Tile_X0Y1_N4END[2]),
    .I2(_0194_),
    .I3(Tile_X0Y0_S4END[6]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .Z(_0077_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0530_ (.I0(Q_SRAM1),
    .I1(_0077_),
    .I2(Q_SRAM2),
    .I3(_0001_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG13 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0531_ (.I0(Tile_X0Y1_N1END[1]),
    .I1(Tile_X0Y1_N4END[1]),
    .I2(_0184_),
    .I3(Tile_X0Y0_S4END[5]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q ),
    .Z(_0078_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0532_ (.I0(Q_SRAM1),
    .I1(_0078_),
    .I2(Q_SRAM2),
    .I3(_0000_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG14 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0533_ (.I0(Tile_X0Y1_N1END[0]),
    .I1(Tile_X0Y1_N4END[0]),
    .I2(_0011_),
    .I3(Tile_X0Y0_S4END[4]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .Z(_0079_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0534_ (.I0(Q_SRAM0),
    .I1(Q_SRAM3),
    .I2(_0079_),
    .I3(_0165_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG15 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0535_ (.I0(Tile_X0Y1_N4END[0]),
    .I1(Tile_X0Y0_S4END[4]),
    .I2(_0072_),
    .I3(_0205_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0536_ (.I0(Tile_X0Y1_N4END[1]),
    .I1(Tile_X0Y0_S4END[5]),
    .I2(_0073_),
    .I3(_0195_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0537_ (.I0(Tile_X0Y1_N4END[2]),
    .I1(Tile_X0Y0_S4END[6]),
    .I2(_0074_),
    .I3(_0185_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0538_ (.I0(Tile_X0Y1_N4END[3]),
    .I1(Tile_X0Y0_S4END[7]),
    .I2(_0075_),
    .I3(_0012_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0539_ (.I0(Q_SRAM3),
    .I1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .I2(_0072_),
    .I3(_0165_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0540_ (.I0(Q_SRAM2),
    .I1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .I2(_0073_),
    .I3(_0000_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0541_ (.I0(Q_SRAM1),
    .I1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .I2(_0074_),
    .I3(_0001_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0542_ (.I0(Q_SRAM0),
    .I1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .I2(_0075_),
    .I3(_0002_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0543_ (.I0(Q_SRAM0),
    .I1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .I2(_0076_),
    .I3(_0003_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG8 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0544_ (.I0(Q_SRAM1),
    .I1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .I2(_0077_),
    .I3(_0004_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG9 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0545_ (.I0(Q_SRAM2),
    .I1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .I2(_0078_),
    .I3(_0005_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG10 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0546_ (.I0(Q_SRAM3),
    .I1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .I2(_0079_),
    .I3(_0006_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG11 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0547_ (.A1(_0160_),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .A3(_0165_),
    .ZN(_0080_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0548_ (.A1(Tile_X0Y1_E2MID[0]),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .ZN(_0081_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0549_ (.A1(Tile_X0Y1_E2END[0]),
    .A2(_0160_),
    .ZN(_0082_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0550_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .A2(_0081_),
    .A3(_0082_),
    .B(_0080_),
    .ZN(net1),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0551_ (.A1(_0161_),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .A3(_0000_),
    .ZN(_0083_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0552_ (.A1(Tile_X0Y1_E2MID[1]),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .ZN(_0084_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0553_ (.A1(Tile_X0Y1_E2END[1]),
    .A2(_0161_),
    .ZN(_0085_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0554_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .A2(_0084_),
    .A3(_0085_),
    .B(_0083_),
    .ZN(net2),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0555_ (.A1(_0162_),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .A3(_0001_),
    .ZN(_0086_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0556_ (.A1(Tile_X0Y1_E2MID[2]),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .ZN(_0087_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0557_ (.A1(Tile_X0Y1_E2END[2]),
    .A2(_0162_),
    .ZN(_0088_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0558_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .A2(_0087_),
    .A3(_0088_),
    .B(_0086_),
    .ZN(net3),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0559_ (.A1(_0163_),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q ),
    .A3(_0002_),
    .ZN(_0089_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0560_ (.A1(Tile_X0Y1_E2MID[3]),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .ZN(_0090_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0561_ (.A1(Tile_X0Y1_E2END[3]),
    .A2(_0163_),
    .ZN(_0091_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0562_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q ),
    .A2(_0090_),
    .A3(_0091_),
    .B(_0089_),
    .ZN(net4),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0563_ (.I0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .I1(_0012_),
    .I2(_0075_),
    .I3(_0165_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .Z(_0092_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0564_ (.I0(Tile_X0Y1_E1END[0]),
    .I1(Tile_X0Y1_E6END[8]),
    .I2(Tile_X0Y1_EE4END[0]),
    .I3(_0079_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .Z(_0093_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0565_ (.I0(_0093_),
    .I1(_0092_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_8.A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0566_ (.I0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .I1(_0185_),
    .I2(_0074_),
    .I3(_0000_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .Z(_0094_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0567_ (.I0(Tile_X0Y1_E1END[1]),
    .I1(Tile_X0Y1_E6END[9]),
    .I2(Tile_X0Y1_EE4END[1]),
    .I3(_0078_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .Z(_0095_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0568_ (.I0(_0095_),
    .I1(_0094_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_9.A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0569_ (.I0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .I1(_0195_),
    .I2(_0073_),
    .I3(_0001_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q ),
    .Z(_0096_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0570_ (.I0(Tile_X0Y1_E1END[2]),
    .I1(Tile_X0Y1_E6END[10]),
    .I2(Tile_X0Y1_EE4END[2]),
    .I3(_0077_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q ),
    .Z(_0097_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0571_ (.I0(_0097_),
    .I1(_0096_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_10.A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0572_ (.I0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .I1(_0205_),
    .I2(_0072_),
    .I3(_0002_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .Z(_0098_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0573_ (.I0(Tile_X0Y1_E1END[3]),
    .I1(Tile_X0Y1_E6END[11]),
    .I2(Tile_X0Y1_EE4END[3]),
    .I3(_0076_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .Z(_0099_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0574_ (.I0(_0099_),
    .I1(_0098_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q ),
    .Z(\Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_11.A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0575_ (.I0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .I1(_0012_),
    .I2(_0075_),
    .I3(_0003_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q ),
    .Z(_0100_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0576_ (.I0(Tile_X0Y1_E1END[0]),
    .I1(Tile_X0Y1_EE4END[12]),
    .I2(Tile_X0Y1_E6END[4]),
    .I3(_0079_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q ),
    .Z(_0101_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0577_ (.I0(_0101_),
    .I1(_0100_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0578_ (.I0(Tile_X0Y1_E1END[1]),
    .I1(Tile_X0Y1_EE4END[13]),
    .I2(Tile_X0Y1_E6END[5]),
    .I3(_0078_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q ),
    .Z(_0102_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0579_ (.I0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .I1(_0185_),
    .I2(_0074_),
    .I3(_0004_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q ),
    .Z(_0103_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0580_ (.I0(_0102_),
    .I1(_0103_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0581_ (.I0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .I1(_0195_),
    .I2(_0073_),
    .I3(_0005_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q ),
    .Z(_0104_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0582_ (.I0(Tile_X0Y1_E1END[2]),
    .I1(Tile_X0Y1_EE4END[14]),
    .I2(Tile_X0Y1_E6END[6]),
    .I3(_0077_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q ),
    .Z(_0105_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0583_ (.I0(_0105_),
    .I1(_0104_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0584_ (.I0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .I1(_0205_),
    .I2(_0072_),
    .I3(_0006_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q ),
    .Z(_0106_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0585_ (.I0(Tile_X0Y1_E1END[3]),
    .I1(Tile_X0Y1_EE4END[15]),
    .I2(Tile_X0Y1_E6END[7]),
    .I3(_0076_),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .Z(_0107_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0586_ (.I0(_0107_),
    .I1(_0106_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q ),
    .Z(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0587_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .A2(_0164_),
    .ZN(_0108_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0588_ (.I0(Tile_X0Y1_E2END[4]),
    .I1(Tile_X0Y0_S2MID[3]),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .Z(_0109_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _0589_ (.A1(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG0 ),
    .A2(_0108_),
    .B1(_0109_),
    .B2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .C(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .ZN(_0110_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0590_ (.A1(Tile_X0Y1_E2END[5]),
    .A2(_0164_),
    .ZN(_0111_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0591_ (.A1(_0142_),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .B1(_0111_),
    .B2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .C(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .ZN(_0112_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0592_ (.A1(Tile_X0Y1_E2END[3]),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .A3(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .B(_0112_),
    .ZN(_0113_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0593_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .A2(_0110_),
    .A3(_0113_),
    .ZN(_0114_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0594_ (.I0(Tile_X0Y1_E2MID[3]),
    .I1(Tile_X0Y1_E2MID[6]),
    .I2(Tile_X0Y1_E2END[1]),
    .I3(Tile_X0Y1_E2END[2]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .Z(_0115_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0595_ (.A1(_0140_),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .ZN(_0116_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0596_ (.A1(Tile_X0Y1_E2MID[0]),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .B(_0108_),
    .C(_0116_),
    .ZN(_0117_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0597_ (.A1(Tile_X0Y1_N2END[2]),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .B(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .C(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .ZN(_0118_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0598_ (.A1(_0139_),
    .A2(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .B(_0118_),
    .ZN(_0119_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0599_ (.A1(_0164_),
    .A2(_0115_),
    .B(_0119_),
    .ZN(_0120_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0600_ (.A1(_0117_),
    .A2(_0120_),
    .ZN(_0121_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0601_ (.A1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .A2(_0121_),
    .B(_0114_),
    .ZN(_0122_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0602_ (.I(_0122_),
    .ZN(net20),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0603_ (.I0(Tile_X0Y1_E6END[0]),
    .I1(_0079_),
    .I2(Tile_X0Y1_E6END[4]),
    .I3(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .Z(_0123_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0604_ (.I0(Tile_X0Y1_EE4END[0]),
    .I1(Tile_X0Y1_EE4END[4]),
    .I2(Tile_X0Y1_EE4END[8]),
    .I3(Tile_X0Y1_EE4END[12]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .Z(_0124_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0605_ (.I0(_0124_),
    .I1(_0123_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .Z(net274),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0606_ (.I0(Tile_X0Y1_E6END[1]),
    .I1(_0078_),
    .I2(Tile_X0Y1_E6END[5]),
    .I3(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .Z(_0125_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0607_ (.I0(Tile_X0Y1_EE4END[1]),
    .I1(Tile_X0Y1_EE4END[5]),
    .I2(Tile_X0Y1_EE4END[9]),
    .I3(Tile_X0Y1_EE4END[13]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .Z(_0126_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0608_ (.I0(_0126_),
    .I1(_0125_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .Z(net275),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0609_ (.I0(Tile_X0Y1_E6END[2]),
    .I1(_0077_),
    .I2(Tile_X0Y1_E6END[6]),
    .I3(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .Z(_0127_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0610_ (.I0(Tile_X0Y1_EE4END[2]),
    .I1(Tile_X0Y1_EE4END[6]),
    .I2(Tile_X0Y1_EE4END[10]),
    .I3(Tile_X0Y1_EE4END[14]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .Z(_0128_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0611_ (.I0(_0128_),
    .I1(_0127_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .Z(net276),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0612_ (.I0(Tile_X0Y1_E6END[3]),
    .I1(_0076_),
    .I2(Tile_X0Y1_E6END[7]),
    .I3(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .Z(_0129_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0613_ (.I0(Tile_X0Y1_EE4END[3]),
    .I1(Tile_X0Y1_EE4END[7]),
    .I2(Tile_X0Y1_EE4END[11]),
    .I3(Tile_X0Y1_EE4END[15]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .Z(_0130_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0614_ (.I0(_0130_),
    .I1(_0129_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q ),
    .Z(net277),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0615_ (.I0(Tile_X0Y1_E6END[0]),
    .I1(_0079_),
    .I2(Tile_X0Y1_E6END[4]),
    .I3(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .Z(_0131_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0616_ (.I0(Tile_X0Y1_EE4END[0]),
    .I1(Tile_X0Y1_EE4END[4]),
    .I2(Tile_X0Y1_EE4END[8]),
    .I3(Tile_X0Y1_EE4END[12]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .Z(_0132_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0617_ (.I0(_0132_),
    .I1(_0131_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .Z(net12),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0618_ (.I0(Tile_X0Y1_E6END[1]),
    .I1(_0078_),
    .I2(Tile_X0Y1_E6END[5]),
    .I3(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .Z(_0133_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0619_ (.I0(Tile_X0Y1_EE4END[1]),
    .I1(Tile_X0Y1_EE4END[5]),
    .I2(Tile_X0Y1_EE4END[9]),
    .I3(Tile_X0Y1_EE4END[13]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .Z(_0134_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0620_ (.I0(_0134_),
    .I1(_0133_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .Z(net13),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0621_ (.I0(Tile_X0Y1_E6END[2]),
    .I1(_0077_),
    .I2(Tile_X0Y1_E6END[6]),
    .I3(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .Z(_0135_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0622_ (.I0(Tile_X0Y1_EE4END[2]),
    .I1(Tile_X0Y1_EE4END[6]),
    .I2(Tile_X0Y1_EE4END[10]),
    .I3(Tile_X0Y1_EE4END[14]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q ),
    .Z(_0136_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0623_ (.I0(_0136_),
    .I1(_0135_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .Z(net14),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0624_ (.I0(Tile_X0Y1_E6END[3]),
    .I1(_0076_),
    .I2(Tile_X0Y1_E6END[7]),
    .I3(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .Z(_0137_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0625_ (.I0(Tile_X0Y1_EE4END[3]),
    .I1(Tile_X0Y1_EE4END[7]),
    .I2(Tile_X0Y1_EE4END[11]),
    .I3(Tile_X0Y1_EE4END[15]),
    .S0(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .S1(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .Z(_0138_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0626_ (.I0(_0138_),
    .I1(_0137_),
    .S(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .Z(net15),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0627_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0628_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0629_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0630_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0631_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0632_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0633_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0634_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0635_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0636_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0637_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0638_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0639_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0640_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0641_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0642_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0643_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0644_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0645_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0646_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0647_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0648_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0649_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0650_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0651_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0652_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0653_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0654_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0655_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0656_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0657_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0658_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0659_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0660_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0661_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0662_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0663_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0664_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0665_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0666_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0667_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0668_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0669_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0670_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0671_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0672_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0673_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0674_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0675_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0676_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0677_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0678_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0679_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0680_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0681_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0682_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0683_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0684_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0685_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0686_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0687_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0688_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0689_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0690_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0691_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0692_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0693_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0694_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0695_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0696_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0697_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0698_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0699_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0700_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0701_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0702_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0703_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0704_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0705_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0706_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0707_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0708_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0709_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0710_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0711_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0712_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0713_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0714_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0715_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0716_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0717_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0718_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0719_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0720_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0721_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0722_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0723_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0724_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0725_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0726_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0727_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0728_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0729_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0730_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0731_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0732_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0733_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0734_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0735_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0736_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0737_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0738_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0739_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0740_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0741_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0742_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0743_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0744_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0745_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0746_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0747_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0748_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0749_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0750_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0751_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0752_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0753_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0754_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0755_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0756_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0757_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0758_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0759_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0760_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0761_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0762_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0763_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0764_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0765_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0766_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0767_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0768_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0769_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0770_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0771_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0772_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0773_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0774_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0775_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0776_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0777_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0778_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0779_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0780_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0781_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0782_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0783_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0784_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0785_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0786_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0787_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0788_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0789_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0790_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0791_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0792_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0793_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0794_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0795_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0796_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0797_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0798_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0799_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0800_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0801_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0802_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0803_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0804_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0805_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0806_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0807_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0808_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0809_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0810_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0811_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0812_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0813_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0814_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0815_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0816_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0817_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0818_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0819_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0820_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0821_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0822_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0823_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0824_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0825_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0826_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0827_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0828_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0829_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0830_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0831_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0832_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0833_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0834_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0835_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0836_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0837_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0838_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0839_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0840_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0841_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0842_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0843_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0844_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0845_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0846_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0847_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0848_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0849_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0850_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0851_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0852_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0853_ (.D(Tile_X0Y0_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0854_ (.D(Tile_X0Y0_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0855_ (.D(Tile_X0Y0_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0856_ (.D(Tile_X0Y0_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0857_ (.D(Tile_X0Y0_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0858_ (.D(Tile_X0Y0_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0859_ (.D(Tile_X0Y0_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0860_ (.D(Tile_X0Y0_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0861_ (.D(Tile_X0Y0_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0862_ (.D(Tile_X0Y0_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0863_ (.D(Tile_X0Y0_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0864_ (.D(Tile_X0Y0_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0865_ (.D(Tile_X0Y0_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0866_ (.D(Tile_X0Y0_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0867_ (.D(Tile_X0Y0_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0868_ (.D(Tile_X0Y0_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0869_ (.D(Tile_X0Y0_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0870_ (.D(Tile_X0Y0_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0871_ (.D(Tile_X0Y0_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0872_ (.D(Tile_X0Y0_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0873_ (.D(Tile_X0Y0_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0874_ (.D(Tile_X0Y0_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0875_ (.D(Tile_X0Y0_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0876_ (.D(Tile_X0Y0_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0877_ (.D(Tile_X0Y0_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0878_ (.D(Tile_X0Y0_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0879_ (.D(Tile_X0Y0_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0880_ (.D(Tile_X0Y0_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0881_ (.D(Tile_X0Y0_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0882_ (.D(Tile_X0Y0_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0883_ (.D(Tile_X0Y0_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame8_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0884_ (.D(Tile_X0Y0_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame8_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0885_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0886_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0887_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0888_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0889_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0890_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0891_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0892_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0893_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0894_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0895_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0896_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0897_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0898_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0899_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0900_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0901_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0902_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0903_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0904_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0905_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0906_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0907_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0908_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0909_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0910_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0911_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0912_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0913_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0914_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0915_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0916_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0917_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0918_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0919_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0920_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0921_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0922_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0923_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0924_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0925_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0926_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0927_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0928_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0929_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0930_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0931_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0932_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0933_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0934_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0935_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0936_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0937_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0938_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0939_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0940_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0941_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0942_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0943_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0944_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0945_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0946_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0947_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0948_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0949_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0950_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0951_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0952_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0953_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0954_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0955_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0956_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0957_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0958_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0959_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0960_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0961_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0962_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0963_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0964_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0965_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0966_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0967_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0968_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0969_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0970_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0971_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0972_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0973_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0974_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0975_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0976_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0977_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0978_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0979_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0980_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0981_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0982_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0983_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0984_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0985_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0986_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0987_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0988_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0989_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0990_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0991_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0992_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0993_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0994_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0995_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0996_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0997_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0998_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _0999_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1000_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1001_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1002_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1003_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1004_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1005_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1006_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1007_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1008_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1009_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1010_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1011_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1012_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1013_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1014_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1015_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1016_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1017_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1018_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1019_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1020_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1021_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1022_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1023_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1024_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1025_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1026_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1027_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1028_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1029_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1030_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1031_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1032_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1033_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1034_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1035_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1036_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1037_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1038_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1039_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1040_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1041_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1042_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1043_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1044_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1045_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1046_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1047_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1048_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1049_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1050_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1051_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1052_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1053_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1054_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1055_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1056_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1057_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1058_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1059_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1060_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1061_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1062_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1063_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1064_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1065_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1066_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1067_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1068_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1069_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1070_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1071_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1072_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1073_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1074_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1075_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1076_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1077_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1078_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1079_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1080_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1081_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1082_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1083_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1084_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1085_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1086_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1087_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1088_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1089_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1090_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1091_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1092_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1093_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1094_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1095_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1096_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1097_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1098_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1099_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1100_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1101_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1102_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1103_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1104_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1105_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1106_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1107_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1108_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1109_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1110_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1111_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1112_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1113_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1114_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1115_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1116_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1117_ (.D(Tile_X0Y1_FrameData[23]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1118_ (.D(Tile_X0Y1_FrameData[22]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1119_ (.D(Tile_X0Y1_FrameData[21]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1120_ (.D(Tile_X0Y1_FrameData[20]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1121_ (.D(Tile_X0Y1_FrameData[19]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1122_ (.D(Tile_X0Y1_FrameData[18]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1123_ (.D(Tile_X0Y1_FrameData[17]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1124_ (.D(Tile_X0Y1_FrameData[16]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1125_ (.D(Tile_X0Y1_FrameData[15]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1126_ (.D(Tile_X0Y1_FrameData[14]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1127_ (.D(Tile_X0Y1_FrameData[13]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1128_ (.D(Tile_X0Y1_FrameData[12]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1129_ (.D(Tile_X0Y1_FrameData[11]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1130_ (.D(Tile_X0Y1_FrameData[10]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1131_ (.D(Tile_X0Y1_FrameData[9]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1132_ (.D(Tile_X0Y1_FrameData[8]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1133_ (.D(Tile_X0Y1_FrameData[7]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1134_ (.D(Tile_X0Y1_FrameData[6]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1135_ (.D(Tile_X0Y1_FrameData[5]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1136_ (.D(Tile_X0Y1_FrameData[4]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1137_ (.D(Tile_X0Y1_FrameData[3]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1138_ (.D(Tile_X0Y1_FrameData[2]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1139_ (.D(Tile_X0Y1_FrameData[1]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1140_ (.D(Tile_X0Y1_FrameData[0]),
    .E(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1141_ (.D(Tile_X0Y1_FrameData[31]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1142_ (.D(Tile_X0Y1_FrameData[30]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1143_ (.D(Tile_X0Y1_FrameData[29]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1144_ (.D(Tile_X0Y1_FrameData[28]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1145_ (.D(Tile_X0Y1_FrameData[27]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1146_ (.D(Tile_X0Y1_FrameData[26]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1147_ (.D(Tile_X0Y1_FrameData[25]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1148_ (.D(Tile_X0Y1_FrameData[24]),
    .E(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1149_ (.I(clknet_1_0__leaf_Tile_X0Y1_UserCLK),
    .Z(net11),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1150_ (.I(Tile_X0Y0_FrameData[0]),
    .Z(net21),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1151_ (.I(Tile_X0Y0_FrameData[1]),
    .Z(net32),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1152_ (.I(Tile_X0Y0_FrameData[2]),
    .Z(net43),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1153_ (.I(Tile_X0Y0_FrameData[3]),
    .Z(net46),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1154_ (.I(Tile_X0Y0_FrameData[4]),
    .Z(net47),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1155_ (.I(Tile_X0Y0_FrameData[5]),
    .Z(net48),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1156_ (.I(Tile_X0Y0_FrameData[6]),
    .Z(net49),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1157_ (.I(Tile_X0Y0_FrameData[7]),
    .Z(net50),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1158_ (.I(Tile_X0Y0_FrameData[8]),
    .Z(net51),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1159_ (.I(Tile_X0Y0_FrameData[9]),
    .Z(net52),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1160_ (.I(Tile_X0Y0_FrameData[10]),
    .Z(net22),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1161_ (.I(Tile_X0Y0_FrameData[11]),
    .Z(net23),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1162_ (.I(Tile_X0Y0_FrameData[12]),
    .Z(net24),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1163_ (.I(Tile_X0Y0_FrameData[13]),
    .Z(net25),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1164_ (.I(Tile_X0Y0_FrameData[14]),
    .Z(net26),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1165_ (.I(Tile_X0Y0_FrameData[15]),
    .Z(net27),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1166_ (.I(Tile_X0Y0_FrameData[16]),
    .Z(net28),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1167_ (.I(Tile_X0Y0_FrameData[17]),
    .Z(net29),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1168_ (.I(Tile_X0Y0_FrameData[18]),
    .Z(net30),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1169_ (.I(Tile_X0Y0_FrameData[19]),
    .Z(net31),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1170_ (.I(Tile_X0Y0_FrameData[20]),
    .Z(net33),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1171_ (.I(Tile_X0Y0_FrameData[21]),
    .Z(net34),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1172_ (.I(Tile_X0Y0_FrameData[22]),
    .Z(net35),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1173_ (.I(Tile_X0Y0_FrameData[23]),
    .Z(net36),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1174_ (.I(Tile_X0Y0_FrameData[24]),
    .Z(net37),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1175_ (.I(Tile_X0Y0_FrameData[25]),
    .Z(net38),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1176_ (.I(Tile_X0Y0_FrameData[26]),
    .Z(net39),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1177_ (.I(Tile_X0Y0_FrameData[27]),
    .Z(net40),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1178_ (.I(Tile_X0Y0_FrameData[28]),
    .Z(net41),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1179_ (.I(Tile_X0Y0_FrameData[29]),
    .Z(net42),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1180_ (.I(Tile_X0Y0_FrameData[30]),
    .Z(net44),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1181_ (.I(Tile_X0Y0_FrameData[31]),
    .Z(net45),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1182_ (.I(Tile_X0Y1_FrameStrobe[0]),
    .Z(net53),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1183_ (.I(Tile_X0Y1_FrameStrobe[1]),
    .Z(net64),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1184_ (.I(Tile_X0Y1_FrameStrobe[2]),
    .Z(net65),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1185_ (.I(Tile_X0Y1_FrameStrobe[3]),
    .Z(net66),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1186_ (.I(Tile_X0Y1_FrameStrobe[4]),
    .Z(net67),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1187_ (.I(Tile_X0Y1_FrameStrobe[5]),
    .Z(net68),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1188_ (.I(Tile_X0Y1_FrameStrobe[6]),
    .Z(net69),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1189_ (.I(Tile_X0Y1_FrameStrobe[7]),
    .Z(net70),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1190_ (.I(Tile_X0Y1_FrameStrobe[8]),
    .Z(net71),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1191_ (.I(Tile_X0Y1_FrameStrobe[9]),
    .Z(net72),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1192_ (.I(Tile_X0Y1_FrameStrobe[10]),
    .Z(net54),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1193_ (.I(Tile_X0Y1_FrameStrobe[11]),
    .Z(net55),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1194_ (.I(Tile_X0Y1_FrameStrobe[12]),
    .Z(net56),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1195_ (.I(Tile_X0Y1_FrameStrobe[13]),
    .Z(net57),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1196_ (.I(Tile_X0Y1_FrameStrobe[14]),
    .Z(net58),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1197_ (.I(Tile_X0Y1_FrameStrobe[15]),
    .Z(net59),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1198_ (.I(Tile_X0Y1_FrameStrobe[16]),
    .Z(net60),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1199_ (.I(Tile_X0Y1_FrameStrobe[17]),
    .Z(net61),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1200_ (.I(Tile_X0Y1_FrameStrobe[18]),
    .Z(net62),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1201_ (.I(Tile_X0Y1_FrameStrobe[19]),
    .Z(net63),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1202_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG0 ),
    .Z(net73),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1203_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG1 ),
    .Z(net74),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1204_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG2 ),
    .Z(net75),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1205_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG3 ),
    .Z(net76),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1206_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG0 ),
    .Z(net77),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1207_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG1 ),
    .Z(net78),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1208_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG2 ),
    .Z(net79),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1209_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG3 ),
    .Z(net80),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1210_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG4 ),
    .Z(net81),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1211_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG5 ),
    .Z(net82),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1212_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG6 ),
    .Z(net83),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1213_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG7 ),
    .Z(net84),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1214_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb0 ),
    .Z(net85),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1215_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb1 ),
    .Z(net86),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1216_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb2 ),
    .Z(net87),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1217_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb3 ),
    .Z(net88),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1218_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb4 ),
    .Z(net89),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1219_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb5 ),
    .Z(net90),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1220_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb6 ),
    .Z(net91),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1221_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb7 ),
    .Z(net92),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1222_ (.I(Tile_X0Y1_N4END[8]),
    .Z(net93),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1223_ (.I(Tile_X0Y1_N4END[9]),
    .Z(net100),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1224_ (.I(Tile_X0Y1_N4END[10]),
    .Z(net101),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1225_ (.I(Tile_X0Y1_N4END[11]),
    .Z(net102),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1226_ (.I(Tile_X0Y1_N4END[12]),
    .Z(net103),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1227_ (.I(Tile_X0Y1_N4END[13]),
    .Z(net104),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1228_ (.I(Tile_X0Y1_N4END[14]),
    .Z(net105),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1229_ (.I(Tile_X0Y1_N4END[15]),
    .Z(net106),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1230_ (.I(\Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_8.A ),
    .Z(net107),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1231_ (.I(\Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_9.A ),
    .Z(net108),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1232_ (.I(\Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_10.A ),
    .Z(net94),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1233_ (.I(\Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_11.A ),
    .Z(net95),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1234_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG0 ),
    .Z(net96),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1235_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG1 ),
    .Z(net97),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1236_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG2 ),
    .Z(net98),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1237_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG3 ),
    .Z(net99),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1238_ (.I(clknet_1_1__leaf_Tile_X0Y1_UserCLK),
    .Z(net109),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1239_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG0 ),
    .Z(net110),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1240_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG1 ),
    .Z(net111),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1241_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG2 ),
    .Z(net112),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1242_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG3 ),
    .Z(net113),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1243_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG0 ),
    .Z(net114),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1244_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG1 ),
    .Z(net115),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1245_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG2 ),
    .Z(net116),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1246_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG3 ),
    .Z(net117),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1247_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG4 ),
    .Z(net118),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1248_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG5 ),
    .Z(net119),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1249_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG6 ),
    .Z(net120),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1250_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG7 ),
    .Z(net121),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1251_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb0 ),
    .Z(net122),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1252_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb1 ),
    .Z(net123),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1253_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb2 ),
    .Z(net124),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1254_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb3 ),
    .Z(net125),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1255_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb4 ),
    .Z(net126),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1256_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb5 ),
    .Z(net127),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1257_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb6 ),
    .Z(net128),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1258_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb7 ),
    .Z(net129),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1259_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG0 ),
    .Z(net130),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1260_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG1 ),
    .Z(net133),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1261_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG2 ),
    .Z(net134),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1262_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG3 ),
    .Z(net135),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1263_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG4 ),
    .Z(net136),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1264_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG5 ),
    .Z(net137),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1265_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG6 ),
    .Z(net138),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1266_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG7 ),
    .Z(net139),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1267_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG8 ),
    .Z(net140),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1268_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG9 ),
    .Z(net141),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1269_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG10 ),
    .Z(net131),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1270_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG11 ),
    .Z(net132),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1271_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG0 ),
    .Z(net142),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1272_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG1 ),
    .Z(net149),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1273_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG2 ),
    .Z(net150),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1274_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG3 ),
    .Z(net151),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1275_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG4 ),
    .Z(net152),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1276_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG5 ),
    .Z(net153),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1277_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG6 ),
    .Z(net154),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1278_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG7 ),
    .Z(net155),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1279_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG8 ),
    .Z(net156),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1280_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG9 ),
    .Z(net157),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1281_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG10 ),
    .Z(net143),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1282_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG11 ),
    .Z(net144),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1283_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG12 ),
    .Z(net145),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1284_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG13 ),
    .Z(net146),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1285_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG14 ),
    .Z(net147),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1286_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG15 ),
    .Z(net148),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1287_ (.I(Tile_X0Y1_FrameData[0]),
    .Z(net158),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1288_ (.I(Tile_X0Y1_FrameData[1]),
    .Z(net169),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1289_ (.I(Tile_X0Y1_FrameData[2]),
    .Z(net180),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1290_ (.I(Tile_X0Y1_FrameData[3]),
    .Z(net183),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1291_ (.I(Tile_X0Y1_FrameData[4]),
    .Z(net184),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1292_ (.I(Tile_X0Y1_FrameData[5]),
    .Z(net185),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1293_ (.I(Tile_X0Y1_FrameData[6]),
    .Z(net186),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1294_ (.I(Tile_X0Y1_FrameData[7]),
    .Z(net187),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1295_ (.I(Tile_X0Y1_FrameData[8]),
    .Z(net188),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1296_ (.I(Tile_X0Y1_FrameData[9]),
    .Z(net189),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1297_ (.I(Tile_X0Y1_FrameData[10]),
    .Z(net159),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1298_ (.I(Tile_X0Y1_FrameData[11]),
    .Z(net160),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1299_ (.I(Tile_X0Y1_FrameData[12]),
    .Z(net161),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1300_ (.I(Tile_X0Y1_FrameData[13]),
    .Z(net162),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1301_ (.I(Tile_X0Y1_FrameData[14]),
    .Z(net163),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1302_ (.I(Tile_X0Y1_FrameData[15]),
    .Z(net164),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1303_ (.I(Tile_X0Y1_FrameData[16]),
    .Z(net165),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1304_ (.I(Tile_X0Y1_FrameData[17]),
    .Z(net166),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1305_ (.I(Tile_X0Y1_FrameData[18]),
    .Z(net167),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1306_ (.I(Tile_X0Y1_FrameData[19]),
    .Z(net168),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1307_ (.I(Tile_X0Y1_FrameData[20]),
    .Z(net170),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1308_ (.I(Tile_X0Y1_FrameData[21]),
    .Z(net171),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1309_ (.I(Tile_X0Y1_FrameData[22]),
    .Z(net172),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1310_ (.I(Tile_X0Y1_FrameData[23]),
    .Z(net173),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1311_ (.I(Tile_X0Y1_FrameData[24]),
    .Z(net174),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1312_ (.I(Tile_X0Y1_FrameData[25]),
    .Z(net175),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1313_ (.I(Tile_X0Y1_FrameData[26]),
    .Z(net176),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1314_ (.I(Tile_X0Y1_FrameData[27]),
    .Z(net177),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1315_ (.I(Tile_X0Y1_FrameData[28]),
    .Z(net178),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1316_ (.I(Tile_X0Y1_FrameData[29]),
    .Z(net179),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1317_ (.I(Tile_X0Y1_FrameData[30]),
    .Z(net181),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1318_ (.I(Tile_X0Y1_FrameData[31]),
    .Z(net182),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1319_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG0 ),
    .Z(net190),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1320_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG1 ),
    .Z(net191),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1321_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG2 ),
    .Z(net192),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1322_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG3 ),
    .Z(net193),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1323_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG0 ),
    .Z(net194),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1324_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG1 ),
    .Z(net195),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1325_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG2 ),
    .Z(net196),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1326_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG3 ),
    .Z(net197),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1327_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG4 ),
    .Z(net198),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1328_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG5 ),
    .Z(net199),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1329_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG6 ),
    .Z(net200),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1330_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG7 ),
    .Z(net201),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1331_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG0 ),
    .Z(net202),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1332_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG1 ),
    .Z(net203),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1333_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG2 ),
    .Z(net204),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1334_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG3 ),
    .Z(net205),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1335_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG4 ),
    .Z(net206),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1336_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG5 ),
    .Z(net207),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1337_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG6 ),
    .Z(net208),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1338_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG7 ),
    .Z(net209),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1339_ (.I(Tile_X0Y0_S4END[8]),
    .Z(net210),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1340_ (.I(Tile_X0Y0_S4END[9]),
    .Z(net217),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1341_ (.I(Tile_X0Y0_S4END[10]),
    .Z(net218),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1342_ (.I(Tile_X0Y0_S4END[11]),
    .Z(net219),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1343_ (.I(Tile_X0Y0_S4END[12]),
    .Z(net220),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1344_ (.I(Tile_X0Y0_S4END[13]),
    .Z(net221),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1345_ (.I(Tile_X0Y0_S4END[14]),
    .Z(net222),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1346_ (.I(Tile_X0Y0_S4END[15]),
    .Z(net223),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1347_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG0 ),
    .Z(net224),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1348_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG1 ),
    .Z(net225),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1349_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG2 ),
    .Z(net211),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1350_ (.I(\Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG3 ),
    .Z(net212),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1351_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG0 ),
    .Z(net213),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1352_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG1 ),
    .Z(net214),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1353_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG2 ),
    .Z(net215),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1354_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG3 ),
    .Z(net216),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1355_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG0 ),
    .Z(net226),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1356_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG1 ),
    .Z(net227),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1357_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG2 ),
    .Z(net228),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1358_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG3 ),
    .Z(net229),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1359_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG0 ),
    .Z(net230),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1360_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG1 ),
    .Z(net231),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1361_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG2 ),
    .Z(net232),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1362_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG3 ),
    .Z(net233),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1363_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG4 ),
    .Z(net234),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1364_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG5 ),
    .Z(net235),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1365_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG6 ),
    .Z(net236),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1366_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG7 ),
    .Z(net237),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1367_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb0 ),
    .Z(net238),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1368_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb1 ),
    .Z(net239),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1369_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb2 ),
    .Z(net240),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1370_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb3 ),
    .Z(net241),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1371_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb4 ),
    .Z(net242),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1372_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb5 ),
    .Z(net243),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1373_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb6 ),
    .Z(net244),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1374_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb7 ),
    .Z(net245),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1375_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG0 ),
    .Z(net246),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1376_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG1 ),
    .Z(net249),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1377_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG2 ),
    .Z(net250),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1378_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG3 ),
    .Z(net251),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1379_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG4 ),
    .Z(net252),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1380_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG5 ),
    .Z(net253),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1381_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG6 ),
    .Z(net254),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1382_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG7 ),
    .Z(net255),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1383_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG8 ),
    .Z(net256),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1384_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG9 ),
    .Z(net257),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1385_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG10 ),
    .Z(net247),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1386_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG11 ),
    .Z(net248),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1387_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG0 ),
    .Z(net258),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1388_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG1 ),
    .Z(net265),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1389_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG2 ),
    .Z(net266),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1390_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG3 ),
    .Z(net267),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1391_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG4 ),
    .Z(net268),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1392_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG5 ),
    .Z(net269),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1393_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG6 ),
    .Z(net270),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1394_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG7 ),
    .Z(net271),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1395_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG8 ),
    .Z(net272),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1396_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG9 ),
    .Z(net273),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1397_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG10 ),
    .Z(net259),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1398_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG11 ),
    .Z(net260),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1399_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG12 ),
    .Z(net261),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1400_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG13 ),
    .Z(net262),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1401_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG14 ),
    .Z(net263),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1402_ (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG15 ),
    .Z(net264),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_144 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_145 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_146 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_147 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_148 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_149 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_150 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_151 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_152 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_153 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_154 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_155 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_156 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_157 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_158 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_159 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_160 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_161 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_162 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_163 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_164 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_165 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_166 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_167 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_168 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_169 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_170 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_171 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_172 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_173 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_174 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_175 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_176 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_177 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_178 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_179 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_180 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_181 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_182 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_183 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_184 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_185 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_186 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_187 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_188 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_189 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_190 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_191 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_192 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_193 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_194 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_195 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_196 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_197 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_198 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_199 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_200 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_201 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_202 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_203 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_204 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_205 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_206 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_207 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_208 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_209 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_210 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_211 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_212 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_213 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_214 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_215 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_216 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_217 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_218 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_219 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_220 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_221 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_222 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_223 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_224 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_225 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_226 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_227 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_228 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_229 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_230 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_231 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_232 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_233 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_234 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_235 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_236 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_237 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_238 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_239 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_240 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_241 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_242 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_243 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_244 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_245 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_246 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_247 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_248 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_249 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_250 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_251 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_252 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_253 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_254 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_255 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_256 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_257 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_258 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_259 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_260 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_261 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_262 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_263 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_264 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_265 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_266 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_267 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_268 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_269 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_270 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_271 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_272 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_273 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_274 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_275 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_276 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_277 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_278 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_279 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_280 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_281 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_282 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_283 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_284 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_285 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_286 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_287 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_288 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_289 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_290 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_291 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_292 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_293 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_294 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_295 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_296 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_297 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_298 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_299 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_300 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_301 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_302 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_303 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_304 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_305 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_306 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_307 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_308 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_309 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_310 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_311 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_312 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_313 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_314 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_315 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_316 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_317 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_318 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_319 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_320 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_321 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_322 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_323 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_324 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_325 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_326 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_327 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_328 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_329 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_330 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_331 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_332 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_333 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_334 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_335 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_336 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_337 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_338 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_339 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_340 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_341 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_342 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_343 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_344 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_345 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_346 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_347 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_348 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_349 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_350 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_351 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_352 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_353 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_354 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_355 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_356 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_357 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_358 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_359 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_360 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_361 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_362 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_363 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_364 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_365 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_366 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_367 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_368 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_369 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_370 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_371 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_372 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_373 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_374 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_375 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_376 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_377 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_378 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_379 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_380 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_381 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_382 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_383 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_384 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_385 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_386 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_387 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_388 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_389 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_390 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_391 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_392 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_393 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_394 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_395 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_396 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_397 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_398 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_399 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_400 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_401 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_402 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_403 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_404 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_405 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_406 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_407 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_408 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_409 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_410 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_411 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_412 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_413 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_414 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_415 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_416 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_417 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_418 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_419 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_420 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_421 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_422 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_423 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_424 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_425 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_426 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_427 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_428 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_429 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_430 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_431 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_432 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_433 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_434 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_435 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_436 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_437 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_438 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_439 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_440 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_441 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_442 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_443 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_444 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_445 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_446 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_447 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_448 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_449 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_450 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_451 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_452 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_453 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_454 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_455 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_456 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_457 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_458 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_459 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_460 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_461 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_462 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_463 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_464 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_465 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_466 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_467 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_468 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_469 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_470 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_471 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_472 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_473 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_474 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_475 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_476 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_477 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_478 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_479 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_480 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_481 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_482 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_483 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_484 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_485 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_486 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_487 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_488 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_489 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_490 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_491 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_492 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_493 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_494 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_495 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_496 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_497 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_498 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_499 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_500 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_501 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_502 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_503 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_504 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_505 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_506 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_507 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_508 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_509 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_510 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_511 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_512 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_513 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_514 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_515 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_516 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_517 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_518 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_519 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_520 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_521 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_522 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_523 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_524 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_525 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_526 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_527 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_528 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_529 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_530 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_531 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_532 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_533 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_534 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_535 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_536 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_537 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_538 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_539 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_540 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_541 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_542 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_543 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_544 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_545 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_546 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_547 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_548 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_549 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_550 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_551 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_552 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_553 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_554 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_555 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_556 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_557 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_558 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_559 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_560 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_561 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_562 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_563 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_564 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_565 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_566 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_567 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_568 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_569 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_570 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_571 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_572 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_573 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_574 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_575 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_576 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_577 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_578 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_579 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_580 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_581 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_582 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_583 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_584 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_585 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_586 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_587 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_588 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_589 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_590 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_591 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_592 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_593 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_594 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_595 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_596 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_597 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_598 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_599 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_600 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_601 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_602 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_603 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_604 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_605 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_606 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_607 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_608 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_609 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_610 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_611 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_612 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_613 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_614 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_615 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_616 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_617 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_618 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_619 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_620 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_621 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_622 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_623 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_624 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_625 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_626 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_627 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_628 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_629 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_630 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_631 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_632 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_633 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_634 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_635 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_636 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_637 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_638 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_639 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_640 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_641 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_642 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_643 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_644 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_645 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_646 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_647 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_648 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_649 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_650 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_651 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_652 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_653 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_654 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_655 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_656 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_657 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_658 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_659 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_660 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_661 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_662 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_663 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_664 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_665 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_666 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_667 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_668 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_669 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_670 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_671 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_672 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_673 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_674 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_675 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_676 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_677 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_678 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_679 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_680 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_681 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_682 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_683 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_684 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_685 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_686 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_687 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_688 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_689 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_690 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_691 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_692 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_693 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_694 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_695 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_696 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_697 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_698 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_699 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_700 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_701 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_702 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_703 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_704 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_705 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_706 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_707 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_708 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_709 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_710 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_711 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_712 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_713 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_714 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_715 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_716 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_717 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_718 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_719 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_720 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_721 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_722 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_723 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_724 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_725 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_726 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_727 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_728 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_729 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_730 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_731 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_732 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_733 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_734 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_735 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_736 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_737 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_738 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_739 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_740 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_741 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_742 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_743 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_744 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_745 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_746 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_747 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_748 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_749 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_750 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_751 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_752 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_753 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_754 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_755 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_756 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_757 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_758 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_759 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_760 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_761 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_762 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_763 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_764 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_765 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_766 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_767 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_768 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_769 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_770 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_771 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_772 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_773 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_774 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_775 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_776 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_777 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_778 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_779 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_780 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_781 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_782 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_783 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_784 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_785 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_786 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_787 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_788 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_789 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_790 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_791 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_792 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_793 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_794 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_795 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_796 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_797 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_798 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output1 (.I(net1),
    .Z(A_SRAM0),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output2 (.I(net2),
    .Z(A_SRAM1),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output3 (.I(net3),
    .Z(A_SRAM2),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output4 (.I(net4),
    .Z(A_SRAM3),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output5 (.I(net5),
    .Z(A_SRAM4),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output6 (.I(net6),
    .Z(A_SRAM5),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output7 (.I(net7),
    .Z(A_SRAM6),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output8 (.I(net8),
    .Z(A_SRAM7),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output9 (.I(net9),
    .Z(A_SRAM8),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output10 (.I(net10),
    .Z(CEN_SRAM),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output11 (.I(net11),
    .Z(CLK_SRAM),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output12 (.I(net12),
    .Z(D_SRAM0),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output13 (.I(net13),
    .Z(D_SRAM1),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output14 (.I(net14),
    .Z(D_SRAM2),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output15 (.I(net15),
    .Z(D_SRAM3),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output16 (.I(net16),
    .Z(D_SRAM4),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output17 (.I(net17),
    .Z(D_SRAM5),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output18 (.I(net18),
    .Z(D_SRAM6),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output19 (.I(net19),
    .Z(D_SRAM7),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output20 (.I(net20),
    .Z(GWEN_SRAM),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output21 (.I(net21),
    .Z(Tile_X0Y0_FrameData_O[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output22 (.I(net22),
    .Z(Tile_X0Y0_FrameData_O[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output23 (.I(net23),
    .Z(Tile_X0Y0_FrameData_O[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output24 (.I(net24),
    .Z(Tile_X0Y0_FrameData_O[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output25 (.I(net25),
    .Z(Tile_X0Y0_FrameData_O[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output26 (.I(net26),
    .Z(Tile_X0Y0_FrameData_O[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output27 (.I(net27),
    .Z(Tile_X0Y0_FrameData_O[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output28 (.I(net28),
    .Z(Tile_X0Y0_FrameData_O[16]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output29 (.I(net29),
    .Z(Tile_X0Y0_FrameData_O[17]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output30 (.I(net30),
    .Z(Tile_X0Y0_FrameData_O[18]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output31 (.I(net31),
    .Z(Tile_X0Y0_FrameData_O[19]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output32 (.I(net32),
    .Z(Tile_X0Y0_FrameData_O[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output33 (.I(net33),
    .Z(Tile_X0Y0_FrameData_O[20]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output34 (.I(net34),
    .Z(Tile_X0Y0_FrameData_O[21]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output35 (.I(net35),
    .Z(Tile_X0Y0_FrameData_O[22]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output36 (.I(net36),
    .Z(Tile_X0Y0_FrameData_O[23]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output37 (.I(net37),
    .Z(Tile_X0Y0_FrameData_O[24]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output38 (.I(net38),
    .Z(Tile_X0Y0_FrameData_O[25]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output39 (.I(net39),
    .Z(Tile_X0Y0_FrameData_O[26]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output40 (.I(net40),
    .Z(Tile_X0Y0_FrameData_O[27]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output41 (.I(net41),
    .Z(Tile_X0Y0_FrameData_O[28]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output42 (.I(net42),
    .Z(Tile_X0Y0_FrameData_O[29]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output43 (.I(net43),
    .Z(Tile_X0Y0_FrameData_O[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output44 (.I(net44),
    .Z(Tile_X0Y0_FrameData_O[30]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output45 (.I(net45),
    .Z(Tile_X0Y0_FrameData_O[31]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output46 (.I(net46),
    .Z(Tile_X0Y0_FrameData_O[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output47 (.I(net47),
    .Z(Tile_X0Y0_FrameData_O[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output48 (.I(net48),
    .Z(Tile_X0Y0_FrameData_O[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output49 (.I(net49),
    .Z(Tile_X0Y0_FrameData_O[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output50 (.I(net50),
    .Z(Tile_X0Y0_FrameData_O[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output51 (.I(net51),
    .Z(Tile_X0Y0_FrameData_O[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output52 (.I(net52),
    .Z(Tile_X0Y0_FrameData_O[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output53 (.I(net53),
    .Z(Tile_X0Y0_FrameStrobe_O[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output54 (.I(net54),
    .Z(Tile_X0Y0_FrameStrobe_O[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output55 (.I(net55),
    .Z(Tile_X0Y0_FrameStrobe_O[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output56 (.I(net56),
    .Z(Tile_X0Y0_FrameStrobe_O[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output57 (.I(net57),
    .Z(Tile_X0Y0_FrameStrobe_O[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output58 (.I(net58),
    .Z(Tile_X0Y0_FrameStrobe_O[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output59 (.I(net59),
    .Z(Tile_X0Y0_FrameStrobe_O[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output60 (.I(net60),
    .Z(Tile_X0Y0_FrameStrobe_O[16]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output61 (.I(net61),
    .Z(Tile_X0Y0_FrameStrobe_O[17]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output62 (.I(net62),
    .Z(Tile_X0Y0_FrameStrobe_O[18]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output63 (.I(net63),
    .Z(Tile_X0Y0_FrameStrobe_O[19]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output64 (.I(net64),
    .Z(Tile_X0Y0_FrameStrobe_O[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output65 (.I(net65),
    .Z(Tile_X0Y0_FrameStrobe_O[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output66 (.I(net66),
    .Z(Tile_X0Y0_FrameStrobe_O[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output67 (.I(net67),
    .Z(Tile_X0Y0_FrameStrobe_O[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output68 (.I(net68),
    .Z(Tile_X0Y0_FrameStrobe_O[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output69 (.I(net69),
    .Z(Tile_X0Y0_FrameStrobe_O[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output70 (.I(net70),
    .Z(Tile_X0Y0_FrameStrobe_O[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output71 (.I(net71),
    .Z(Tile_X0Y0_FrameStrobe_O[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output72 (.I(net72),
    .Z(Tile_X0Y0_FrameStrobe_O[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output73 (.I(net73),
    .Z(Tile_X0Y0_N1BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output74 (.I(net74),
    .Z(Tile_X0Y0_N1BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output75 (.I(net75),
    .Z(Tile_X0Y0_N1BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output76 (.I(net76),
    .Z(Tile_X0Y0_N1BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output77 (.I(net77),
    .Z(Tile_X0Y0_N2BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output78 (.I(net78),
    .Z(Tile_X0Y0_N2BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output79 (.I(net79),
    .Z(Tile_X0Y0_N2BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output80 (.I(net80),
    .Z(Tile_X0Y0_N2BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output81 (.I(net81),
    .Z(Tile_X0Y0_N2BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output82 (.I(net82),
    .Z(Tile_X0Y0_N2BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output83 (.I(net83),
    .Z(Tile_X0Y0_N2BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output84 (.I(net84),
    .Z(Tile_X0Y0_N2BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output85 (.I(net85),
    .Z(Tile_X0Y0_N2BEGb[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output86 (.I(net86),
    .Z(Tile_X0Y0_N2BEGb[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output87 (.I(net87),
    .Z(Tile_X0Y0_N2BEGb[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output88 (.I(net88),
    .Z(Tile_X0Y0_N2BEGb[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output89 (.I(net89),
    .Z(Tile_X0Y0_N2BEGb[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output90 (.I(net90),
    .Z(Tile_X0Y0_N2BEGb[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output91 (.I(net91),
    .Z(Tile_X0Y0_N2BEGb[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output92 (.I(net92),
    .Z(Tile_X0Y0_N2BEGb[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output93 (.I(net93),
    .Z(Tile_X0Y0_N4BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output94 (.I(net94),
    .Z(Tile_X0Y0_N4BEG[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output95 (.I(net95),
    .Z(Tile_X0Y0_N4BEG[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output96 (.I(net96),
    .Z(Tile_X0Y0_N4BEG[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output97 (.I(net97),
    .Z(Tile_X0Y0_N4BEG[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output98 (.I(net98),
    .Z(Tile_X0Y0_N4BEG[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output99 (.I(net99),
    .Z(Tile_X0Y0_N4BEG[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output100 (.I(net100),
    .Z(Tile_X0Y0_N4BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output101 (.I(net101),
    .Z(Tile_X0Y0_N4BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output102 (.I(net102),
    .Z(Tile_X0Y0_N4BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output103 (.I(net103),
    .Z(Tile_X0Y0_N4BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output104 (.I(net104),
    .Z(Tile_X0Y0_N4BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output105 (.I(net105),
    .Z(Tile_X0Y0_N4BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output106 (.I(net106),
    .Z(Tile_X0Y0_N4BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output107 (.I(net107),
    .Z(Tile_X0Y0_N4BEG[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output108 (.I(net108),
    .Z(Tile_X0Y0_N4BEG[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output109 (.I(net109),
    .Z(Tile_X0Y0_UserCLKo),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output110 (.I(net110),
    .Z(Tile_X0Y0_W1BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output111 (.I(net111),
    .Z(Tile_X0Y0_W1BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output112 (.I(net112),
    .Z(Tile_X0Y0_W1BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output113 (.I(net113),
    .Z(Tile_X0Y0_W1BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output114 (.I(net114),
    .Z(Tile_X0Y0_W2BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output115 (.I(net115),
    .Z(Tile_X0Y0_W2BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output116 (.I(net116),
    .Z(Tile_X0Y0_W2BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output117 (.I(net117),
    .Z(Tile_X0Y0_W2BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output118 (.I(net118),
    .Z(Tile_X0Y0_W2BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output119 (.I(net119),
    .Z(Tile_X0Y0_W2BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output120 (.I(net120),
    .Z(Tile_X0Y0_W2BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output121 (.I(net121),
    .Z(Tile_X0Y0_W2BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output122 (.I(net122),
    .Z(Tile_X0Y0_W2BEGb[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output123 (.I(net123),
    .Z(Tile_X0Y0_W2BEGb[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output124 (.I(net124),
    .Z(Tile_X0Y0_W2BEGb[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output125 (.I(net125),
    .Z(Tile_X0Y0_W2BEGb[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output126 (.I(net126),
    .Z(Tile_X0Y0_W2BEGb[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output127 (.I(net127),
    .Z(Tile_X0Y0_W2BEGb[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output128 (.I(net128),
    .Z(Tile_X0Y0_W2BEGb[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output129 (.I(net129),
    .Z(Tile_X0Y0_W2BEGb[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output130 (.I(net130),
    .Z(Tile_X0Y0_W6BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output131 (.I(net131),
    .Z(Tile_X0Y0_W6BEG[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output132 (.I(net132),
    .Z(Tile_X0Y0_W6BEG[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output133 (.I(net133),
    .Z(Tile_X0Y0_W6BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output134 (.I(net134),
    .Z(Tile_X0Y0_W6BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output135 (.I(net135),
    .Z(Tile_X0Y0_W6BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output136 (.I(net136),
    .Z(Tile_X0Y0_W6BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output137 (.I(net137),
    .Z(Tile_X0Y0_W6BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output138 (.I(net138),
    .Z(Tile_X0Y0_W6BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output139 (.I(net139),
    .Z(Tile_X0Y0_W6BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output140 (.I(net140),
    .Z(Tile_X0Y0_W6BEG[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output141 (.I(net141),
    .Z(Tile_X0Y0_W6BEG[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output142 (.I(net142),
    .Z(Tile_X0Y0_WW4BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output143 (.I(net143),
    .Z(Tile_X0Y0_WW4BEG[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output144 (.I(net144),
    .Z(Tile_X0Y0_WW4BEG[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output145 (.I(net145),
    .Z(Tile_X0Y0_WW4BEG[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output146 (.I(net146),
    .Z(Tile_X0Y0_WW4BEG[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output147 (.I(net147),
    .Z(Tile_X0Y0_WW4BEG[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output148 (.I(net148),
    .Z(Tile_X0Y0_WW4BEG[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output149 (.I(net149),
    .Z(Tile_X0Y0_WW4BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output150 (.I(net150),
    .Z(Tile_X0Y0_WW4BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output151 (.I(net151),
    .Z(Tile_X0Y0_WW4BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output152 (.I(net152),
    .Z(Tile_X0Y0_WW4BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output153 (.I(net153),
    .Z(Tile_X0Y0_WW4BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output154 (.I(net154),
    .Z(Tile_X0Y0_WW4BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output155 (.I(net155),
    .Z(Tile_X0Y0_WW4BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output156 (.I(net156),
    .Z(Tile_X0Y0_WW4BEG[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output157 (.I(net157),
    .Z(Tile_X0Y0_WW4BEG[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output158 (.I(net158),
    .Z(Tile_X0Y1_FrameData_O[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output159 (.I(net159),
    .Z(Tile_X0Y1_FrameData_O[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output160 (.I(net160),
    .Z(Tile_X0Y1_FrameData_O[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output161 (.I(net161),
    .Z(Tile_X0Y1_FrameData_O[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output162 (.I(net162),
    .Z(Tile_X0Y1_FrameData_O[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output163 (.I(net163),
    .Z(Tile_X0Y1_FrameData_O[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output164 (.I(net164),
    .Z(Tile_X0Y1_FrameData_O[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output165 (.I(net165),
    .Z(Tile_X0Y1_FrameData_O[16]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output166 (.I(net166),
    .Z(Tile_X0Y1_FrameData_O[17]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output167 (.I(net167),
    .Z(Tile_X0Y1_FrameData_O[18]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output168 (.I(net168),
    .Z(Tile_X0Y1_FrameData_O[19]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output169 (.I(net169),
    .Z(Tile_X0Y1_FrameData_O[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output170 (.I(net170),
    .Z(Tile_X0Y1_FrameData_O[20]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output171 (.I(net171),
    .Z(Tile_X0Y1_FrameData_O[21]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output172 (.I(net172),
    .Z(Tile_X0Y1_FrameData_O[22]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output173 (.I(net173),
    .Z(Tile_X0Y1_FrameData_O[23]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output174 (.I(net174),
    .Z(Tile_X0Y1_FrameData_O[24]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output175 (.I(net175),
    .Z(Tile_X0Y1_FrameData_O[25]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output176 (.I(net176),
    .Z(Tile_X0Y1_FrameData_O[26]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output177 (.I(net177),
    .Z(Tile_X0Y1_FrameData_O[27]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output178 (.I(net178),
    .Z(Tile_X0Y1_FrameData_O[28]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output179 (.I(net179),
    .Z(Tile_X0Y1_FrameData_O[29]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output180 (.I(net180),
    .Z(Tile_X0Y1_FrameData_O[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output181 (.I(net181),
    .Z(Tile_X0Y1_FrameData_O[30]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output182 (.I(net182),
    .Z(Tile_X0Y1_FrameData_O[31]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output183 (.I(net183),
    .Z(Tile_X0Y1_FrameData_O[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output184 (.I(net184),
    .Z(Tile_X0Y1_FrameData_O[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output185 (.I(net185),
    .Z(Tile_X0Y1_FrameData_O[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output186 (.I(net186),
    .Z(Tile_X0Y1_FrameData_O[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output187 (.I(net187),
    .Z(Tile_X0Y1_FrameData_O[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output188 (.I(net188),
    .Z(Tile_X0Y1_FrameData_O[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output189 (.I(net189),
    .Z(Tile_X0Y1_FrameData_O[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output190 (.I(net190),
    .Z(Tile_X0Y1_S1BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output191 (.I(net191),
    .Z(Tile_X0Y1_S1BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output192 (.I(net192),
    .Z(Tile_X0Y1_S1BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output193 (.I(net193),
    .Z(Tile_X0Y1_S1BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output194 (.I(net194),
    .Z(Tile_X0Y1_S2BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output195 (.I(net195),
    .Z(Tile_X0Y1_S2BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output196 (.I(net196),
    .Z(Tile_X0Y1_S2BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output197 (.I(net197),
    .Z(Tile_X0Y1_S2BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output198 (.I(net198),
    .Z(Tile_X0Y1_S2BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output199 (.I(net199),
    .Z(Tile_X0Y1_S2BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output200 (.I(net200),
    .Z(Tile_X0Y1_S2BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output201 (.I(net201),
    .Z(Tile_X0Y1_S2BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output202 (.I(net202),
    .Z(Tile_X0Y1_S2BEGb[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output203 (.I(net203),
    .Z(Tile_X0Y1_S2BEGb[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output204 (.I(net204),
    .Z(Tile_X0Y1_S2BEGb[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output205 (.I(net205),
    .Z(Tile_X0Y1_S2BEGb[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output206 (.I(net206),
    .Z(Tile_X0Y1_S2BEGb[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output207 (.I(net207),
    .Z(Tile_X0Y1_S2BEGb[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output208 (.I(net208),
    .Z(Tile_X0Y1_S2BEGb[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output209 (.I(net209),
    .Z(Tile_X0Y1_S2BEGb[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output210 (.I(net210),
    .Z(Tile_X0Y1_S4BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output211 (.I(net211),
    .Z(Tile_X0Y1_S4BEG[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output212 (.I(net212),
    .Z(Tile_X0Y1_S4BEG[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output213 (.I(net213),
    .Z(Tile_X0Y1_S4BEG[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output214 (.I(net214),
    .Z(Tile_X0Y1_S4BEG[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output215 (.I(net215),
    .Z(Tile_X0Y1_S4BEG[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output216 (.I(net216),
    .Z(Tile_X0Y1_S4BEG[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output217 (.I(net217),
    .Z(Tile_X0Y1_S4BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output218 (.I(net218),
    .Z(Tile_X0Y1_S4BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output219 (.I(net219),
    .Z(Tile_X0Y1_S4BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output220 (.I(net220),
    .Z(Tile_X0Y1_S4BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output221 (.I(net221),
    .Z(Tile_X0Y1_S4BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output222 (.I(net222),
    .Z(Tile_X0Y1_S4BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output223 (.I(net223),
    .Z(Tile_X0Y1_S4BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output224 (.I(net224),
    .Z(Tile_X0Y1_S4BEG[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output225 (.I(net225),
    .Z(Tile_X0Y1_S4BEG[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output226 (.I(net226),
    .Z(Tile_X0Y1_W1BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output227 (.I(net227),
    .Z(Tile_X0Y1_W1BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output228 (.I(net228),
    .Z(Tile_X0Y1_W1BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output229 (.I(net229),
    .Z(Tile_X0Y1_W1BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output230 (.I(net230),
    .Z(Tile_X0Y1_W2BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output231 (.I(net231),
    .Z(Tile_X0Y1_W2BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output232 (.I(net232),
    .Z(Tile_X0Y1_W2BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output233 (.I(net233),
    .Z(Tile_X0Y1_W2BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output234 (.I(net234),
    .Z(Tile_X0Y1_W2BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output235 (.I(net235),
    .Z(Tile_X0Y1_W2BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output236 (.I(net236),
    .Z(Tile_X0Y1_W2BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output237 (.I(net237),
    .Z(Tile_X0Y1_W2BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output238 (.I(net238),
    .Z(Tile_X0Y1_W2BEGb[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output239 (.I(net239),
    .Z(Tile_X0Y1_W2BEGb[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output240 (.I(net240),
    .Z(Tile_X0Y1_W2BEGb[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output241 (.I(net241),
    .Z(Tile_X0Y1_W2BEGb[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output242 (.I(net242),
    .Z(Tile_X0Y1_W2BEGb[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output243 (.I(net243),
    .Z(Tile_X0Y1_W2BEGb[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output244 (.I(net244),
    .Z(Tile_X0Y1_W2BEGb[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output245 (.I(net245),
    .Z(Tile_X0Y1_W2BEGb[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output246 (.I(net246),
    .Z(Tile_X0Y1_W6BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output247 (.I(net247),
    .Z(Tile_X0Y1_W6BEG[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output248 (.I(net248),
    .Z(Tile_X0Y1_W6BEG[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output249 (.I(net249),
    .Z(Tile_X0Y1_W6BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output250 (.I(net250),
    .Z(Tile_X0Y1_W6BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output251 (.I(net251),
    .Z(Tile_X0Y1_W6BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output252 (.I(net252),
    .Z(Tile_X0Y1_W6BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output253 (.I(net253),
    .Z(Tile_X0Y1_W6BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output254 (.I(net254),
    .Z(Tile_X0Y1_W6BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output255 (.I(net255),
    .Z(Tile_X0Y1_W6BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output256 (.I(net256),
    .Z(Tile_X0Y1_W6BEG[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output257 (.I(net257),
    .Z(Tile_X0Y1_W6BEG[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output258 (.I(net258),
    .Z(Tile_X0Y1_WW4BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output259 (.I(net259),
    .Z(Tile_X0Y1_WW4BEG[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output260 (.I(net260),
    .Z(Tile_X0Y1_WW4BEG[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output261 (.I(net261),
    .Z(Tile_X0Y1_WW4BEG[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output262 (.I(net262),
    .Z(Tile_X0Y1_WW4BEG[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output263 (.I(net263),
    .Z(Tile_X0Y1_WW4BEG[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output264 (.I(net264),
    .Z(Tile_X0Y1_WW4BEG[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output265 (.I(net265),
    .Z(Tile_X0Y1_WW4BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output266 (.I(net266),
    .Z(Tile_X0Y1_WW4BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output267 (.I(net267),
    .Z(Tile_X0Y1_WW4BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output268 (.I(net268),
    .Z(Tile_X0Y1_WW4BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output269 (.I(net269),
    .Z(Tile_X0Y1_WW4BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output270 (.I(net270),
    .Z(Tile_X0Y1_WW4BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output271 (.I(net271),
    .Z(Tile_X0Y1_WW4BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output272 (.I(net272),
    .Z(Tile_X0Y1_WW4BEG[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output273 (.I(net273),
    .Z(Tile_X0Y1_WW4BEG[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output274 (.I(net274),
    .Z(WEN_SRAM0),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output275 (.I(net275),
    .Z(WEN_SRAM1),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output276 (.I(net276),
    .Z(WEN_SRAM2),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output277 (.I(net277),
    .Z(WEN_SRAM3),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output278 (.I(net278),
    .Z(WEN_SRAM4),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output279 (.I(net279),
    .Z(WEN_SRAM5),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output280 (.I(net280),
    .Z(WEN_SRAM6),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output281 (.I(net281),
    .Z(WEN_SRAM7),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_Tile_X0Y1_UserCLK (.I(Tile_X0Y1_UserCLK),
    .Z(clknet_0_Tile_X0Y1_UserCLK),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_Tile_X0Y1_UserCLK (.I(clknet_0_Tile_X0Y1_UserCLK),
    .Z(clknet_1_0__leaf_Tile_X0Y1_UserCLK),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_Tile_X0Y1_UserCLK (.I(clknet_0_Tile_X0Y1_UserCLK),
    .Z(clknet_1_1__leaf_Tile_X0Y1_UserCLK),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(Tile_X0Y0_S2END[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(Tile_X0Y0_S2MID[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_3 (.I(Tile_X0Y0_S2MID[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_4 (.I(Tile_X0Y0_S2MID[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_5 (.I(Tile_X0Y0_S2MID[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_6 (.I(Tile_X0Y0_S2MID[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_7 (.I(Tile_X0Y0_S2MID[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_8 (.I(Tile_X0Y1_FrameStrobe[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_9 (.I(Tile_X0Y1_FrameStrobe[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_10 (.I(Tile_X0Y1_FrameStrobe[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_11 (.I(Tile_X0Y1_FrameStrobe[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_12 (.I(Tile_X0Y1_FrameStrobe[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_13 (.I(Tile_X0Y1_FrameStrobe[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_14 (.I(Tile_X0Y1_FrameStrobe[16]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_15 (.I(Tile_X0Y1_FrameStrobe[16]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_16 (.I(Tile_X0Y1_FrameStrobe[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_17 (.I(Tile_X0Y1_N2END[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_18 (.I(Tile_X0Y1_N2END[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_19 (.I(Tile_X0Y1_N2END[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_20 (.I(Tile_X0Y1_N2MID[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_21 (.I(Tile_X0Y1_N2MID[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_22 (.I(Tile_X0Y1_N2MID[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_23 (.I(Tile_X0Y1_N2MID[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_24 (.I(Tile_X0Y1_N2MID[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_25 (.I(Tile_X0Y1_N2MID[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_26 (.I(Tile_X0Y1_N2MID[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_27 (.I(Tile_X0Y1_N2MID[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_28 (.I(Tile_X0Y1_N2MID[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_29 (.I(Tile_X0Y1_N2MID[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_30 (.I(Tile_X0Y1_N4END[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_31 (.I(Tile_X0Y1_N4END[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_32 (.I(Tile_X0Y1_N4END[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_33 (.I(Tile_X0Y1_N4END[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_34 (.I(Tile_X0Y1_N4END[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_35 (.I(Tile_X0Y1_N4END[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_36 (.I(Tile_X0Y1_N4END[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_37 (.I(Tile_X0Y1_N4END[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_38 (.I(Tile_X0Y1_N4END[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_39 (.I(Tile_X0Y1_N4END[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_40 (.I(Tile_X0Y1_N4END[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_41 (.I(Tile_X0Y1_N4END[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_42 (.I(Tile_X0Y1_N4END[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_43 (.I(Tile_X0Y1_N4END[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_44 (.I(Tile_X0Y1_N4END[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_45 (.I(Tile_X0Y1_N4END[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_46 (.I(Tile_X0Y1_FrameStrobe[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_47 (.I(Tile_X0Y1_FrameStrobe[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_48 (.I(Tile_X0Y1_N2MID[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_49 (.I(Tile_X0Y1_N2MID[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_50 (.I(Q_SRAM5),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_51 (.I(Tile_X0Y0_S4END[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_52 (.I(Tile_X0Y1_FrameStrobe[17]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_53 (.I(Tile_X0Y1_FrameStrobe[17]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_54 (.I(Tile_X0Y1_FrameStrobe[18]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_55 (.I(Tile_X0Y1_FrameStrobe[18]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_56 (.I(Tile_X0Y1_FrameStrobe[19]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_57 (.I(Tile_X0Y1_FrameStrobe[19]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_58 (.I(Tile_X0Y1_FrameStrobe[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_59 (.I(\Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_60 (.I(Tile_X0Y1_N4END[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_61 (.I(Tile_X0Y1_N4END[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_62 (.I(net212),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_63 (.I(net225),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_64 (.I(net225),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_65 (.I(net278),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_66 (.I(Tile_X0Y0_S4END[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_67 (.I(Tile_X0Y0_S4END[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_68 (.I(Tile_X0Y0_S4END[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_69 (.I(Tile_X0Y0_S4END[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_70 (.I(Tile_X0Y0_S4END[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_258 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_250 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_236 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_239 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_265 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_240 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_240 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_261 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_256 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_261 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_259 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_239 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_235 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_235 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_236 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_240 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_235 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_239 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_259 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_236 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_245 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_253 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_259 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_265 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_258 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_265 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
endmodule
