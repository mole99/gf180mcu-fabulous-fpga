VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO N_term_single
  CLASS BLOCK ;
  FOREIGN N_term_single ;
  ORIGIN 0.000 0.000 ;
  SIZE 287.280 BY 71.120 ;
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 0.000 120.400 0.560 ;
    END
  END Ci
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 0.000 0.560 0.560 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 22.400 0.560 22.960 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 24.640 0.560 25.200 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 26.880 0.560 27.440 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 29.120 0.560 29.680 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 31.360 0.560 31.920 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.600 0.560 34.160 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 35.840 0.560 36.400 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 38.080 0.560 38.640 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.320 0.560 40.880 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.560 0.560 43.120 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2.240 0.560 2.800 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 44.800 0.560 45.360 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.040 0.560 47.600 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 49.280 0.560 49.840 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 51.520 0.560 52.080 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.760 0.560 54.320 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 56.000 0.560 56.560 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 58.240 0.560 58.800 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.480 0.560 61.040 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 62.720 0.560 63.280 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 64.960 0.560 65.520 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 4.480 0.560 5.040 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 67.200 0.560 67.760 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 69.440 0.560 70.000 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 6.720 0.560 7.280 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 8.960 0.560 9.520 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 11.200 0.560 11.760 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 13.440 0.560 14.000 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.680 0.560 16.240 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 17.920 0.560 18.480 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.160 0.560 20.720 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 0.000 287.280 0.560 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 22.400 287.280 22.960 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 24.640 287.280 25.200 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 26.880 287.280 27.440 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 29.120 287.280 29.680 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 31.360 287.280 31.920 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 33.600 287.280 34.160 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 35.840 287.280 36.400 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 38.080 287.280 38.640 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 40.320 287.280 40.880 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 42.560 287.280 43.120 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 2.240 287.280 2.800 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 44.800 287.280 45.360 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 47.040 287.280 47.600 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 49.280 287.280 49.840 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 51.520 287.280 52.080 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 53.760 287.280 54.320 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 56.000 287.280 56.560 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 58.240 287.280 58.800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 60.480 287.280 61.040 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 62.720 287.280 63.280 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 64.960 287.280 65.520 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 4.480 287.280 5.040 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 67.200 287.280 67.760 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 69.440 287.280 70.000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 6.720 287.280 7.280 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 8.960 287.280 9.520 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 11.200 287.280 11.760 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 13.440 287.280 14.000 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 15.680 287.280 16.240 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 17.920 287.280 18.480 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 20.160 287.280 20.720 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 240.800 0.000 241.360 0.560 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 0.000 263.760 0.560 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 0.000 266.000 0.560 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 0.000 268.240 0.560 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 0.000 270.480 0.560 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 0.000 272.720 0.560 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 274.400 0.000 274.960 0.560 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 0.000 277.200 0.560 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 0.000 279.440 0.560 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 0.000 281.680 0.560 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 283.360 0.000 283.920 0.560 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 243.040 0.000 243.600 0.560 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 0.000 245.840 0.560 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 0.000 248.080 0.560 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 0.000 250.320 0.560 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 0.000 252.560 0.560 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 254.240 0.000 254.800 0.560 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 0.000 257.040 0.560 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 0.000 259.280 0.560 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 0.000 261.520 0.560 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 22.400 70.560 22.960 71.120 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 156.800 70.560 157.360 71.120 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 170.240 70.560 170.800 71.120 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 183.680 70.560 184.240 71.120 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 70.560 197.680 71.120 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 210.560 70.560 211.120 71.120 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 224.000 70.560 224.560 71.120 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 237.440 70.560 238.000 71.120 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 250.880 70.560 251.440 71.120 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 264.320 70.560 264.880 71.120 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 277.760 70.560 278.320 71.120 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 35.840 70.560 36.400 71.120 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 70.560 49.840 71.120 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 70.560 63.280 71.120 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 70.560 76.720 71.120 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 70.560 90.160 71.120 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 70.560 103.600 71.120 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 70.560 117.040 71.120 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 129.920 70.560 130.480 71.120 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 143.360 70.560 143.920 71.120 ;
    END
  END FrameStrobe_O[9]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 0.560 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.600 0.000 6.160 0.560 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.840 0.000 8.400 0.560 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 0.000 10.640 0.560 ;
    END
  END N1END[3]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 0.560 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 0.000 33.040 0.560 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 0.000 35.280 0.560 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 0.560 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 0.000 39.760 0.560 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 0.000 42.000 0.560 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 0.560 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 0.000 46.480 0.560 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 12.320 0.000 12.880 0.560 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 14.560 0.000 15.120 0.560 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 0.000 17.360 0.560 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 19.040 0.000 19.600 0.560 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 21.280 0.000 21.840 0.560 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 0.560 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 0.000 26.320 0.560 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 0.000 28.560 0.560 ;
    END
  END N2MID[7]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 0.000 48.720 0.560 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 0.560 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 0.000 73.360 0.560 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 0.000 75.600 0.560 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 0.560 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 0.000 80.080 0.560 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 0.000 82.320 0.560 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 0.560 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 0.000 53.200 0.560 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 0.000 55.440 0.560 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 0.000 57.680 0.560 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 0.000 59.920 0.560 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 0.000 62.160 0.560 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 0.560 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 0.000 66.640 0.560 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 0.000 68.880 0.560 ;
    END
  END N4END[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 0.560 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 0.000 106.960 0.560 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 0.000 109.200 0.560 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 0.560 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 0.000 113.680 0.560 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 0.000 115.920 0.560 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 0.000 118.160 0.560 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 0.000 86.800 0.560 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 0.000 89.040 0.560 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 0.560 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 0.000 93.520 0.560 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 0.000 95.760 0.560 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 0.560 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 0.000 100.240 0.560 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 0.000 102.480 0.560 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 0.560 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 0.000 122.640 0.560 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 0.560 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 0.000 127.120 0.560 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 0.000 129.360 0.560 ;
    END
  END S1BEG[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 0.560 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 0.000 133.840 0.560 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 0.000 136.080 0.560 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 0.000 138.320 0.560 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 0.000 140.560 0.560 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 0.000 142.800 0.560 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 0.560 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 0.000 147.280 0.560 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 0.000 149.520 0.560 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 0.000 151.760 0.560 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 0.000 154.000 0.560 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 0.000 156.240 0.560 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 0.560 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 0.000 160.720 0.560 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 0.000 162.960 0.560 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 0.560 ;
    END
  END S2BEGb[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 0.560 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 0.000 189.840 0.560 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 0.000 192.080 0.560 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 0.000 194.320 0.560 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 0.000 196.560 0.560 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 0.000 198.800 0.560 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 200.480 0.000 201.040 0.560 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 169.120 0.000 169.680 0.560 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 0.000 171.920 0.560 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 0.000 174.160 0.560 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 0.000 176.400 0.560 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 0.000 178.640 0.560 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 0.000 180.880 0.560 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 0.000 183.120 0.560 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 0.000 185.360 0.560 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 0.000 187.600 0.560 ;
    END
  END S4BEG[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 0.000 203.280 0.560 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 0.000 225.680 0.560 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 0.000 227.920 0.560 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 0.000 230.160 0.560 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 0.000 232.400 0.560 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 0.000 234.640 0.560 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 0.000 236.880 0.560 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 0.000 205.520 0.560 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 0.000 207.760 0.560 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 0.000 210.000 0.560 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 0.560 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 0.000 214.480 0.560 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 216.160 0.000 216.720 0.560 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 0.000 218.960 0.560 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 220.640 0.000 221.200 0.560 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 0.000 223.440 0.560 ;
    END
  END SS4BEG[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 0.000 239.120 0.560 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 8.960 70.560 9.520 71.120 ;
    END
  END UserCLKo
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.880 0.000 20.480 71.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 118.880 0.000 120.480 71.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.880 0.000 220.480 71.120 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.180 0.000 23.780 71.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.180 0.000 123.780 71.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 222.180 0.000 223.780 71.120 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 2.930 3.490 284.350 67.070 ;
      LAYER Metal1 ;
        RECT 3.360 3.620 283.920 66.940 ;
      LAYER Metal2 ;
        RECT 1.820 70.260 8.660 70.560 ;
        RECT 9.820 70.260 22.100 70.560 ;
        RECT 23.260 70.260 35.540 70.560 ;
        RECT 36.700 70.260 48.980 70.560 ;
        RECT 50.140 70.260 62.420 70.560 ;
        RECT 63.580 70.260 75.860 70.560 ;
        RECT 77.020 70.260 89.300 70.560 ;
        RECT 90.460 70.260 102.740 70.560 ;
        RECT 103.900 70.260 116.180 70.560 ;
        RECT 117.340 70.260 129.620 70.560 ;
        RECT 130.780 70.260 143.060 70.560 ;
        RECT 144.220 70.260 156.500 70.560 ;
        RECT 157.660 70.260 169.940 70.560 ;
        RECT 171.100 70.260 183.380 70.560 ;
        RECT 184.540 70.260 196.820 70.560 ;
        RECT 197.980 70.260 210.260 70.560 ;
        RECT 211.420 70.260 223.700 70.560 ;
        RECT 224.860 70.260 237.140 70.560 ;
        RECT 238.300 70.260 250.580 70.560 ;
        RECT 251.740 70.260 264.020 70.560 ;
        RECT 265.180 70.260 277.460 70.560 ;
        RECT 278.620 70.260 286.580 70.560 ;
        RECT 1.820 0.860 286.580 70.260 ;
        RECT 1.820 0.090 3.060 0.860 ;
        RECT 4.220 0.090 5.300 0.860 ;
        RECT 6.460 0.090 7.540 0.860 ;
        RECT 8.700 0.090 9.780 0.860 ;
        RECT 10.940 0.090 12.020 0.860 ;
        RECT 13.180 0.090 14.260 0.860 ;
        RECT 15.420 0.090 16.500 0.860 ;
        RECT 17.660 0.090 18.740 0.860 ;
        RECT 19.900 0.090 20.980 0.860 ;
        RECT 22.140 0.090 23.220 0.860 ;
        RECT 24.380 0.090 25.460 0.860 ;
        RECT 26.620 0.090 27.700 0.860 ;
        RECT 28.860 0.090 29.940 0.860 ;
        RECT 31.100 0.090 32.180 0.860 ;
        RECT 33.340 0.090 34.420 0.860 ;
        RECT 35.580 0.090 36.660 0.860 ;
        RECT 37.820 0.090 38.900 0.860 ;
        RECT 40.060 0.090 41.140 0.860 ;
        RECT 42.300 0.090 43.380 0.860 ;
        RECT 44.540 0.090 45.620 0.860 ;
        RECT 46.780 0.090 47.860 0.860 ;
        RECT 49.020 0.090 50.100 0.860 ;
        RECT 51.260 0.090 52.340 0.860 ;
        RECT 53.500 0.090 54.580 0.860 ;
        RECT 55.740 0.090 56.820 0.860 ;
        RECT 57.980 0.090 59.060 0.860 ;
        RECT 60.220 0.090 61.300 0.860 ;
        RECT 62.460 0.090 63.540 0.860 ;
        RECT 64.700 0.090 65.780 0.860 ;
        RECT 66.940 0.090 68.020 0.860 ;
        RECT 69.180 0.090 70.260 0.860 ;
        RECT 71.420 0.090 72.500 0.860 ;
        RECT 73.660 0.090 74.740 0.860 ;
        RECT 75.900 0.090 76.980 0.860 ;
        RECT 78.140 0.090 79.220 0.860 ;
        RECT 80.380 0.090 81.460 0.860 ;
        RECT 82.620 0.090 83.700 0.860 ;
        RECT 84.860 0.090 85.940 0.860 ;
        RECT 87.100 0.090 88.180 0.860 ;
        RECT 89.340 0.090 90.420 0.860 ;
        RECT 91.580 0.090 92.660 0.860 ;
        RECT 93.820 0.090 94.900 0.860 ;
        RECT 96.060 0.090 97.140 0.860 ;
        RECT 98.300 0.090 99.380 0.860 ;
        RECT 100.540 0.090 101.620 0.860 ;
        RECT 102.780 0.090 103.860 0.860 ;
        RECT 105.020 0.090 106.100 0.860 ;
        RECT 107.260 0.090 108.340 0.860 ;
        RECT 109.500 0.090 110.580 0.860 ;
        RECT 111.740 0.090 112.820 0.860 ;
        RECT 113.980 0.090 115.060 0.860 ;
        RECT 116.220 0.090 117.300 0.860 ;
        RECT 118.460 0.090 119.540 0.860 ;
        RECT 120.700 0.090 121.780 0.860 ;
        RECT 122.940 0.090 124.020 0.860 ;
        RECT 125.180 0.090 126.260 0.860 ;
        RECT 127.420 0.090 128.500 0.860 ;
        RECT 129.660 0.090 130.740 0.860 ;
        RECT 131.900 0.090 132.980 0.860 ;
        RECT 134.140 0.090 135.220 0.860 ;
        RECT 136.380 0.090 137.460 0.860 ;
        RECT 138.620 0.090 139.700 0.860 ;
        RECT 140.860 0.090 141.940 0.860 ;
        RECT 143.100 0.090 144.180 0.860 ;
        RECT 145.340 0.090 146.420 0.860 ;
        RECT 147.580 0.090 148.660 0.860 ;
        RECT 149.820 0.090 150.900 0.860 ;
        RECT 152.060 0.090 153.140 0.860 ;
        RECT 154.300 0.090 155.380 0.860 ;
        RECT 156.540 0.090 157.620 0.860 ;
        RECT 158.780 0.090 159.860 0.860 ;
        RECT 161.020 0.090 162.100 0.860 ;
        RECT 163.260 0.090 164.340 0.860 ;
        RECT 165.500 0.090 166.580 0.860 ;
        RECT 167.740 0.090 168.820 0.860 ;
        RECT 169.980 0.090 171.060 0.860 ;
        RECT 172.220 0.090 173.300 0.860 ;
        RECT 174.460 0.090 175.540 0.860 ;
        RECT 176.700 0.090 177.780 0.860 ;
        RECT 178.940 0.090 180.020 0.860 ;
        RECT 181.180 0.090 182.260 0.860 ;
        RECT 183.420 0.090 184.500 0.860 ;
        RECT 185.660 0.090 186.740 0.860 ;
        RECT 187.900 0.090 188.980 0.860 ;
        RECT 190.140 0.090 191.220 0.860 ;
        RECT 192.380 0.090 193.460 0.860 ;
        RECT 194.620 0.090 195.700 0.860 ;
        RECT 196.860 0.090 197.940 0.860 ;
        RECT 199.100 0.090 200.180 0.860 ;
        RECT 201.340 0.090 202.420 0.860 ;
        RECT 203.580 0.090 204.660 0.860 ;
        RECT 205.820 0.090 206.900 0.860 ;
        RECT 208.060 0.090 209.140 0.860 ;
        RECT 210.300 0.090 211.380 0.860 ;
        RECT 212.540 0.090 213.620 0.860 ;
        RECT 214.780 0.090 215.860 0.860 ;
        RECT 217.020 0.090 218.100 0.860 ;
        RECT 219.260 0.090 220.340 0.860 ;
        RECT 221.500 0.090 222.580 0.860 ;
        RECT 223.740 0.090 224.820 0.860 ;
        RECT 225.980 0.090 227.060 0.860 ;
        RECT 228.220 0.090 229.300 0.860 ;
        RECT 230.460 0.090 231.540 0.860 ;
        RECT 232.700 0.090 233.780 0.860 ;
        RECT 234.940 0.090 236.020 0.860 ;
        RECT 237.180 0.090 238.260 0.860 ;
        RECT 239.420 0.090 240.500 0.860 ;
        RECT 241.660 0.090 242.740 0.860 ;
        RECT 243.900 0.090 244.980 0.860 ;
        RECT 246.140 0.090 247.220 0.860 ;
        RECT 248.380 0.090 249.460 0.860 ;
        RECT 250.620 0.090 251.700 0.860 ;
        RECT 252.860 0.090 253.940 0.860 ;
        RECT 255.100 0.090 256.180 0.860 ;
        RECT 257.340 0.090 258.420 0.860 ;
        RECT 259.580 0.090 260.660 0.860 ;
        RECT 261.820 0.090 262.900 0.860 ;
        RECT 264.060 0.090 265.140 0.860 ;
        RECT 266.300 0.090 267.380 0.860 ;
        RECT 268.540 0.090 269.620 0.860 ;
        RECT 270.780 0.090 271.860 0.860 ;
        RECT 273.020 0.090 274.100 0.860 ;
        RECT 275.260 0.090 276.340 0.860 ;
        RECT 277.500 0.090 278.580 0.860 ;
        RECT 279.740 0.090 280.820 0.860 ;
        RECT 281.980 0.090 283.060 0.860 ;
        RECT 284.220 0.090 286.580 0.860 ;
      LAYER Metal3 ;
        RECT 0.560 70.300 286.720 70.420 ;
        RECT 0.860 69.140 286.420 70.300 ;
        RECT 0.560 68.060 286.720 69.140 ;
        RECT 0.860 66.900 286.420 68.060 ;
        RECT 0.560 65.820 286.720 66.900 ;
        RECT 0.860 64.660 286.420 65.820 ;
        RECT 0.560 63.580 286.720 64.660 ;
        RECT 0.860 62.420 286.420 63.580 ;
        RECT 0.560 61.340 286.720 62.420 ;
        RECT 0.860 60.180 286.420 61.340 ;
        RECT 0.560 59.100 286.720 60.180 ;
        RECT 0.860 57.940 286.420 59.100 ;
        RECT 0.560 56.860 286.720 57.940 ;
        RECT 0.860 55.700 286.420 56.860 ;
        RECT 0.560 54.620 286.720 55.700 ;
        RECT 0.860 53.460 286.420 54.620 ;
        RECT 0.560 52.380 286.720 53.460 ;
        RECT 0.860 51.220 286.420 52.380 ;
        RECT 0.560 50.140 286.720 51.220 ;
        RECT 0.860 48.980 286.420 50.140 ;
        RECT 0.560 47.900 286.720 48.980 ;
        RECT 0.860 46.740 286.420 47.900 ;
        RECT 0.560 45.660 286.720 46.740 ;
        RECT 0.860 44.500 286.420 45.660 ;
        RECT 0.560 43.420 286.720 44.500 ;
        RECT 0.860 42.260 286.420 43.420 ;
        RECT 0.560 41.180 286.720 42.260 ;
        RECT 0.860 40.020 286.420 41.180 ;
        RECT 0.560 38.940 286.720 40.020 ;
        RECT 0.860 37.780 286.420 38.940 ;
        RECT 0.560 36.700 286.720 37.780 ;
        RECT 0.860 35.540 286.420 36.700 ;
        RECT 0.560 34.460 286.720 35.540 ;
        RECT 0.860 33.300 286.420 34.460 ;
        RECT 0.560 32.220 286.720 33.300 ;
        RECT 0.860 31.060 286.420 32.220 ;
        RECT 0.560 29.980 286.720 31.060 ;
        RECT 0.860 28.820 286.420 29.980 ;
        RECT 0.560 27.740 286.720 28.820 ;
        RECT 0.860 26.580 286.420 27.740 ;
        RECT 0.560 25.500 286.720 26.580 ;
        RECT 0.860 24.340 286.420 25.500 ;
        RECT 0.560 23.260 286.720 24.340 ;
        RECT 0.860 22.100 286.420 23.260 ;
        RECT 0.560 21.020 286.720 22.100 ;
        RECT 0.860 19.860 286.420 21.020 ;
        RECT 0.560 18.780 286.720 19.860 ;
        RECT 0.860 17.620 286.420 18.780 ;
        RECT 0.560 16.540 286.720 17.620 ;
        RECT 0.860 15.380 286.420 16.540 ;
        RECT 0.560 14.300 286.720 15.380 ;
        RECT 0.860 13.140 286.420 14.300 ;
        RECT 0.560 12.060 286.720 13.140 ;
        RECT 0.860 10.900 286.420 12.060 ;
        RECT 0.560 9.820 286.720 10.900 ;
        RECT 0.860 8.660 286.420 9.820 ;
        RECT 0.560 7.580 286.720 8.660 ;
        RECT 0.860 6.420 286.420 7.580 ;
        RECT 0.560 5.340 286.720 6.420 ;
        RECT 0.860 4.180 286.420 5.340 ;
        RECT 0.560 3.100 286.720 4.180 ;
        RECT 0.860 1.940 286.420 3.100 ;
        RECT 0.560 0.860 286.720 1.940 ;
        RECT 0.860 0.140 286.420 0.860 ;
      LAYER Metal4 ;
        RECT 20.860 0.090 21.880 62.630 ;
        RECT 24.080 0.090 118.580 62.630 ;
        RECT 120.780 0.090 121.880 62.630 ;
        RECT 124.080 0.090 218.580 62.630 ;
        RECT 220.780 0.090 221.880 62.630 ;
        RECT 224.080 0.090 224.420 62.630 ;
  END
END N_term_single
END LIBRARY

